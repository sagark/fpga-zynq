module BTB(input clk, input reset,
    input  io_req_valid,
    input [42:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output[42:0] io_resp_bits_target,
    output[5:0] io_resp_bits_entry,
    output[6:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_update_valid,
    input  io_update_bits_prediction_valid,
    input  io_update_bits_prediction_bits_taken,
    input [42:0] io_update_bits_prediction_bits_target,
    input [5:0] io_update_bits_prediction_bits_entry,
    input [6:0] io_update_bits_prediction_bits_bht_history,
    input [1:0] io_update_bits_prediction_bits_bht_value,
    input [42:0] io_update_bits_pc,
    input [42:0] io_update_bits_target,
    input [42:0] io_update_bits_returnAddr,
    input  io_update_bits_taken,
    input  io_update_bits_isJump,
    input  io_update_bits_isCall,
    input  io_update_bits_isReturn,
    input  io_update_bits_mispredict,
    input  io_invalidate
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg [42:0] R4;
  wire[42:0] T5;
  wire T6;
  wire T7;
  wire updateTarget;
  reg  R8;
  wire T9;
  wire T10;
  reg  R11;
  wire T12;
  wire updateValid;
  reg  updateHit;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  R18;
  wire T1590;
  wire[1:0] T19;
  wire[1:0] T20;
  reg [1:0] T21 [127:0];
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  reg [6:0] R38;
  wire[6:0] T39;
  wire[6:0] T40;
  wire[6:0] T41;
  wire[5:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[61:0] T47;
  reg [61:0] isJump;
  wire[61:0] T1591;
  wire[63:0] T48;
  wire[63:0] T1592;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T1593;
  wire[61:0] T52;
  wire[63:0] T53;
  wire[5:0] T54;
  reg [5:0] R55;
  wire[5:0] T1594;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg [5:0] R63;
  wire[5:0] T64;
  wire[63:0] T1595;
  wire T65;
  wire T66;
  reg  R67;
  wire T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T1596;
  wire[61:0] hits;
  wire[61:0] T71;
  wire[61:0] T72;
  wire[30:0] T73;
  wire[15:0] T74;
  wire[7:0] T75;
  wire[3:0] T76;
  wire[1:0] T77;
  wire T78;
  wire[5:0] T79;
  wire[5:0] pageHit;
  reg [5:0] pageValid;
  wire[5:0] T1597;
  wire[7:0] T1598;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T1599;
  wire[7:0] T82;
  wire[7:0] pageReplEn;
  wire[7:0] tgtPageReplEn;
  wire[7:0] tgtPageRepl;
  wire[7:0] T1600;
  wire[5:0] T83;
  wire[5:0] T1601;
  wire T84;
  wire[5:0] T85;
  wire[4:0] T86;
  wire[7:0] idxPageUpdateOH;
  wire[7:0] idxPageRepl;
  wire[7:0] T87;
  reg [2:0] R88;
  wire[2:0] T1602;
  wire[2:0] T89;
  wire[2:0] T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire T94;
  wire[7:0] T1603;
  wire[5:0] updatePageHit;
  wire[5:0] T95;
  wire[5:0] T96;
  wire[2:0] T97;
  wire[1:0] T98;
  wire T99;
  wire[29:0] T100;
  reg [42:0] R101;
  wire[42:0] T102;
  wire[29:0] T103;
  reg [29:0] pages [5:0];
  wire[29:0] T104;
  wire[29:0] T105;
  wire[29:0] T106;
  wire[29:0] T107;
  wire T108;
  wire[7:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire[29:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire[29:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[29:0] T122;
  wire[29:0] T123;
  wire[29:0] T124;
  wire[29:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire[29:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[29:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[29:0] T139;
  wire T140;
  wire[29:0] T141;
  wire[2:0] T142;
  wire[1:0] T143;
  wire T144;
  wire[29:0] T145;
  wire T146;
  wire[29:0] T147;
  wire T148;
  wire[29:0] T149;
  wire useUpdatePageHit;
  wire samePage;
  wire[29:0] T150;
  wire[29:0] T151;
  wire doTgtPageRepl;
  wire T152;
  wire usePageHit;
  wire[7:0] T153;
  wire[7:0] T154;
  wire[7:0] T1604;
  wire T155;
  wire T156;
  wire[7:0] idxPageReplEn;
  wire[7:0] T1605;
  wire T157;
  wire[5:0] T158;
  wire[5:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[29:0] T163;
  wire[29:0] T164;
  wire T165;
  wire[29:0] T166;
  wire T167;
  wire[29:0] T168;
  wire[2:0] T169;
  wire[1:0] T170;
  wire T171;
  wire[29:0] T172;
  wire T173;
  wire[29:0] T174;
  wire T175;
  wire[29:0] T176;
  wire[5:0] idxPagesOH_0;
  wire[7:0] T177;
  wire[2:0] T178;
  reg [2:0] idxPages [61:0];
  wire[2:0] T179;
  wire[2:0] T1606;
  wire[1:0] T1607;
  wire T1608;
  wire[1:0] T1609;
  wire[1:0] T1610;
  wire[3:0] T1611;
  wire[3:0] T1612;
  wire[3:0] T1613;
  wire[1:0] T1614;
  wire T1615;
  wire T1616;
  wire T180;
  wire T181;
  wire T182;
  wire[5:0] T183;
  wire[5:0] idxPagesOH_1;
  wire[7:0] T184;
  wire[2:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[5:0] T188;
  wire[5:0] idxPagesOH_2;
  wire[7:0] T189;
  wire[2:0] T190;
  wire T191;
  wire[5:0] T192;
  wire[5:0] idxPagesOH_3;
  wire[7:0] T193;
  wire[2:0] T194;
  wire[3:0] T195;
  wire[1:0] T196;
  wire T197;
  wire[5:0] T198;
  wire[5:0] idxPagesOH_4;
  wire[7:0] T199;
  wire[2:0] T200;
  wire T201;
  wire[5:0] T202;
  wire[5:0] idxPagesOH_5;
  wire[7:0] T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[5:0] T207;
  wire[5:0] idxPagesOH_6;
  wire[7:0] T208;
  wire[2:0] T209;
  wire T210;
  wire[5:0] T211;
  wire[5:0] idxPagesOH_7;
  wire[7:0] T212;
  wire[2:0] T213;
  wire[7:0] T214;
  wire[3:0] T215;
  wire[1:0] T216;
  wire T217;
  wire[5:0] T218;
  wire[5:0] idxPagesOH_8;
  wire[7:0] T219;
  wire[2:0] T220;
  wire T221;
  wire[5:0] T222;
  wire[5:0] idxPagesOH_9;
  wire[7:0] T223;
  wire[2:0] T224;
  wire[1:0] T225;
  wire T226;
  wire[5:0] T227;
  wire[5:0] idxPagesOH_10;
  wire[7:0] T228;
  wire[2:0] T229;
  wire T230;
  wire[5:0] T231;
  wire[5:0] idxPagesOH_11;
  wire[7:0] T232;
  wire[2:0] T233;
  wire[3:0] T234;
  wire[1:0] T235;
  wire T236;
  wire[5:0] T237;
  wire[5:0] idxPagesOH_12;
  wire[7:0] T238;
  wire[2:0] T239;
  wire T240;
  wire[5:0] T241;
  wire[5:0] idxPagesOH_13;
  wire[7:0] T242;
  wire[2:0] T243;
  wire[1:0] T244;
  wire T245;
  wire[5:0] T246;
  wire[5:0] idxPagesOH_14;
  wire[7:0] T247;
  wire[2:0] T248;
  wire T249;
  wire[5:0] T250;
  wire[5:0] idxPagesOH_15;
  wire[7:0] T251;
  wire[2:0] T252;
  wire[14:0] T253;
  wire[7:0] T254;
  wire[3:0] T255;
  wire[1:0] T256;
  wire T257;
  wire[5:0] T258;
  wire[5:0] idxPagesOH_16;
  wire[7:0] T259;
  wire[2:0] T260;
  wire T261;
  wire[5:0] T262;
  wire[5:0] idxPagesOH_17;
  wire[7:0] T263;
  wire[2:0] T264;
  wire[1:0] T265;
  wire T266;
  wire[5:0] T267;
  wire[5:0] idxPagesOH_18;
  wire[7:0] T268;
  wire[2:0] T269;
  wire T270;
  wire[5:0] T271;
  wire[5:0] idxPagesOH_19;
  wire[7:0] T272;
  wire[2:0] T273;
  wire[3:0] T274;
  wire[1:0] T275;
  wire T276;
  wire[5:0] T277;
  wire[5:0] idxPagesOH_20;
  wire[7:0] T278;
  wire[2:0] T279;
  wire T280;
  wire[5:0] T281;
  wire[5:0] idxPagesOH_21;
  wire[7:0] T282;
  wire[2:0] T283;
  wire[1:0] T284;
  wire T285;
  wire[5:0] T286;
  wire[5:0] idxPagesOH_22;
  wire[7:0] T287;
  wire[2:0] T288;
  wire T289;
  wire[5:0] T290;
  wire[5:0] idxPagesOH_23;
  wire[7:0] T291;
  wire[2:0] T292;
  wire[6:0] T293;
  wire[3:0] T294;
  wire[1:0] T295;
  wire T296;
  wire[5:0] T297;
  wire[5:0] idxPagesOH_24;
  wire[7:0] T298;
  wire[2:0] T299;
  wire T300;
  wire[5:0] T301;
  wire[5:0] idxPagesOH_25;
  wire[7:0] T302;
  wire[2:0] T303;
  wire[1:0] T304;
  wire T305;
  wire[5:0] T306;
  wire[5:0] idxPagesOH_26;
  wire[7:0] T307;
  wire[2:0] T308;
  wire T309;
  wire[5:0] T310;
  wire[5:0] idxPagesOH_27;
  wire[7:0] T311;
  wire[2:0] T312;
  wire[2:0] T313;
  wire[1:0] T314;
  wire T315;
  wire[5:0] T316;
  wire[5:0] idxPagesOH_28;
  wire[7:0] T317;
  wire[2:0] T318;
  wire T319;
  wire[5:0] T320;
  wire[5:0] idxPagesOH_29;
  wire[7:0] T321;
  wire[2:0] T322;
  wire T323;
  wire[5:0] T324;
  wire[5:0] idxPagesOH_30;
  wire[7:0] T325;
  wire[2:0] T326;
  wire[30:0] T327;
  wire[15:0] T328;
  wire[7:0] T329;
  wire[3:0] T330;
  wire[1:0] T331;
  wire T332;
  wire[5:0] T333;
  wire[5:0] idxPagesOH_31;
  wire[7:0] T334;
  wire[2:0] T335;
  wire T336;
  wire[5:0] T337;
  wire[5:0] idxPagesOH_32;
  wire[7:0] T338;
  wire[2:0] T339;
  wire[1:0] T340;
  wire T341;
  wire[5:0] T342;
  wire[5:0] idxPagesOH_33;
  wire[7:0] T343;
  wire[2:0] T344;
  wire T345;
  wire[5:0] T346;
  wire[5:0] idxPagesOH_34;
  wire[7:0] T347;
  wire[2:0] T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire T351;
  wire[5:0] T352;
  wire[5:0] idxPagesOH_35;
  wire[7:0] T353;
  wire[2:0] T354;
  wire T355;
  wire[5:0] T356;
  wire[5:0] idxPagesOH_36;
  wire[7:0] T357;
  wire[2:0] T358;
  wire[1:0] T359;
  wire T360;
  wire[5:0] T361;
  wire[5:0] idxPagesOH_37;
  wire[7:0] T362;
  wire[2:0] T363;
  wire T364;
  wire[5:0] T365;
  wire[5:0] idxPagesOH_38;
  wire[7:0] T366;
  wire[2:0] T367;
  wire[7:0] T368;
  wire[3:0] T369;
  wire[1:0] T370;
  wire T371;
  wire[5:0] T372;
  wire[5:0] idxPagesOH_39;
  wire[7:0] T373;
  wire[2:0] T374;
  wire T375;
  wire[5:0] T376;
  wire[5:0] idxPagesOH_40;
  wire[7:0] T377;
  wire[2:0] T378;
  wire[1:0] T379;
  wire T380;
  wire[5:0] T381;
  wire[5:0] idxPagesOH_41;
  wire[7:0] T382;
  wire[2:0] T383;
  wire T384;
  wire[5:0] T385;
  wire[5:0] idxPagesOH_42;
  wire[7:0] T386;
  wire[2:0] T387;
  wire[3:0] T388;
  wire[1:0] T389;
  wire T390;
  wire[5:0] T391;
  wire[5:0] idxPagesOH_43;
  wire[7:0] T392;
  wire[2:0] T393;
  wire T394;
  wire[5:0] T395;
  wire[5:0] idxPagesOH_44;
  wire[7:0] T396;
  wire[2:0] T397;
  wire[1:0] T398;
  wire T399;
  wire[5:0] T400;
  wire[5:0] idxPagesOH_45;
  wire[7:0] T401;
  wire[2:0] T402;
  wire T403;
  wire[5:0] T404;
  wire[5:0] idxPagesOH_46;
  wire[7:0] T405;
  wire[2:0] T406;
  wire[14:0] T407;
  wire[7:0] T408;
  wire[3:0] T409;
  wire[1:0] T410;
  wire T411;
  wire[5:0] T412;
  wire[5:0] idxPagesOH_47;
  wire[7:0] T413;
  wire[2:0] T414;
  wire T415;
  wire[5:0] T416;
  wire[5:0] idxPagesOH_48;
  wire[7:0] T417;
  wire[2:0] T418;
  wire[1:0] T419;
  wire T420;
  wire[5:0] T421;
  wire[5:0] idxPagesOH_49;
  wire[7:0] T422;
  wire[2:0] T423;
  wire T424;
  wire[5:0] T425;
  wire[5:0] idxPagesOH_50;
  wire[7:0] T426;
  wire[2:0] T427;
  wire[3:0] T428;
  wire[1:0] T429;
  wire T430;
  wire[5:0] T431;
  wire[5:0] idxPagesOH_51;
  wire[7:0] T432;
  wire[2:0] T433;
  wire T434;
  wire[5:0] T435;
  wire[5:0] idxPagesOH_52;
  wire[7:0] T436;
  wire[2:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[5:0] T440;
  wire[5:0] idxPagesOH_53;
  wire[7:0] T441;
  wire[2:0] T442;
  wire T443;
  wire[5:0] T444;
  wire[5:0] idxPagesOH_54;
  wire[7:0] T445;
  wire[2:0] T446;
  wire[6:0] T447;
  wire[3:0] T448;
  wire[1:0] T449;
  wire T450;
  wire[5:0] T451;
  wire[5:0] idxPagesOH_55;
  wire[7:0] T452;
  wire[2:0] T453;
  wire T454;
  wire[5:0] T455;
  wire[5:0] idxPagesOH_56;
  wire[7:0] T456;
  wire[2:0] T457;
  wire[1:0] T458;
  wire T459;
  wire[5:0] T460;
  wire[5:0] idxPagesOH_57;
  wire[7:0] T461;
  wire[2:0] T462;
  wire T463;
  wire[5:0] T464;
  wire[5:0] idxPagesOH_58;
  wire[7:0] T465;
  wire[2:0] T466;
  wire[2:0] T467;
  wire[1:0] T468;
  wire T469;
  wire[5:0] T470;
  wire[5:0] idxPagesOH_59;
  wire[7:0] T471;
  wire[2:0] T472;
  wire T473;
  wire[5:0] T474;
  wire[5:0] idxPagesOH_60;
  wire[7:0] T475;
  wire[2:0] T476;
  wire T477;
  wire[5:0] T478;
  wire[5:0] idxPagesOH_61;
  wire[7:0] T479;
  wire[2:0] T480;
  wire[61:0] T481;
  wire[61:0] T482;
  wire[61:0] T483;
  wire[30:0] T484;
  wire[15:0] T485;
  wire[7:0] T486;
  wire[3:0] T487;
  wire[1:0] T488;
  wire T489;
  wire[12:0] T490;
  wire[12:0] T491;
  reg [12:0] idxs [61:0];
  wire[12:0] T492;
  wire[12:0] T1617;
  wire T493;
  wire T494;
  wire T495;
  wire[12:0] T496;
  wire[1:0] T497;
  wire T498;
  wire[12:0] T499;
  wire T500;
  wire[12:0] T501;
  wire[3:0] T502;
  wire[1:0] T503;
  wire T504;
  wire[12:0] T505;
  wire T506;
  wire[12:0] T507;
  wire[1:0] T508;
  wire T509;
  wire[12:0] T510;
  wire T511;
  wire[12:0] T512;
  wire[7:0] T513;
  wire[3:0] T514;
  wire[1:0] T515;
  wire T516;
  wire[12:0] T517;
  wire T518;
  wire[12:0] T519;
  wire[1:0] T520;
  wire T521;
  wire[12:0] T522;
  wire T523;
  wire[12:0] T524;
  wire[3:0] T525;
  wire[1:0] T526;
  wire T527;
  wire[12:0] T528;
  wire T529;
  wire[12:0] T530;
  wire[1:0] T531;
  wire T532;
  wire[12:0] T533;
  wire T534;
  wire[12:0] T535;
  wire[14:0] T536;
  wire[7:0] T537;
  wire[3:0] T538;
  wire[1:0] T539;
  wire T540;
  wire[12:0] T541;
  wire T542;
  wire[12:0] T543;
  wire[1:0] T544;
  wire T545;
  wire[12:0] T546;
  wire T547;
  wire[12:0] T548;
  wire[3:0] T549;
  wire[1:0] T550;
  wire T551;
  wire[12:0] T552;
  wire T553;
  wire[12:0] T554;
  wire[1:0] T555;
  wire T556;
  wire[12:0] T557;
  wire T558;
  wire[12:0] T559;
  wire[6:0] T560;
  wire[3:0] T561;
  wire[1:0] T562;
  wire T563;
  wire[12:0] T564;
  wire T565;
  wire[12:0] T566;
  wire[1:0] T567;
  wire T568;
  wire[12:0] T569;
  wire T570;
  wire[12:0] T571;
  wire[2:0] T572;
  wire[1:0] T573;
  wire T574;
  wire[12:0] T575;
  wire T576;
  wire[12:0] T577;
  wire T578;
  wire[12:0] T579;
  wire[30:0] T580;
  wire[15:0] T581;
  wire[7:0] T582;
  wire[3:0] T583;
  wire[1:0] T584;
  wire T585;
  wire[12:0] T586;
  wire T587;
  wire[12:0] T588;
  wire[1:0] T589;
  wire T590;
  wire[12:0] T591;
  wire T592;
  wire[12:0] T593;
  wire[3:0] T594;
  wire[1:0] T595;
  wire T596;
  wire[12:0] T597;
  wire T598;
  wire[12:0] T599;
  wire[1:0] T600;
  wire T601;
  wire[12:0] T602;
  wire T603;
  wire[12:0] T604;
  wire[7:0] T605;
  wire[3:0] T606;
  wire[1:0] T607;
  wire T608;
  wire[12:0] T609;
  wire T610;
  wire[12:0] T611;
  wire[1:0] T612;
  wire T613;
  wire[12:0] T614;
  wire T615;
  wire[12:0] T616;
  wire[3:0] T617;
  wire[1:0] T618;
  wire T619;
  wire[12:0] T620;
  wire T621;
  wire[12:0] T622;
  wire[1:0] T623;
  wire T624;
  wire[12:0] T625;
  wire T626;
  wire[12:0] T627;
  wire[14:0] T628;
  wire[7:0] T629;
  wire[3:0] T630;
  wire[1:0] T631;
  wire T632;
  wire[12:0] T633;
  wire T634;
  wire[12:0] T635;
  wire[1:0] T636;
  wire T637;
  wire[12:0] T638;
  wire T639;
  wire[12:0] T640;
  wire[3:0] T641;
  wire[1:0] T642;
  wire T643;
  wire[12:0] T644;
  wire T645;
  wire[12:0] T646;
  wire[1:0] T647;
  wire T648;
  wire[12:0] T649;
  wire T650;
  wire[12:0] T651;
  wire[6:0] T652;
  wire[3:0] T653;
  wire[1:0] T654;
  wire T655;
  wire[12:0] T656;
  wire T657;
  wire[12:0] T658;
  wire[1:0] T659;
  wire T660;
  wire[12:0] T661;
  wire T662;
  wire[12:0] T663;
  wire[2:0] T664;
  wire[1:0] T665;
  wire T666;
  wire[12:0] T667;
  wire T668;
  wire[12:0] T669;
  wire T670;
  wire[12:0] T671;
  reg [61:0] idxValid;
  wire[61:0] T1618;
  wire[63:0] T1619;
  wire[63:0] T672;
  wire[63:0] T673;
  wire[63:0] T1620;
  wire[61:0] T674;
  wire[61:0] T675;
  wire[61:0] T676;
  wire[61:0] T677;
  wire[61:0] T678;
  wire[30:0] T679;
  wire[15:0] T680;
  wire[7:0] T681;
  wire[3:0] T682;
  wire[1:0] T683;
  wire T684;
  wire[7:0] T685;
  wire[7:0] T1621;
  wire[5:0] T686;
  wire[5:0] tgtPagesOH_0;
  wire[7:0] T687;
  wire[2:0] T688;
  reg [2:0] tgtPages [61:0];
  wire[2:0] T689;
  wire[2:0] T1622;
  wire[1:0] T1623;
  wire T1624;
  wire[1:0] T1625;
  wire[1:0] T1626;
  wire[3:0] T1627;
  wire[3:0] T1628;
  wire[7:0] T690;
  wire[7:0] T1629;
  wire[3:0] T1630;
  wire[1:0] T1631;
  wire T1632;
  wire T1633;
  wire T691;
  wire T692;
  wire T693;
  wire[7:0] T694;
  wire[7:0] T1634;
  wire[5:0] T695;
  wire[5:0] tgtPagesOH_1;
  wire[7:0] T696;
  wire[2:0] T697;
  wire[1:0] T698;
  wire T699;
  wire[7:0] T700;
  wire[7:0] T1635;
  wire[5:0] T701;
  wire[5:0] tgtPagesOH_2;
  wire[7:0] T702;
  wire[2:0] T703;
  wire T704;
  wire[7:0] T705;
  wire[7:0] T1636;
  wire[5:0] T706;
  wire[5:0] tgtPagesOH_3;
  wire[7:0] T707;
  wire[2:0] T708;
  wire[3:0] T709;
  wire[1:0] T710;
  wire T711;
  wire[7:0] T712;
  wire[7:0] T1637;
  wire[5:0] T713;
  wire[5:0] tgtPagesOH_4;
  wire[7:0] T714;
  wire[2:0] T715;
  wire T716;
  wire[7:0] T717;
  wire[7:0] T1638;
  wire[5:0] T718;
  wire[5:0] tgtPagesOH_5;
  wire[7:0] T719;
  wire[2:0] T720;
  wire[1:0] T721;
  wire T722;
  wire[7:0] T723;
  wire[7:0] T1639;
  wire[5:0] T724;
  wire[5:0] tgtPagesOH_6;
  wire[7:0] T725;
  wire[2:0] T726;
  wire T727;
  wire[7:0] T728;
  wire[7:0] T1640;
  wire[5:0] T729;
  wire[5:0] tgtPagesOH_7;
  wire[7:0] T730;
  wire[2:0] T731;
  wire[7:0] T732;
  wire[3:0] T733;
  wire[1:0] T734;
  wire T735;
  wire[7:0] T736;
  wire[7:0] T1641;
  wire[5:0] T737;
  wire[5:0] tgtPagesOH_8;
  wire[7:0] T738;
  wire[2:0] T739;
  wire T740;
  wire[7:0] T741;
  wire[7:0] T1642;
  wire[5:0] T742;
  wire[5:0] tgtPagesOH_9;
  wire[7:0] T743;
  wire[2:0] T744;
  wire[1:0] T745;
  wire T746;
  wire[7:0] T747;
  wire[7:0] T1643;
  wire[5:0] T748;
  wire[5:0] tgtPagesOH_10;
  wire[7:0] T749;
  wire[2:0] T750;
  wire T751;
  wire[7:0] T752;
  wire[7:0] T1644;
  wire[5:0] T753;
  wire[5:0] tgtPagesOH_11;
  wire[7:0] T754;
  wire[2:0] T755;
  wire[3:0] T756;
  wire[1:0] T757;
  wire T758;
  wire[7:0] T759;
  wire[7:0] T1645;
  wire[5:0] T760;
  wire[5:0] tgtPagesOH_12;
  wire[7:0] T761;
  wire[2:0] T762;
  wire T763;
  wire[7:0] T764;
  wire[7:0] T1646;
  wire[5:0] T765;
  wire[5:0] tgtPagesOH_13;
  wire[7:0] T766;
  wire[2:0] T767;
  wire[1:0] T768;
  wire T769;
  wire[7:0] T770;
  wire[7:0] T1647;
  wire[5:0] T771;
  wire[5:0] tgtPagesOH_14;
  wire[7:0] T772;
  wire[2:0] T773;
  wire T774;
  wire[7:0] T775;
  wire[7:0] T1648;
  wire[5:0] T776;
  wire[5:0] tgtPagesOH_15;
  wire[7:0] T777;
  wire[2:0] T778;
  wire[14:0] T779;
  wire[7:0] T780;
  wire[3:0] T781;
  wire[1:0] T782;
  wire T783;
  wire[7:0] T784;
  wire[7:0] T1649;
  wire[5:0] T785;
  wire[5:0] tgtPagesOH_16;
  wire[7:0] T786;
  wire[2:0] T787;
  wire T788;
  wire[7:0] T789;
  wire[7:0] T1650;
  wire[5:0] T790;
  wire[5:0] tgtPagesOH_17;
  wire[7:0] T791;
  wire[2:0] T792;
  wire[1:0] T793;
  wire T794;
  wire[7:0] T795;
  wire[7:0] T1651;
  wire[5:0] T796;
  wire[5:0] tgtPagesOH_18;
  wire[7:0] T797;
  wire[2:0] T798;
  wire T799;
  wire[7:0] T800;
  wire[7:0] T1652;
  wire[5:0] T801;
  wire[5:0] tgtPagesOH_19;
  wire[7:0] T802;
  wire[2:0] T803;
  wire[3:0] T804;
  wire[1:0] T805;
  wire T806;
  wire[7:0] T807;
  wire[7:0] T1653;
  wire[5:0] T808;
  wire[5:0] tgtPagesOH_20;
  wire[7:0] T809;
  wire[2:0] T810;
  wire T811;
  wire[7:0] T812;
  wire[7:0] T1654;
  wire[5:0] T813;
  wire[5:0] tgtPagesOH_21;
  wire[7:0] T814;
  wire[2:0] T815;
  wire[1:0] T816;
  wire T817;
  wire[7:0] T818;
  wire[7:0] T1655;
  wire[5:0] T819;
  wire[5:0] tgtPagesOH_22;
  wire[7:0] T820;
  wire[2:0] T821;
  wire T822;
  wire[7:0] T823;
  wire[7:0] T1656;
  wire[5:0] T824;
  wire[5:0] tgtPagesOH_23;
  wire[7:0] T825;
  wire[2:0] T826;
  wire[6:0] T827;
  wire[3:0] T828;
  wire[1:0] T829;
  wire T830;
  wire[7:0] T831;
  wire[7:0] T1657;
  wire[5:0] T832;
  wire[5:0] tgtPagesOH_24;
  wire[7:0] T833;
  wire[2:0] T834;
  wire T835;
  wire[7:0] T836;
  wire[7:0] T1658;
  wire[5:0] T837;
  wire[5:0] tgtPagesOH_25;
  wire[7:0] T838;
  wire[2:0] T839;
  wire[1:0] T840;
  wire T841;
  wire[7:0] T842;
  wire[7:0] T1659;
  wire[5:0] T843;
  wire[5:0] tgtPagesOH_26;
  wire[7:0] T844;
  wire[2:0] T845;
  wire T846;
  wire[7:0] T847;
  wire[7:0] T1660;
  wire[5:0] T848;
  wire[5:0] tgtPagesOH_27;
  wire[7:0] T849;
  wire[2:0] T850;
  wire[2:0] T851;
  wire[1:0] T852;
  wire T853;
  wire[7:0] T854;
  wire[7:0] T1661;
  wire[5:0] T855;
  wire[5:0] tgtPagesOH_28;
  wire[7:0] T856;
  wire[2:0] T857;
  wire T858;
  wire[7:0] T859;
  wire[7:0] T1662;
  wire[5:0] T860;
  wire[5:0] tgtPagesOH_29;
  wire[7:0] T861;
  wire[2:0] T862;
  wire T863;
  wire[7:0] T864;
  wire[7:0] T1663;
  wire[5:0] T865;
  wire[5:0] tgtPagesOH_30;
  wire[7:0] T866;
  wire[2:0] T867;
  wire[30:0] T868;
  wire[15:0] T869;
  wire[7:0] T870;
  wire[3:0] T871;
  wire[1:0] T872;
  wire T873;
  wire[7:0] T874;
  wire[7:0] T1664;
  wire[5:0] T875;
  wire[5:0] tgtPagesOH_31;
  wire[7:0] T876;
  wire[2:0] T877;
  wire T878;
  wire[7:0] T879;
  wire[7:0] T1665;
  wire[5:0] T880;
  wire[5:0] tgtPagesOH_32;
  wire[7:0] T881;
  wire[2:0] T882;
  wire[1:0] T883;
  wire T884;
  wire[7:0] T885;
  wire[7:0] T1666;
  wire[5:0] T886;
  wire[5:0] tgtPagesOH_33;
  wire[7:0] T887;
  wire[2:0] T888;
  wire T889;
  wire[7:0] T890;
  wire[7:0] T1667;
  wire[5:0] T891;
  wire[5:0] tgtPagesOH_34;
  wire[7:0] T892;
  wire[2:0] T893;
  wire[3:0] T894;
  wire[1:0] T895;
  wire T896;
  wire[7:0] T897;
  wire[7:0] T1668;
  wire[5:0] T898;
  wire[5:0] tgtPagesOH_35;
  wire[7:0] T899;
  wire[2:0] T900;
  wire T901;
  wire[7:0] T902;
  wire[7:0] T1669;
  wire[5:0] T903;
  wire[5:0] tgtPagesOH_36;
  wire[7:0] T904;
  wire[2:0] T905;
  wire[1:0] T906;
  wire T907;
  wire[7:0] T908;
  wire[7:0] T1670;
  wire[5:0] T909;
  wire[5:0] tgtPagesOH_37;
  wire[7:0] T910;
  wire[2:0] T911;
  wire T912;
  wire[7:0] T913;
  wire[7:0] T1671;
  wire[5:0] T914;
  wire[5:0] tgtPagesOH_38;
  wire[7:0] T915;
  wire[2:0] T916;
  wire[7:0] T917;
  wire[3:0] T918;
  wire[1:0] T919;
  wire T920;
  wire[7:0] T921;
  wire[7:0] T1672;
  wire[5:0] T922;
  wire[5:0] tgtPagesOH_39;
  wire[7:0] T923;
  wire[2:0] T924;
  wire T925;
  wire[7:0] T926;
  wire[7:0] T1673;
  wire[5:0] T927;
  wire[5:0] tgtPagesOH_40;
  wire[7:0] T928;
  wire[2:0] T929;
  wire[1:0] T930;
  wire T931;
  wire[7:0] T932;
  wire[7:0] T1674;
  wire[5:0] T933;
  wire[5:0] tgtPagesOH_41;
  wire[7:0] T934;
  wire[2:0] T935;
  wire T936;
  wire[7:0] T937;
  wire[7:0] T1675;
  wire[5:0] T938;
  wire[5:0] tgtPagesOH_42;
  wire[7:0] T939;
  wire[2:0] T940;
  wire[3:0] T941;
  wire[1:0] T942;
  wire T943;
  wire[7:0] T944;
  wire[7:0] T1676;
  wire[5:0] T945;
  wire[5:0] tgtPagesOH_43;
  wire[7:0] T946;
  wire[2:0] T947;
  wire T948;
  wire[7:0] T949;
  wire[7:0] T1677;
  wire[5:0] T950;
  wire[5:0] tgtPagesOH_44;
  wire[7:0] T951;
  wire[2:0] T952;
  wire[1:0] T953;
  wire T954;
  wire[7:0] T955;
  wire[7:0] T1678;
  wire[5:0] T956;
  wire[5:0] tgtPagesOH_45;
  wire[7:0] T957;
  wire[2:0] T958;
  wire T959;
  wire[7:0] T960;
  wire[7:0] T1679;
  wire[5:0] T961;
  wire[5:0] tgtPagesOH_46;
  wire[7:0] T962;
  wire[2:0] T963;
  wire[14:0] T964;
  wire[7:0] T965;
  wire[3:0] T966;
  wire[1:0] T967;
  wire T968;
  wire[7:0] T969;
  wire[7:0] T1680;
  wire[5:0] T970;
  wire[5:0] tgtPagesOH_47;
  wire[7:0] T971;
  wire[2:0] T972;
  wire T973;
  wire[7:0] T974;
  wire[7:0] T1681;
  wire[5:0] T975;
  wire[5:0] tgtPagesOH_48;
  wire[7:0] T976;
  wire[2:0] T977;
  wire[1:0] T978;
  wire T979;
  wire[7:0] T980;
  wire[7:0] T1682;
  wire[5:0] T981;
  wire[5:0] tgtPagesOH_49;
  wire[7:0] T982;
  wire[2:0] T983;
  wire T984;
  wire[7:0] T985;
  wire[7:0] T1683;
  wire[5:0] T986;
  wire[5:0] tgtPagesOH_50;
  wire[7:0] T987;
  wire[2:0] T988;
  wire[3:0] T989;
  wire[1:0] T990;
  wire T991;
  wire[7:0] T992;
  wire[7:0] T1684;
  wire[5:0] T993;
  wire[5:0] tgtPagesOH_51;
  wire[7:0] T994;
  wire[2:0] T995;
  wire T996;
  wire[7:0] T997;
  wire[7:0] T1685;
  wire[5:0] T998;
  wire[5:0] tgtPagesOH_52;
  wire[7:0] T999;
  wire[2:0] T1000;
  wire[1:0] T1001;
  wire T1002;
  wire[7:0] T1003;
  wire[7:0] T1686;
  wire[5:0] T1004;
  wire[5:0] tgtPagesOH_53;
  wire[7:0] T1005;
  wire[2:0] T1006;
  wire T1007;
  wire[7:0] T1008;
  wire[7:0] T1687;
  wire[5:0] T1009;
  wire[5:0] tgtPagesOH_54;
  wire[7:0] T1010;
  wire[2:0] T1011;
  wire[6:0] T1012;
  wire[3:0] T1013;
  wire[1:0] T1014;
  wire T1015;
  wire[7:0] T1016;
  wire[7:0] T1688;
  wire[5:0] T1017;
  wire[5:0] tgtPagesOH_55;
  wire[7:0] T1018;
  wire[2:0] T1019;
  wire T1020;
  wire[7:0] T1021;
  wire[7:0] T1689;
  wire[5:0] T1022;
  wire[5:0] tgtPagesOH_56;
  wire[7:0] T1023;
  wire[2:0] T1024;
  wire[1:0] T1025;
  wire T1026;
  wire[7:0] T1027;
  wire[7:0] T1690;
  wire[5:0] T1028;
  wire[5:0] tgtPagesOH_57;
  wire[7:0] T1029;
  wire[2:0] T1030;
  wire T1031;
  wire[7:0] T1032;
  wire[7:0] T1691;
  wire[5:0] T1033;
  wire[5:0] tgtPagesOH_58;
  wire[7:0] T1034;
  wire[2:0] T1035;
  wire[2:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire[7:0] T1039;
  wire[7:0] T1692;
  wire[5:0] T1040;
  wire[5:0] tgtPagesOH_59;
  wire[7:0] T1041;
  wire[2:0] T1042;
  wire T1043;
  wire[7:0] T1044;
  wire[7:0] T1693;
  wire[5:0] T1045;
  wire[5:0] tgtPagesOH_60;
  wire[7:0] T1046;
  wire[2:0] T1047;
  wire T1048;
  wire[7:0] T1049;
  wire[7:0] T1694;
  wire[5:0] T1050;
  wire[5:0] tgtPagesOH_61;
  wire[7:0] T1051;
  wire[2:0] T1052;
  wire[63:0] T1053;
  wire[63:0] T1054;
  wire[63:0] T1055;
  wire[63:0] T1695;
  wire[61:0] T1056;
  wire[63:0] T1057;
  wire[63:0] T1696;
  wire T1058;
  wire T1059;
  wire[63:0] T1060;
  wire[63:0] T1061;
  wire[63:0] T1697;
  wire T1062;
  wire T1063;
  wire[6:0] T1064;
  wire[5:0] T1065;
  wire T1066;
  wire[6:0] T1067;
  wire[6:0] T1068;
  wire[5:0] T1698;
  wire[4:0] T1699;
  wire[3:0] T1700;
  wire[2:0] T1701;
  wire[1:0] T1702;
  wire T1703;
  wire[1:0] T1704;
  wire[1:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[7:0] T1708;
  wire[7:0] T1709;
  wire[15:0] T1710;
  wire[15:0] T1711;
  wire[31:0] T1712;
  wire[31:0] T1713;
  wire[29:0] T1714;
  wire[15:0] T1715;
  wire[7:0] T1716;
  wire[3:0] T1717;
  wire[1:0] T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire T1723;
  wire[42:0] T1070;
  wire[42:0] T1071;
  wire[42:0] T1072;
  wire[12:0] T1073;
  wire[12:0] T1074;
  wire[12:0] T1075;
  reg [12:0] tgts [61:0];
  wire[12:0] T1076;
  wire[12:0] T1724;
  wire T1077;
  wire T1078;
  wire T1079;
  wire[12:0] T1080;
  wire[12:0] T1081;
  wire[12:0] T1082;
  wire T1083;
  wire[12:0] T1084;
  wire[12:0] T1085;
  wire[12:0] T1086;
  wire T1087;
  wire[12:0] T1088;
  wire[12:0] T1089;
  wire[12:0] T1090;
  wire T1091;
  wire[12:0] T1092;
  wire[12:0] T1093;
  wire[12:0] T1094;
  wire T1095;
  wire[12:0] T1096;
  wire[12:0] T1097;
  wire[12:0] T1098;
  wire T1099;
  wire[12:0] T1100;
  wire[12:0] T1101;
  wire[12:0] T1102;
  wire T1103;
  wire[12:0] T1104;
  wire[12:0] T1105;
  wire[12:0] T1106;
  wire T1107;
  wire[12:0] T1108;
  wire[12:0] T1109;
  wire[12:0] T1110;
  wire T1111;
  wire[12:0] T1112;
  wire[12:0] T1113;
  wire[12:0] T1114;
  wire T1115;
  wire[12:0] T1116;
  wire[12:0] T1117;
  wire[12:0] T1118;
  wire T1119;
  wire[12:0] T1120;
  wire[12:0] T1121;
  wire[12:0] T1122;
  wire T1123;
  wire[12:0] T1124;
  wire[12:0] T1125;
  wire[12:0] T1126;
  wire T1127;
  wire[12:0] T1128;
  wire[12:0] T1129;
  wire[12:0] T1130;
  wire T1131;
  wire[12:0] T1132;
  wire[12:0] T1133;
  wire[12:0] T1134;
  wire T1135;
  wire[12:0] T1136;
  wire[12:0] T1137;
  wire[12:0] T1138;
  wire T1139;
  wire[12:0] T1140;
  wire[12:0] T1141;
  wire[12:0] T1142;
  wire T1143;
  wire[12:0] T1144;
  wire[12:0] T1145;
  wire[12:0] T1146;
  wire T1147;
  wire[12:0] T1148;
  wire[12:0] T1149;
  wire[12:0] T1150;
  wire T1151;
  wire[12:0] T1152;
  wire[12:0] T1153;
  wire[12:0] T1154;
  wire T1155;
  wire[12:0] T1156;
  wire[12:0] T1157;
  wire[12:0] T1158;
  wire T1159;
  wire[12:0] T1160;
  wire[12:0] T1161;
  wire[12:0] T1162;
  wire T1163;
  wire[12:0] T1164;
  wire[12:0] T1165;
  wire[12:0] T1166;
  wire T1167;
  wire[12:0] T1168;
  wire[12:0] T1169;
  wire[12:0] T1170;
  wire T1171;
  wire[12:0] T1172;
  wire[12:0] T1173;
  wire[12:0] T1174;
  wire T1175;
  wire[12:0] T1176;
  wire[12:0] T1177;
  wire[12:0] T1178;
  wire T1179;
  wire[12:0] T1180;
  wire[12:0] T1181;
  wire[12:0] T1182;
  wire T1183;
  wire[12:0] T1184;
  wire[12:0] T1185;
  wire[12:0] T1186;
  wire T1187;
  wire[12:0] T1188;
  wire[12:0] T1189;
  wire[12:0] T1190;
  wire T1191;
  wire[12:0] T1192;
  wire[12:0] T1193;
  wire[12:0] T1194;
  wire T1195;
  wire[12:0] T1196;
  wire[12:0] T1197;
  wire[12:0] T1198;
  wire T1199;
  wire[12:0] T1200;
  wire[12:0] T1201;
  wire[12:0] T1202;
  wire T1203;
  wire[12:0] T1204;
  wire[12:0] T1205;
  wire[12:0] T1206;
  wire T1207;
  wire[12:0] T1208;
  wire[12:0] T1209;
  wire[12:0] T1210;
  wire T1211;
  wire[12:0] T1212;
  wire[12:0] T1213;
  wire[12:0] T1214;
  wire T1215;
  wire[12:0] T1216;
  wire[12:0] T1217;
  wire[12:0] T1218;
  wire T1219;
  wire[12:0] T1220;
  wire[12:0] T1221;
  wire[12:0] T1222;
  wire T1223;
  wire[12:0] T1224;
  wire[12:0] T1225;
  wire[12:0] T1226;
  wire T1227;
  wire[12:0] T1228;
  wire[12:0] T1229;
  wire[12:0] T1230;
  wire T1231;
  wire[12:0] T1232;
  wire[12:0] T1233;
  wire[12:0] T1234;
  wire T1235;
  wire[12:0] T1236;
  wire[12:0] T1237;
  wire[12:0] T1238;
  wire T1239;
  wire[12:0] T1240;
  wire[12:0] T1241;
  wire[12:0] T1242;
  wire T1243;
  wire[12:0] T1244;
  wire[12:0] T1245;
  wire[12:0] T1246;
  wire T1247;
  wire[12:0] T1248;
  wire[12:0] T1249;
  wire[12:0] T1250;
  wire T1251;
  wire[12:0] T1252;
  wire[12:0] T1253;
  wire[12:0] T1254;
  wire T1255;
  wire[12:0] T1256;
  wire[12:0] T1257;
  wire[12:0] T1258;
  wire T1259;
  wire[12:0] T1260;
  wire[12:0] T1261;
  wire[12:0] T1262;
  wire T1263;
  wire[12:0] T1264;
  wire[12:0] T1265;
  wire[12:0] T1266;
  wire T1267;
  wire[12:0] T1268;
  wire[12:0] T1269;
  wire[12:0] T1270;
  wire T1271;
  wire[12:0] T1272;
  wire[12:0] T1273;
  wire[12:0] T1274;
  wire T1275;
  wire[12:0] T1276;
  wire[12:0] T1277;
  wire[12:0] T1278;
  wire T1279;
  wire[12:0] T1280;
  wire[12:0] T1281;
  wire[12:0] T1282;
  wire T1283;
  wire[12:0] T1284;
  wire[12:0] T1285;
  wire[12:0] T1286;
  wire T1287;
  wire[12:0] T1288;
  wire[12:0] T1289;
  wire[12:0] T1290;
  wire T1291;
  wire[12:0] T1292;
  wire[12:0] T1293;
  wire[12:0] T1294;
  wire T1295;
  wire[12:0] T1296;
  wire[12:0] T1297;
  wire[12:0] T1298;
  wire T1299;
  wire[12:0] T1300;
  wire[12:0] T1301;
  wire[12:0] T1302;
  wire T1303;
  wire[12:0] T1304;
  wire[12:0] T1305;
  wire[12:0] T1306;
  wire T1307;
  wire[12:0] T1308;
  wire[12:0] T1309;
  wire[12:0] T1310;
  wire T1311;
  wire[12:0] T1312;
  wire[12:0] T1313;
  wire[12:0] T1314;
  wire T1315;
  wire[12:0] T1316;
  wire[12:0] T1317;
  wire[12:0] T1318;
  wire T1319;
  wire[12:0] T1320;
  wire[12:0] T1321;
  wire T1322;
  wire[29:0] T1323;
  wire[29:0] T1324;
  wire[29:0] T1325;
  wire T1326;
  wire[5:0] T1327;
  wire[5:0] T1328;
  wire T1329;
  wire[5:0] T1330;
  wire[5:0] T1331;
  wire T1332;
  wire[5:0] T1333;
  wire[5:0] T1334;
  wire T1335;
  wire[5:0] T1336;
  wire[5:0] T1337;
  wire T1338;
  wire[5:0] T1339;
  wire[5:0] T1340;
  wire T1341;
  wire[5:0] T1342;
  wire[5:0] T1343;
  wire T1344;
  wire[5:0] T1345;
  wire[5:0] T1346;
  wire T1347;
  wire[5:0] T1348;
  wire[5:0] T1349;
  wire T1350;
  wire[5:0] T1351;
  wire[5:0] T1352;
  wire T1353;
  wire[5:0] T1354;
  wire[5:0] T1355;
  wire T1356;
  wire[5:0] T1357;
  wire[5:0] T1358;
  wire T1359;
  wire[5:0] T1360;
  wire[5:0] T1361;
  wire T1362;
  wire[5:0] T1363;
  wire[5:0] T1364;
  wire T1365;
  wire[5:0] T1366;
  wire[5:0] T1367;
  wire T1368;
  wire[5:0] T1369;
  wire[5:0] T1370;
  wire T1371;
  wire[5:0] T1372;
  wire[5:0] T1373;
  wire T1374;
  wire[5:0] T1375;
  wire[5:0] T1376;
  wire T1377;
  wire[5:0] T1378;
  wire[5:0] T1379;
  wire T1380;
  wire[5:0] T1381;
  wire[5:0] T1382;
  wire T1383;
  wire[5:0] T1384;
  wire[5:0] T1385;
  wire T1386;
  wire[5:0] T1387;
  wire[5:0] T1388;
  wire T1389;
  wire[5:0] T1390;
  wire[5:0] T1391;
  wire T1392;
  wire[5:0] T1393;
  wire[5:0] T1394;
  wire T1395;
  wire[5:0] T1396;
  wire[5:0] T1397;
  wire T1398;
  wire[5:0] T1399;
  wire[5:0] T1400;
  wire T1401;
  wire[5:0] T1402;
  wire[5:0] T1403;
  wire T1404;
  wire[5:0] T1405;
  wire[5:0] T1406;
  wire T1407;
  wire[5:0] T1408;
  wire[5:0] T1409;
  wire T1410;
  wire[5:0] T1411;
  wire[5:0] T1412;
  wire T1413;
  wire[5:0] T1414;
  wire[5:0] T1415;
  wire T1416;
  wire[5:0] T1417;
  wire[5:0] T1418;
  wire T1419;
  wire[5:0] T1420;
  wire[5:0] T1421;
  wire T1422;
  wire[5:0] T1423;
  wire[5:0] T1424;
  wire T1425;
  wire[5:0] T1426;
  wire[5:0] T1427;
  wire T1428;
  wire[5:0] T1429;
  wire[5:0] T1430;
  wire T1431;
  wire[5:0] T1432;
  wire[5:0] T1433;
  wire T1434;
  wire[5:0] T1435;
  wire[5:0] T1436;
  wire T1437;
  wire[5:0] T1438;
  wire[5:0] T1439;
  wire T1440;
  wire[5:0] T1441;
  wire[5:0] T1442;
  wire T1443;
  wire[5:0] T1444;
  wire[5:0] T1445;
  wire T1446;
  wire[5:0] T1447;
  wire[5:0] T1448;
  wire T1449;
  wire[5:0] T1450;
  wire[5:0] T1451;
  wire T1452;
  wire[5:0] T1453;
  wire[5:0] T1454;
  wire T1455;
  wire[5:0] T1456;
  wire[5:0] T1457;
  wire T1458;
  wire[5:0] T1459;
  wire[5:0] T1460;
  wire T1461;
  wire[5:0] T1462;
  wire[5:0] T1463;
  wire T1464;
  wire[5:0] T1465;
  wire[5:0] T1466;
  wire T1467;
  wire[5:0] T1468;
  wire[5:0] T1469;
  wire T1470;
  wire[5:0] T1471;
  wire[5:0] T1472;
  wire T1473;
  wire[5:0] T1474;
  wire[5:0] T1475;
  wire T1476;
  wire[5:0] T1477;
  wire[5:0] T1478;
  wire T1479;
  wire[5:0] T1480;
  wire[5:0] T1481;
  wire T1482;
  wire[5:0] T1483;
  wire[5:0] T1484;
  wire T1485;
  wire[5:0] T1486;
  wire[5:0] T1487;
  wire T1488;
  wire[5:0] T1489;
  wire[5:0] T1490;
  wire T1491;
  wire[5:0] T1492;
  wire[5:0] T1493;
  wire T1494;
  wire[5:0] T1495;
  wire[5:0] T1496;
  wire T1497;
  wire[5:0] T1498;
  wire[5:0] T1499;
  wire T1500;
  wire[5:0] T1501;
  wire[5:0] T1502;
  wire T1503;
  wire[5:0] T1504;
  wire[5:0] T1505;
  wire T1506;
  wire[5:0] T1507;
  wire[5:0] T1508;
  wire T1509;
  wire[5:0] T1510;
  wire T1511;
  wire[29:0] T1512;
  wire[29:0] T1513;
  wire[29:0] T1514;
  wire T1515;
  wire[29:0] T1516;
  wire[29:0] T1517;
  wire[29:0] T1518;
  wire T1519;
  wire[29:0] T1520;
  wire[29:0] T1521;
  wire[29:0] T1522;
  wire T1523;
  wire[29:0] T1524;
  wire[29:0] T1525;
  wire[29:0] T1526;
  wire T1527;
  wire[29:0] T1528;
  wire[29:0] T1529;
  wire T1530;
  wire[42:0] T1531;
  reg [42:0] R1532;
  wire[42:0] T1533;
  wire T1534;
  wire T1535;
  wire[1:0] T1536;
  wire T1537;
  wire T1538;
  reg  R1539;
  wire T1725;
  wire T1540;
  wire T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire T1545;
  reg [1:0] R1546;
  wire[1:0] T1726;
  wire[1:0] T1547;
  wire[1:0] T1548;
  wire[1:0] T1549;
  wire[1:0] T1550;
  wire T1551;
  wire T1552;
  wire[1:0] T1553;
  wire T1554;
  wire T1555;
  wire T1556;
  wire T1557;
  wire T1558;
  reg [42:0] R1559;
  wire[42:0] T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire T1564;
  wire T1565;
  wire[61:0] T1566;
  reg [61:0] useRAS;
  wire[61:0] T1727;
  wire[63:0] T1567;
  wire[63:0] T1728;
  wire[63:0] T1568;
  wire[63:0] T1569;
  wire[63:0] T1570;
  wire[63:0] T1729;
  wire[61:0] T1571;
  wire[63:0] T1572;
  wire[63:0] T1730;
  wire T1573;
  wire T1574;
  reg  R1575;
  wire T1576;
  wire[63:0] T1577;
  wire[63:0] T1578;
  wire[63:0] T1731;
  wire T1579;
  wire T1580;
  wire T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire T1585;
  wire[61:0] T1586;
  wire T1587;
  wire T1588;
  wire T1589;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R8 = {1{$random}};
    R11 = {1{$random}};
    updateHit = {1{$random}};
    R18 = {1{$random}};
    for (initvar = 0; initvar < 128; initvar = initvar+1)
      T21[initvar] = {1{$random}};
    R38 = {1{$random}};
    isJump = {2{$random}};
    R55 = {1{$random}};
    R63 = {1{$random}};
    R67 = {1{$random}};
    pageValid = {1{$random}};
    R88 = {1{$random}};
    R101 = {2{$random}};
    for (initvar = 0; initvar < 6; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {2{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R1532 = {2{$random}};
    R1539 = {1{$random}};
    R1546 = {1{$random}};
    R1559 = {2{$random}};
    useRAS = {2{$random}};
    R1575 = {1{$random}};
  end
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_update_valid ? io_update_bits_target : R4;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T14 & updateTarget;
  assign updateTarget = T10 & R8;
  assign T9 = io_update_valid ? io_update_bits_taken : R8;
  assign T10 = updateValid & R11;
  assign T12 = io_update_valid ? io_update_bits_mispredict : R11;
  assign updateValid = R11 | updateHit;
  assign T13 = io_update_valid ? io_update_bits_prediction_valid : updateHit;
  assign T14 = R18 & T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = updateValid & T17;
  assign T17 = updateTarget ^ 1'h1;
  assign T1590 = reset ? 1'h0 : io_update_valid;
  assign io_resp_bits_bht_value = T19;
  assign T19 = T20;
  assign T20 = T21[T37];
  assign T23 = {io_update_bits_taken, T24};
  assign T24 = T29 | T25;
  assign T25 = T26 & io_update_bits_taken;
  assign T26 = T28 | T27;
  assign T27 = io_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T28 = io_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T29 = T31 & T30;
  assign T30 = io_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T31 = io_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T32 = T34 & T33;
  assign T33 = io_update_bits_isJump ^ 1'h1;
  assign T34 = io_update_valid & io_update_bits_prediction_valid;
  assign T35 = T36 ^ io_update_bits_prediction_bits_bht_history;
  assign T36 = io_update_bits_pc[4'h8:2'h2];
  assign T37 = T1067 ^ R38;
  assign T39 = T1066 ? T1064 : T40;
  assign T40 = T44 ? T41 : R38;
  assign T41 = {T43, T42};
  assign T42 = R38[3'h6:1'h1];
  assign T43 = T19[1'h0:1'h0];
  assign T44 = T1062 & T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 != 62'h0;
  assign T47 = hits & isJump;
  assign T1591 = T48[6'h3d:1'h0];
  assign T48 = T7 ? T49 : T1592;
  assign T1592 = {2'h0, isJump};
  assign T49 = T69 | T50;
  assign T50 = T1595 & T51;
  assign T51 = T53 | T1593;
  assign T1593 = {2'h0, T52};
  assign T52 = isJump ^ isJump;
  assign T53 = 1'h1 << T54;
  assign T54 = updateHit ? R63 : R55;
  assign T1594 = reset ? 6'h0 : T56;
  assign T56 = T60 ? T57 : R55;
  assign T57 = T59 ? 6'h0 : T58;
  assign T58 = R55 + 6'h1;
  assign T59 = R55 == 6'h3d;
  assign T60 = T14 & T61;
  assign T61 = T62 & updateValid;
  assign T62 = updateHit ^ 1'h1;
  assign T64 = io_update_valid ? io_update_bits_prediction_bits_entry : R63;
  assign T1595 = T65 ? 64'hffffffffffffffff : 64'h0;
  assign T65 = T66;
  assign T66 = R67;
  assign T68 = io_update_valid ? io_update_bits_isJump : R67;
  assign T69 = T1596 & T70;
  assign T70 = ~ T51;
  assign T1596 = {2'h0, isJump};
  assign hits = T481 & T71;
  assign T71 = T72;
  assign T72 = {T327, T73};
  assign T73 = {T253, T74};
  assign T74 = {T214, T75};
  assign T75 = {T195, T76};
  assign T76 = {T186, T77};
  assign T77 = {T182, T78};
  assign T78 = T79 != 6'h0;
  assign T79 = idxPagesOH_0 & pageHit;
  assign pageHit = T158 & pageValid;
  assign T1597 = T1598[3'h5:1'h0];
  assign T1598 = reset ? 8'h0 : T80;
  assign T80 = io_invalidate ? 8'h0 : T81;
  assign T81 = T157 ? T82 : T1599;
  assign T1599 = {2'h0, pageValid};
  assign T82 = T1605 | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T1600;
  assign T1600 = {2'h0, T83};
  assign T83 = T85 | T1601;
  assign T1601 = {5'h0, T84};
  assign T84 = idxPageUpdateOH[3'h5:3'h5];
  assign T85 = T86 << 1'h1;
  assign T86 = idxPageUpdateOH[3'h4:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? T1603 : idxPageRepl;
  assign idxPageRepl = T87;
  assign T87 = 1'h1 << R88;
  assign T1602 = reset ? 3'h0 : T89;
  assign T89 = T93 ? T90 : R88;
  assign T90 = T92 ? 3'h0 : T91;
  assign T91 = R88 + 3'h1;
  assign T92 = R88 == 3'h5;
  assign T93 = R18 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = updateTarget & T94;
  assign T94 = useUpdatePageHit ^ 1'h1;
  assign T1603 = {2'h0, updatePageHit};
  assign updatePageHit = T95 & pageValid;
  assign T95 = T96;
  assign T96 = {T142, T97};
  assign T97 = {T140, T98};
  assign T98 = {T138, T99};
  assign T99 = T103 == T100;
  assign T100 = R101 >> 4'hd;
  assign T102 = io_update_valid ? io_update_bits_pc : R101;
  assign T103 = pages[3'h0];
  assign T105 = T108 ? T107 : T106;
  assign T106 = R101 >> 4'hd;
  assign T107 = io_req_bits_addr >> 4'hd;
  assign T108 = T109 != 8'h0;
  assign T109 = idxPageUpdateOH & 8'h15;
  assign T110 = T14 & T111;
  assign T111 = T113 & T112;
  assign T112 = pageReplEn[3'h5:3'h5];
  assign T113 = T108 ? doTgtPageRepl : doIdxPageRepl;
  assign T115 = T14 & T116;
  assign T116 = T113 & T117;
  assign T117 = pageReplEn[2'h3:2'h3];
  assign T119 = T14 & T120;
  assign T120 = T113 & T121;
  assign T121 = pageReplEn[1'h1:1'h1];
  assign T123 = T108 ? T125 : T124;
  assign T124 = io_req_bits_addr >> 4'hd;
  assign T125 = R101 >> 4'hd;
  assign T126 = T14 & T127;
  assign T127 = T129 & T128;
  assign T128 = pageReplEn[3'h4:3'h4];
  assign T129 = T108 ? doIdxPageRepl : doTgtPageRepl;
  assign T131 = T14 & T132;
  assign T132 = T129 & T133;
  assign T133 = pageReplEn[2'h2:2'h2];
  assign T135 = T14 & T136;
  assign T136 = T129 & T137;
  assign T137 = pageReplEn[1'h0:1'h0];
  assign T138 = T139 == T100;
  assign T139 = pages[3'h1];
  assign T140 = T141 == T100;
  assign T141 = pages[3'h2];
  assign T142 = {T148, T143};
  assign T143 = {T146, T144};
  assign T144 = T145 == T100;
  assign T145 = pages[3'h3];
  assign T146 = T147 == T100;
  assign T147 = pages[3'h4];
  assign T148 = T149 == T100;
  assign T149 = pages[3'h5];
  assign useUpdatePageHit = updatePageHit != 6'h0;
  assign samePage = T151 == T150;
  assign T150 = io_req_bits_addr >> 4'hd;
  assign T151 = R101 >> 4'hd;
  assign doTgtPageRepl = T155 & T152;
  assign T152 = usePageHit ^ 1'h1;
  assign usePageHit = T153 != 8'h0;
  assign T153 = T1604 & T154;
  assign T154 = ~ idxPageReplEn;
  assign T1604 = {2'h0, pageHit};
  assign T155 = updateTarget & T156;
  assign T156 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0;
  assign T1605 = {2'h0, pageValid};
  assign T157 = T14 & doPageRepl;
  assign T158 = T159;
  assign T159 = {T169, T160};
  assign T160 = {T167, T161};
  assign T161 = {T165, T162};
  assign T162 = T164 == T163;
  assign T163 = io_req_bits_addr >> 4'hd;
  assign T164 = pages[3'h0];
  assign T165 = T166 == T163;
  assign T166 = pages[3'h1];
  assign T167 = T168 == T163;
  assign T168 = pages[3'h2];
  assign T169 = {T175, T170};
  assign T170 = {T173, T171};
  assign T171 = T172 == T163;
  assign T172 = pages[3'h3];
  assign T173 = T174 == T163;
  assign T174 = pages[3'h4];
  assign T175 = T176 == T163;
  assign T176 = pages[3'h5];
  assign idxPagesOH_0 = T177[3'h5:1'h0];
  assign T177 = 1'h1 << T178;
  assign T178 = idxPages[6'h0];
  assign T1606 = {T1616, T1607};
  assign T1607 = {T1615, T1608};
  assign T1608 = T1609[1'h1:1'h1];
  assign T1609 = T1614 | T1610;
  assign T1610 = T1611[1'h1:1'h0];
  assign T1611 = T1613 | T1612;
  assign T1612 = idxPageUpdateOH[2'h3:1'h0];
  assign T1613 = idxPageUpdateOH[3'h7:3'h4];
  assign T1614 = T1611[2'h3:2'h2];
  assign T1615 = T1614 != 2'h0;
  assign T1616 = T1613 != 4'h0;
  assign T180 = T7 & T181;
  assign T181 = T54 < 6'h3e;
  assign T182 = T183 != 6'h0;
  assign T183 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T184[3'h5:1'h0];
  assign T184 = 1'h1 << T185;
  assign T185 = idxPages[6'h1];
  assign T186 = {T191, T187};
  assign T187 = T188 != 6'h0;
  assign T188 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T189[3'h5:1'h0];
  assign T189 = 1'h1 << T190;
  assign T190 = idxPages[6'h2];
  assign T191 = T192 != 6'h0;
  assign T192 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T193[3'h5:1'h0];
  assign T193 = 1'h1 << T194;
  assign T194 = idxPages[6'h3];
  assign T195 = {T205, T196};
  assign T196 = {T201, T197};
  assign T197 = T198 != 6'h0;
  assign T198 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T199[3'h5:1'h0];
  assign T199 = 1'h1 << T200;
  assign T200 = idxPages[6'h4];
  assign T201 = T202 != 6'h0;
  assign T202 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T203[3'h5:1'h0];
  assign T203 = 1'h1 << T204;
  assign T204 = idxPages[6'h5];
  assign T205 = {T210, T206};
  assign T206 = T207 != 6'h0;
  assign T207 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T208[3'h5:1'h0];
  assign T208 = 1'h1 << T209;
  assign T209 = idxPages[6'h6];
  assign T210 = T211 != 6'h0;
  assign T211 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T212[3'h5:1'h0];
  assign T212 = 1'h1 << T213;
  assign T213 = idxPages[6'h7];
  assign T214 = {T234, T215};
  assign T215 = {T225, T216};
  assign T216 = {T221, T217};
  assign T217 = T218 != 6'h0;
  assign T218 = idxPagesOH_8 & pageHit;
  assign idxPagesOH_8 = T219[3'h5:1'h0];
  assign T219 = 1'h1 << T220;
  assign T220 = idxPages[6'h8];
  assign T221 = T222 != 6'h0;
  assign T222 = idxPagesOH_9 & pageHit;
  assign idxPagesOH_9 = T223[3'h5:1'h0];
  assign T223 = 1'h1 << T224;
  assign T224 = idxPages[6'h9];
  assign T225 = {T230, T226};
  assign T226 = T227 != 6'h0;
  assign T227 = idxPagesOH_10 & pageHit;
  assign idxPagesOH_10 = T228[3'h5:1'h0];
  assign T228 = 1'h1 << T229;
  assign T229 = idxPages[6'ha];
  assign T230 = T231 != 6'h0;
  assign T231 = idxPagesOH_11 & pageHit;
  assign idxPagesOH_11 = T232[3'h5:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = idxPages[6'hb];
  assign T234 = {T244, T235};
  assign T235 = {T240, T236};
  assign T236 = T237 != 6'h0;
  assign T237 = idxPagesOH_12 & pageHit;
  assign idxPagesOH_12 = T238[3'h5:1'h0];
  assign T238 = 1'h1 << T239;
  assign T239 = idxPages[6'hc];
  assign T240 = T241 != 6'h0;
  assign T241 = idxPagesOH_13 & pageHit;
  assign idxPagesOH_13 = T242[3'h5:1'h0];
  assign T242 = 1'h1 << T243;
  assign T243 = idxPages[6'hd];
  assign T244 = {T249, T245};
  assign T245 = T246 != 6'h0;
  assign T246 = idxPagesOH_14 & pageHit;
  assign idxPagesOH_14 = T247[3'h5:1'h0];
  assign T247 = 1'h1 << T248;
  assign T248 = idxPages[6'he];
  assign T249 = T250 != 6'h0;
  assign T250 = idxPagesOH_15 & pageHit;
  assign idxPagesOH_15 = T251[3'h5:1'h0];
  assign T251 = 1'h1 << T252;
  assign T252 = idxPages[6'hf];
  assign T253 = {T293, T254};
  assign T254 = {T274, T255};
  assign T255 = {T265, T256};
  assign T256 = {T261, T257};
  assign T257 = T258 != 6'h0;
  assign T258 = idxPagesOH_16 & pageHit;
  assign idxPagesOH_16 = T259[3'h5:1'h0];
  assign T259 = 1'h1 << T260;
  assign T260 = idxPages[6'h10];
  assign T261 = T262 != 6'h0;
  assign T262 = idxPagesOH_17 & pageHit;
  assign idxPagesOH_17 = T263[3'h5:1'h0];
  assign T263 = 1'h1 << T264;
  assign T264 = idxPages[6'h11];
  assign T265 = {T270, T266};
  assign T266 = T267 != 6'h0;
  assign T267 = idxPagesOH_18 & pageHit;
  assign idxPagesOH_18 = T268[3'h5:1'h0];
  assign T268 = 1'h1 << T269;
  assign T269 = idxPages[6'h12];
  assign T270 = T271 != 6'h0;
  assign T271 = idxPagesOH_19 & pageHit;
  assign idxPagesOH_19 = T272[3'h5:1'h0];
  assign T272 = 1'h1 << T273;
  assign T273 = idxPages[6'h13];
  assign T274 = {T284, T275};
  assign T275 = {T280, T276};
  assign T276 = T277 != 6'h0;
  assign T277 = idxPagesOH_20 & pageHit;
  assign idxPagesOH_20 = T278[3'h5:1'h0];
  assign T278 = 1'h1 << T279;
  assign T279 = idxPages[6'h14];
  assign T280 = T281 != 6'h0;
  assign T281 = idxPagesOH_21 & pageHit;
  assign idxPagesOH_21 = T282[3'h5:1'h0];
  assign T282 = 1'h1 << T283;
  assign T283 = idxPages[6'h15];
  assign T284 = {T289, T285};
  assign T285 = T286 != 6'h0;
  assign T286 = idxPagesOH_22 & pageHit;
  assign idxPagesOH_22 = T287[3'h5:1'h0];
  assign T287 = 1'h1 << T288;
  assign T288 = idxPages[6'h16];
  assign T289 = T290 != 6'h0;
  assign T290 = idxPagesOH_23 & pageHit;
  assign idxPagesOH_23 = T291[3'h5:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = idxPages[6'h17];
  assign T293 = {T313, T294};
  assign T294 = {T304, T295};
  assign T295 = {T300, T296};
  assign T296 = T297 != 6'h0;
  assign T297 = idxPagesOH_24 & pageHit;
  assign idxPagesOH_24 = T298[3'h5:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = idxPages[6'h18];
  assign T300 = T301 != 6'h0;
  assign T301 = idxPagesOH_25 & pageHit;
  assign idxPagesOH_25 = T302[3'h5:1'h0];
  assign T302 = 1'h1 << T303;
  assign T303 = idxPages[6'h19];
  assign T304 = {T309, T305};
  assign T305 = T306 != 6'h0;
  assign T306 = idxPagesOH_26 & pageHit;
  assign idxPagesOH_26 = T307[3'h5:1'h0];
  assign T307 = 1'h1 << T308;
  assign T308 = idxPages[6'h1a];
  assign T309 = T310 != 6'h0;
  assign T310 = idxPagesOH_27 & pageHit;
  assign idxPagesOH_27 = T311[3'h5:1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = idxPages[6'h1b];
  assign T313 = {T323, T314};
  assign T314 = {T319, T315};
  assign T315 = T316 != 6'h0;
  assign T316 = idxPagesOH_28 & pageHit;
  assign idxPagesOH_28 = T317[3'h5:1'h0];
  assign T317 = 1'h1 << T318;
  assign T318 = idxPages[6'h1c];
  assign T319 = T320 != 6'h0;
  assign T320 = idxPagesOH_29 & pageHit;
  assign idxPagesOH_29 = T321[3'h5:1'h0];
  assign T321 = 1'h1 << T322;
  assign T322 = idxPages[6'h1d];
  assign T323 = T324 != 6'h0;
  assign T324 = idxPagesOH_30 & pageHit;
  assign idxPagesOH_30 = T325[3'h5:1'h0];
  assign T325 = 1'h1 << T326;
  assign T326 = idxPages[6'h1e];
  assign T327 = {T407, T328};
  assign T328 = {T368, T329};
  assign T329 = {T349, T330};
  assign T330 = {T340, T331};
  assign T331 = {T336, T332};
  assign T332 = T333 != 6'h0;
  assign T333 = idxPagesOH_31 & pageHit;
  assign idxPagesOH_31 = T334[3'h5:1'h0];
  assign T334 = 1'h1 << T335;
  assign T335 = idxPages[6'h1f];
  assign T336 = T337 != 6'h0;
  assign T337 = idxPagesOH_32 & pageHit;
  assign idxPagesOH_32 = T338[3'h5:1'h0];
  assign T338 = 1'h1 << T339;
  assign T339 = idxPages[6'h20];
  assign T340 = {T345, T341};
  assign T341 = T342 != 6'h0;
  assign T342 = idxPagesOH_33 & pageHit;
  assign idxPagesOH_33 = T343[3'h5:1'h0];
  assign T343 = 1'h1 << T344;
  assign T344 = idxPages[6'h21];
  assign T345 = T346 != 6'h0;
  assign T346 = idxPagesOH_34 & pageHit;
  assign idxPagesOH_34 = T347[3'h5:1'h0];
  assign T347 = 1'h1 << T348;
  assign T348 = idxPages[6'h22];
  assign T349 = {T359, T350};
  assign T350 = {T355, T351};
  assign T351 = T352 != 6'h0;
  assign T352 = idxPagesOH_35 & pageHit;
  assign idxPagesOH_35 = T353[3'h5:1'h0];
  assign T353 = 1'h1 << T354;
  assign T354 = idxPages[6'h23];
  assign T355 = T356 != 6'h0;
  assign T356 = idxPagesOH_36 & pageHit;
  assign idxPagesOH_36 = T357[3'h5:1'h0];
  assign T357 = 1'h1 << T358;
  assign T358 = idxPages[6'h24];
  assign T359 = {T364, T360};
  assign T360 = T361 != 6'h0;
  assign T361 = idxPagesOH_37 & pageHit;
  assign idxPagesOH_37 = T362[3'h5:1'h0];
  assign T362 = 1'h1 << T363;
  assign T363 = idxPages[6'h25];
  assign T364 = T365 != 6'h0;
  assign T365 = idxPagesOH_38 & pageHit;
  assign idxPagesOH_38 = T366[3'h5:1'h0];
  assign T366 = 1'h1 << T367;
  assign T367 = idxPages[6'h26];
  assign T368 = {T388, T369};
  assign T369 = {T379, T370};
  assign T370 = {T375, T371};
  assign T371 = T372 != 6'h0;
  assign T372 = idxPagesOH_39 & pageHit;
  assign idxPagesOH_39 = T373[3'h5:1'h0];
  assign T373 = 1'h1 << T374;
  assign T374 = idxPages[6'h27];
  assign T375 = T376 != 6'h0;
  assign T376 = idxPagesOH_40 & pageHit;
  assign idxPagesOH_40 = T377[3'h5:1'h0];
  assign T377 = 1'h1 << T378;
  assign T378 = idxPages[6'h28];
  assign T379 = {T384, T380};
  assign T380 = T381 != 6'h0;
  assign T381 = idxPagesOH_41 & pageHit;
  assign idxPagesOH_41 = T382[3'h5:1'h0];
  assign T382 = 1'h1 << T383;
  assign T383 = idxPages[6'h29];
  assign T384 = T385 != 6'h0;
  assign T385 = idxPagesOH_42 & pageHit;
  assign idxPagesOH_42 = T386[3'h5:1'h0];
  assign T386 = 1'h1 << T387;
  assign T387 = idxPages[6'h2a];
  assign T388 = {T398, T389};
  assign T389 = {T394, T390};
  assign T390 = T391 != 6'h0;
  assign T391 = idxPagesOH_43 & pageHit;
  assign idxPagesOH_43 = T392[3'h5:1'h0];
  assign T392 = 1'h1 << T393;
  assign T393 = idxPages[6'h2b];
  assign T394 = T395 != 6'h0;
  assign T395 = idxPagesOH_44 & pageHit;
  assign idxPagesOH_44 = T396[3'h5:1'h0];
  assign T396 = 1'h1 << T397;
  assign T397 = idxPages[6'h2c];
  assign T398 = {T403, T399};
  assign T399 = T400 != 6'h0;
  assign T400 = idxPagesOH_45 & pageHit;
  assign idxPagesOH_45 = T401[3'h5:1'h0];
  assign T401 = 1'h1 << T402;
  assign T402 = idxPages[6'h2d];
  assign T403 = T404 != 6'h0;
  assign T404 = idxPagesOH_46 & pageHit;
  assign idxPagesOH_46 = T405[3'h5:1'h0];
  assign T405 = 1'h1 << T406;
  assign T406 = idxPages[6'h2e];
  assign T407 = {T447, T408};
  assign T408 = {T428, T409};
  assign T409 = {T419, T410};
  assign T410 = {T415, T411};
  assign T411 = T412 != 6'h0;
  assign T412 = idxPagesOH_47 & pageHit;
  assign idxPagesOH_47 = T413[3'h5:1'h0];
  assign T413 = 1'h1 << T414;
  assign T414 = idxPages[6'h2f];
  assign T415 = T416 != 6'h0;
  assign T416 = idxPagesOH_48 & pageHit;
  assign idxPagesOH_48 = T417[3'h5:1'h0];
  assign T417 = 1'h1 << T418;
  assign T418 = idxPages[6'h30];
  assign T419 = {T424, T420};
  assign T420 = T421 != 6'h0;
  assign T421 = idxPagesOH_49 & pageHit;
  assign idxPagesOH_49 = T422[3'h5:1'h0];
  assign T422 = 1'h1 << T423;
  assign T423 = idxPages[6'h31];
  assign T424 = T425 != 6'h0;
  assign T425 = idxPagesOH_50 & pageHit;
  assign idxPagesOH_50 = T426[3'h5:1'h0];
  assign T426 = 1'h1 << T427;
  assign T427 = idxPages[6'h32];
  assign T428 = {T438, T429};
  assign T429 = {T434, T430};
  assign T430 = T431 != 6'h0;
  assign T431 = idxPagesOH_51 & pageHit;
  assign idxPagesOH_51 = T432[3'h5:1'h0];
  assign T432 = 1'h1 << T433;
  assign T433 = idxPages[6'h33];
  assign T434 = T435 != 6'h0;
  assign T435 = idxPagesOH_52 & pageHit;
  assign idxPagesOH_52 = T436[3'h5:1'h0];
  assign T436 = 1'h1 << T437;
  assign T437 = idxPages[6'h34];
  assign T438 = {T443, T439};
  assign T439 = T440 != 6'h0;
  assign T440 = idxPagesOH_53 & pageHit;
  assign idxPagesOH_53 = T441[3'h5:1'h0];
  assign T441 = 1'h1 << T442;
  assign T442 = idxPages[6'h35];
  assign T443 = T444 != 6'h0;
  assign T444 = idxPagesOH_54 & pageHit;
  assign idxPagesOH_54 = T445[3'h5:1'h0];
  assign T445 = 1'h1 << T446;
  assign T446 = idxPages[6'h36];
  assign T447 = {T467, T448};
  assign T448 = {T458, T449};
  assign T449 = {T454, T450};
  assign T450 = T451 != 6'h0;
  assign T451 = idxPagesOH_55 & pageHit;
  assign idxPagesOH_55 = T452[3'h5:1'h0];
  assign T452 = 1'h1 << T453;
  assign T453 = idxPages[6'h37];
  assign T454 = T455 != 6'h0;
  assign T455 = idxPagesOH_56 & pageHit;
  assign idxPagesOH_56 = T456[3'h5:1'h0];
  assign T456 = 1'h1 << T457;
  assign T457 = idxPages[6'h38];
  assign T458 = {T463, T459};
  assign T459 = T460 != 6'h0;
  assign T460 = idxPagesOH_57 & pageHit;
  assign idxPagesOH_57 = T461[3'h5:1'h0];
  assign T461 = 1'h1 << T462;
  assign T462 = idxPages[6'h39];
  assign T463 = T464 != 6'h0;
  assign T464 = idxPagesOH_58 & pageHit;
  assign idxPagesOH_58 = T465[3'h5:1'h0];
  assign T465 = 1'h1 << T466;
  assign T466 = idxPages[6'h3a];
  assign T467 = {T477, T468};
  assign T468 = {T473, T469};
  assign T469 = T470 != 6'h0;
  assign T470 = idxPagesOH_59 & pageHit;
  assign idxPagesOH_59 = T471[3'h5:1'h0];
  assign T471 = 1'h1 << T472;
  assign T472 = idxPages[6'h3b];
  assign T473 = T474 != 6'h0;
  assign T474 = idxPagesOH_60 & pageHit;
  assign idxPagesOH_60 = T475[3'h5:1'h0];
  assign T475 = 1'h1 << T476;
  assign T476 = idxPages[6'h3c];
  assign T477 = T478 != 6'h0;
  assign T478 = idxPagesOH_61 & pageHit;
  assign idxPagesOH_61 = T479[3'h5:1'h0];
  assign T479 = 1'h1 << T480;
  assign T480 = idxPages[6'h3d];
  assign T481 = idxValid & T482;
  assign T482 = T483;
  assign T483 = {T580, T484};
  assign T484 = {T536, T485};
  assign T485 = {T513, T486};
  assign T486 = {T502, T487};
  assign T487 = {T497, T488};
  assign T488 = {T495, T489};
  assign T489 = T491 == T490;
  assign T490 = io_req_bits_addr[4'hc:1'h0];
  assign T491 = idxs[6'h0];
  assign T1617 = R101[4'hc:1'h0];
  assign T493 = T7 & T494;
  assign T494 = T54 < 6'h3e;
  assign T495 = T496 == T490;
  assign T496 = idxs[6'h1];
  assign T497 = {T500, T498};
  assign T498 = T499 == T490;
  assign T499 = idxs[6'h2];
  assign T500 = T501 == T490;
  assign T501 = idxs[6'h3];
  assign T502 = {T508, T503};
  assign T503 = {T506, T504};
  assign T504 = T505 == T490;
  assign T505 = idxs[6'h4];
  assign T506 = T507 == T490;
  assign T507 = idxs[6'h5];
  assign T508 = {T511, T509};
  assign T509 = T510 == T490;
  assign T510 = idxs[6'h6];
  assign T511 = T512 == T490;
  assign T512 = idxs[6'h7];
  assign T513 = {T525, T514};
  assign T514 = {T520, T515};
  assign T515 = {T518, T516};
  assign T516 = T517 == T490;
  assign T517 = idxs[6'h8];
  assign T518 = T519 == T490;
  assign T519 = idxs[6'h9];
  assign T520 = {T523, T521};
  assign T521 = T522 == T490;
  assign T522 = idxs[6'ha];
  assign T523 = T524 == T490;
  assign T524 = idxs[6'hb];
  assign T525 = {T531, T526};
  assign T526 = {T529, T527};
  assign T527 = T528 == T490;
  assign T528 = idxs[6'hc];
  assign T529 = T530 == T490;
  assign T530 = idxs[6'hd];
  assign T531 = {T534, T532};
  assign T532 = T533 == T490;
  assign T533 = idxs[6'he];
  assign T534 = T535 == T490;
  assign T535 = idxs[6'hf];
  assign T536 = {T560, T537};
  assign T537 = {T549, T538};
  assign T538 = {T544, T539};
  assign T539 = {T542, T540};
  assign T540 = T541 == T490;
  assign T541 = idxs[6'h10];
  assign T542 = T543 == T490;
  assign T543 = idxs[6'h11];
  assign T544 = {T547, T545};
  assign T545 = T546 == T490;
  assign T546 = idxs[6'h12];
  assign T547 = T548 == T490;
  assign T548 = idxs[6'h13];
  assign T549 = {T555, T550};
  assign T550 = {T553, T551};
  assign T551 = T552 == T490;
  assign T552 = idxs[6'h14];
  assign T553 = T554 == T490;
  assign T554 = idxs[6'h15];
  assign T555 = {T558, T556};
  assign T556 = T557 == T490;
  assign T557 = idxs[6'h16];
  assign T558 = T559 == T490;
  assign T559 = idxs[6'h17];
  assign T560 = {T572, T561};
  assign T561 = {T567, T562};
  assign T562 = {T565, T563};
  assign T563 = T564 == T490;
  assign T564 = idxs[6'h18];
  assign T565 = T566 == T490;
  assign T566 = idxs[6'h19];
  assign T567 = {T570, T568};
  assign T568 = T569 == T490;
  assign T569 = idxs[6'h1a];
  assign T570 = T571 == T490;
  assign T571 = idxs[6'h1b];
  assign T572 = {T578, T573};
  assign T573 = {T576, T574};
  assign T574 = T575 == T490;
  assign T575 = idxs[6'h1c];
  assign T576 = T577 == T490;
  assign T577 = idxs[6'h1d];
  assign T578 = T579 == T490;
  assign T579 = idxs[6'h1e];
  assign T580 = {T628, T581};
  assign T581 = {T605, T582};
  assign T582 = {T594, T583};
  assign T583 = {T589, T584};
  assign T584 = {T587, T585};
  assign T585 = T586 == T490;
  assign T586 = idxs[6'h1f];
  assign T587 = T588 == T490;
  assign T588 = idxs[6'h20];
  assign T589 = {T592, T590};
  assign T590 = T591 == T490;
  assign T591 = idxs[6'h21];
  assign T592 = T593 == T490;
  assign T593 = idxs[6'h22];
  assign T594 = {T600, T595};
  assign T595 = {T598, T596};
  assign T596 = T597 == T490;
  assign T597 = idxs[6'h23];
  assign T598 = T599 == T490;
  assign T599 = idxs[6'h24];
  assign T600 = {T603, T601};
  assign T601 = T602 == T490;
  assign T602 = idxs[6'h25];
  assign T603 = T604 == T490;
  assign T604 = idxs[6'h26];
  assign T605 = {T617, T606};
  assign T606 = {T612, T607};
  assign T607 = {T610, T608};
  assign T608 = T609 == T490;
  assign T609 = idxs[6'h27];
  assign T610 = T611 == T490;
  assign T611 = idxs[6'h28];
  assign T612 = {T615, T613};
  assign T613 = T614 == T490;
  assign T614 = idxs[6'h29];
  assign T615 = T616 == T490;
  assign T616 = idxs[6'h2a];
  assign T617 = {T623, T618};
  assign T618 = {T621, T619};
  assign T619 = T620 == T490;
  assign T620 = idxs[6'h2b];
  assign T621 = T622 == T490;
  assign T622 = idxs[6'h2c];
  assign T623 = {T626, T624};
  assign T624 = T625 == T490;
  assign T625 = idxs[6'h2d];
  assign T626 = T627 == T490;
  assign T627 = idxs[6'h2e];
  assign T628 = {T652, T629};
  assign T629 = {T641, T630};
  assign T630 = {T636, T631};
  assign T631 = {T634, T632};
  assign T632 = T633 == T490;
  assign T633 = idxs[6'h2f];
  assign T634 = T635 == T490;
  assign T635 = idxs[6'h30];
  assign T636 = {T639, T637};
  assign T637 = T638 == T490;
  assign T638 = idxs[6'h31];
  assign T639 = T640 == T490;
  assign T640 = idxs[6'h32];
  assign T641 = {T647, T642};
  assign T642 = {T645, T643};
  assign T643 = T644 == T490;
  assign T644 = idxs[6'h33];
  assign T645 = T646 == T490;
  assign T646 = idxs[6'h34];
  assign T647 = {T650, T648};
  assign T648 = T649 == T490;
  assign T649 = idxs[6'h35];
  assign T650 = T651 == T490;
  assign T651 = idxs[6'h36];
  assign T652 = {T664, T653};
  assign T653 = {T659, T654};
  assign T654 = {T657, T655};
  assign T655 = T656 == T490;
  assign T656 = idxs[6'h37];
  assign T657 = T658 == T490;
  assign T658 = idxs[6'h38];
  assign T659 = {T662, T660};
  assign T660 = T661 == T490;
  assign T661 = idxs[6'h39];
  assign T662 = T663 == T490;
  assign T663 = idxs[6'h3a];
  assign T664 = {T670, T665};
  assign T665 = {T668, T666};
  assign T666 = T667 == T490;
  assign T667 = idxs[6'h3b];
  assign T668 = T669 == T490;
  assign T669 = idxs[6'h3c];
  assign T670 = T671 == T490;
  assign T671 = idxs[6'h3d];
  assign T1618 = T1619[6'h3d:1'h0];
  assign T1619 = reset ? 64'h0 : T672;
  assign T672 = io_invalidate ? 64'h0 : T673;
  assign T673 = T14 ? T1053 : T1620;
  assign T1620 = {2'h0, T674};
  assign T674 = T14 ? T675 : idxValid;
  assign T675 = idxValid & T676;
  assign T676 = ~ T677;
  assign T677 = T678;
  assign T678 = {T868, T679};
  assign T679 = {T779, T680};
  assign T680 = {T732, T681};
  assign T681 = {T709, T682};
  assign T682 = {T698, T683};
  assign T683 = {T693, T684};
  assign T684 = T685 != 8'h0;
  assign T685 = pageReplEn & T1621;
  assign T1621 = {2'h0, T686};
  assign T686 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T687[3'h5:1'h0];
  assign T687 = 1'h1 << T688;
  assign T688 = tgtPages[6'h0];
  assign T1622 = {T1633, T1623};
  assign T1623 = {T1632, T1624};
  assign T1624 = T1625[1'h1:1'h1];
  assign T1625 = T1631 | T1626;
  assign T1626 = T1627[1'h1:1'h0];
  assign T1627 = T1630 | T1628;
  assign T1628 = T690[2'h3:1'h0];
  assign T690 = usePageHit ? T1629 : tgtPageRepl;
  assign T1629 = {2'h0, pageHit};
  assign T1630 = T690[3'h7:3'h4];
  assign T1631 = T1627[2'h3:2'h2];
  assign T1632 = T1631 != 2'h0;
  assign T1633 = T1630 != 4'h0;
  assign T691 = T7 & T692;
  assign T692 = T54 < 6'h3e;
  assign T693 = T694 != 8'h0;
  assign T694 = pageReplEn & T1634;
  assign T1634 = {2'h0, T695};
  assign T695 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T696[3'h5:1'h0];
  assign T696 = 1'h1 << T697;
  assign T697 = tgtPages[6'h1];
  assign T698 = {T704, T699};
  assign T699 = T700 != 8'h0;
  assign T700 = pageReplEn & T1635;
  assign T1635 = {2'h0, T701};
  assign T701 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T702[3'h5:1'h0];
  assign T702 = 1'h1 << T703;
  assign T703 = tgtPages[6'h2];
  assign T704 = T705 != 8'h0;
  assign T705 = pageReplEn & T1636;
  assign T1636 = {2'h0, T706};
  assign T706 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T707[3'h5:1'h0];
  assign T707 = 1'h1 << T708;
  assign T708 = tgtPages[6'h3];
  assign T709 = {T721, T710};
  assign T710 = {T716, T711};
  assign T711 = T712 != 8'h0;
  assign T712 = pageReplEn & T1637;
  assign T1637 = {2'h0, T713};
  assign T713 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T714[3'h5:1'h0];
  assign T714 = 1'h1 << T715;
  assign T715 = tgtPages[6'h4];
  assign T716 = T717 != 8'h0;
  assign T717 = pageReplEn & T1638;
  assign T1638 = {2'h0, T718};
  assign T718 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T719[3'h5:1'h0];
  assign T719 = 1'h1 << T720;
  assign T720 = tgtPages[6'h5];
  assign T721 = {T727, T722};
  assign T722 = T723 != 8'h0;
  assign T723 = pageReplEn & T1639;
  assign T1639 = {2'h0, T724};
  assign T724 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T725[3'h5:1'h0];
  assign T725 = 1'h1 << T726;
  assign T726 = tgtPages[6'h6];
  assign T727 = T728 != 8'h0;
  assign T728 = pageReplEn & T1640;
  assign T1640 = {2'h0, T729};
  assign T729 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T730[3'h5:1'h0];
  assign T730 = 1'h1 << T731;
  assign T731 = tgtPages[6'h7];
  assign T732 = {T756, T733};
  assign T733 = {T745, T734};
  assign T734 = {T740, T735};
  assign T735 = T736 != 8'h0;
  assign T736 = pageReplEn & T1641;
  assign T1641 = {2'h0, T737};
  assign T737 = idxPagesOH_8 | tgtPagesOH_8;
  assign tgtPagesOH_8 = T738[3'h5:1'h0];
  assign T738 = 1'h1 << T739;
  assign T739 = tgtPages[6'h8];
  assign T740 = T741 != 8'h0;
  assign T741 = pageReplEn & T1642;
  assign T1642 = {2'h0, T742};
  assign T742 = idxPagesOH_9 | tgtPagesOH_9;
  assign tgtPagesOH_9 = T743[3'h5:1'h0];
  assign T743 = 1'h1 << T744;
  assign T744 = tgtPages[6'h9];
  assign T745 = {T751, T746};
  assign T746 = T747 != 8'h0;
  assign T747 = pageReplEn & T1643;
  assign T1643 = {2'h0, T748};
  assign T748 = idxPagesOH_10 | tgtPagesOH_10;
  assign tgtPagesOH_10 = T749[3'h5:1'h0];
  assign T749 = 1'h1 << T750;
  assign T750 = tgtPages[6'ha];
  assign T751 = T752 != 8'h0;
  assign T752 = pageReplEn & T1644;
  assign T1644 = {2'h0, T753};
  assign T753 = idxPagesOH_11 | tgtPagesOH_11;
  assign tgtPagesOH_11 = T754[3'h5:1'h0];
  assign T754 = 1'h1 << T755;
  assign T755 = tgtPages[6'hb];
  assign T756 = {T768, T757};
  assign T757 = {T763, T758};
  assign T758 = T759 != 8'h0;
  assign T759 = pageReplEn & T1645;
  assign T1645 = {2'h0, T760};
  assign T760 = idxPagesOH_12 | tgtPagesOH_12;
  assign tgtPagesOH_12 = T761[3'h5:1'h0];
  assign T761 = 1'h1 << T762;
  assign T762 = tgtPages[6'hc];
  assign T763 = T764 != 8'h0;
  assign T764 = pageReplEn & T1646;
  assign T1646 = {2'h0, T765};
  assign T765 = idxPagesOH_13 | tgtPagesOH_13;
  assign tgtPagesOH_13 = T766[3'h5:1'h0];
  assign T766 = 1'h1 << T767;
  assign T767 = tgtPages[6'hd];
  assign T768 = {T774, T769};
  assign T769 = T770 != 8'h0;
  assign T770 = pageReplEn & T1647;
  assign T1647 = {2'h0, T771};
  assign T771 = idxPagesOH_14 | tgtPagesOH_14;
  assign tgtPagesOH_14 = T772[3'h5:1'h0];
  assign T772 = 1'h1 << T773;
  assign T773 = tgtPages[6'he];
  assign T774 = T775 != 8'h0;
  assign T775 = pageReplEn & T1648;
  assign T1648 = {2'h0, T776};
  assign T776 = idxPagesOH_15 | tgtPagesOH_15;
  assign tgtPagesOH_15 = T777[3'h5:1'h0];
  assign T777 = 1'h1 << T778;
  assign T778 = tgtPages[6'hf];
  assign T779 = {T827, T780};
  assign T780 = {T804, T781};
  assign T781 = {T793, T782};
  assign T782 = {T788, T783};
  assign T783 = T784 != 8'h0;
  assign T784 = pageReplEn & T1649;
  assign T1649 = {2'h0, T785};
  assign T785 = idxPagesOH_16 | tgtPagesOH_16;
  assign tgtPagesOH_16 = T786[3'h5:1'h0];
  assign T786 = 1'h1 << T787;
  assign T787 = tgtPages[6'h10];
  assign T788 = T789 != 8'h0;
  assign T789 = pageReplEn & T1650;
  assign T1650 = {2'h0, T790};
  assign T790 = idxPagesOH_17 | tgtPagesOH_17;
  assign tgtPagesOH_17 = T791[3'h5:1'h0];
  assign T791 = 1'h1 << T792;
  assign T792 = tgtPages[6'h11];
  assign T793 = {T799, T794};
  assign T794 = T795 != 8'h0;
  assign T795 = pageReplEn & T1651;
  assign T1651 = {2'h0, T796};
  assign T796 = idxPagesOH_18 | tgtPagesOH_18;
  assign tgtPagesOH_18 = T797[3'h5:1'h0];
  assign T797 = 1'h1 << T798;
  assign T798 = tgtPages[6'h12];
  assign T799 = T800 != 8'h0;
  assign T800 = pageReplEn & T1652;
  assign T1652 = {2'h0, T801};
  assign T801 = idxPagesOH_19 | tgtPagesOH_19;
  assign tgtPagesOH_19 = T802[3'h5:1'h0];
  assign T802 = 1'h1 << T803;
  assign T803 = tgtPages[6'h13];
  assign T804 = {T816, T805};
  assign T805 = {T811, T806};
  assign T806 = T807 != 8'h0;
  assign T807 = pageReplEn & T1653;
  assign T1653 = {2'h0, T808};
  assign T808 = idxPagesOH_20 | tgtPagesOH_20;
  assign tgtPagesOH_20 = T809[3'h5:1'h0];
  assign T809 = 1'h1 << T810;
  assign T810 = tgtPages[6'h14];
  assign T811 = T812 != 8'h0;
  assign T812 = pageReplEn & T1654;
  assign T1654 = {2'h0, T813};
  assign T813 = idxPagesOH_21 | tgtPagesOH_21;
  assign tgtPagesOH_21 = T814[3'h5:1'h0];
  assign T814 = 1'h1 << T815;
  assign T815 = tgtPages[6'h15];
  assign T816 = {T822, T817};
  assign T817 = T818 != 8'h0;
  assign T818 = pageReplEn & T1655;
  assign T1655 = {2'h0, T819};
  assign T819 = idxPagesOH_22 | tgtPagesOH_22;
  assign tgtPagesOH_22 = T820[3'h5:1'h0];
  assign T820 = 1'h1 << T821;
  assign T821 = tgtPages[6'h16];
  assign T822 = T823 != 8'h0;
  assign T823 = pageReplEn & T1656;
  assign T1656 = {2'h0, T824};
  assign T824 = idxPagesOH_23 | tgtPagesOH_23;
  assign tgtPagesOH_23 = T825[3'h5:1'h0];
  assign T825 = 1'h1 << T826;
  assign T826 = tgtPages[6'h17];
  assign T827 = {T851, T828};
  assign T828 = {T840, T829};
  assign T829 = {T835, T830};
  assign T830 = T831 != 8'h0;
  assign T831 = pageReplEn & T1657;
  assign T1657 = {2'h0, T832};
  assign T832 = idxPagesOH_24 | tgtPagesOH_24;
  assign tgtPagesOH_24 = T833[3'h5:1'h0];
  assign T833 = 1'h1 << T834;
  assign T834 = tgtPages[6'h18];
  assign T835 = T836 != 8'h0;
  assign T836 = pageReplEn & T1658;
  assign T1658 = {2'h0, T837};
  assign T837 = idxPagesOH_25 | tgtPagesOH_25;
  assign tgtPagesOH_25 = T838[3'h5:1'h0];
  assign T838 = 1'h1 << T839;
  assign T839 = tgtPages[6'h19];
  assign T840 = {T846, T841};
  assign T841 = T842 != 8'h0;
  assign T842 = pageReplEn & T1659;
  assign T1659 = {2'h0, T843};
  assign T843 = idxPagesOH_26 | tgtPagesOH_26;
  assign tgtPagesOH_26 = T844[3'h5:1'h0];
  assign T844 = 1'h1 << T845;
  assign T845 = tgtPages[6'h1a];
  assign T846 = T847 != 8'h0;
  assign T847 = pageReplEn & T1660;
  assign T1660 = {2'h0, T848};
  assign T848 = idxPagesOH_27 | tgtPagesOH_27;
  assign tgtPagesOH_27 = T849[3'h5:1'h0];
  assign T849 = 1'h1 << T850;
  assign T850 = tgtPages[6'h1b];
  assign T851 = {T863, T852};
  assign T852 = {T858, T853};
  assign T853 = T854 != 8'h0;
  assign T854 = pageReplEn & T1661;
  assign T1661 = {2'h0, T855};
  assign T855 = idxPagesOH_28 | tgtPagesOH_28;
  assign tgtPagesOH_28 = T856[3'h5:1'h0];
  assign T856 = 1'h1 << T857;
  assign T857 = tgtPages[6'h1c];
  assign T858 = T859 != 8'h0;
  assign T859 = pageReplEn & T1662;
  assign T1662 = {2'h0, T860};
  assign T860 = idxPagesOH_29 | tgtPagesOH_29;
  assign tgtPagesOH_29 = T861[3'h5:1'h0];
  assign T861 = 1'h1 << T862;
  assign T862 = tgtPages[6'h1d];
  assign T863 = T864 != 8'h0;
  assign T864 = pageReplEn & T1663;
  assign T1663 = {2'h0, T865};
  assign T865 = idxPagesOH_30 | tgtPagesOH_30;
  assign tgtPagesOH_30 = T866[3'h5:1'h0];
  assign T866 = 1'h1 << T867;
  assign T867 = tgtPages[6'h1e];
  assign T868 = {T964, T869};
  assign T869 = {T917, T870};
  assign T870 = {T894, T871};
  assign T871 = {T883, T872};
  assign T872 = {T878, T873};
  assign T873 = T874 != 8'h0;
  assign T874 = pageReplEn & T1664;
  assign T1664 = {2'h0, T875};
  assign T875 = idxPagesOH_31 | tgtPagesOH_31;
  assign tgtPagesOH_31 = T876[3'h5:1'h0];
  assign T876 = 1'h1 << T877;
  assign T877 = tgtPages[6'h1f];
  assign T878 = T879 != 8'h0;
  assign T879 = pageReplEn & T1665;
  assign T1665 = {2'h0, T880};
  assign T880 = idxPagesOH_32 | tgtPagesOH_32;
  assign tgtPagesOH_32 = T881[3'h5:1'h0];
  assign T881 = 1'h1 << T882;
  assign T882 = tgtPages[6'h20];
  assign T883 = {T889, T884};
  assign T884 = T885 != 8'h0;
  assign T885 = pageReplEn & T1666;
  assign T1666 = {2'h0, T886};
  assign T886 = idxPagesOH_33 | tgtPagesOH_33;
  assign tgtPagesOH_33 = T887[3'h5:1'h0];
  assign T887 = 1'h1 << T888;
  assign T888 = tgtPages[6'h21];
  assign T889 = T890 != 8'h0;
  assign T890 = pageReplEn & T1667;
  assign T1667 = {2'h0, T891};
  assign T891 = idxPagesOH_34 | tgtPagesOH_34;
  assign tgtPagesOH_34 = T892[3'h5:1'h0];
  assign T892 = 1'h1 << T893;
  assign T893 = tgtPages[6'h22];
  assign T894 = {T906, T895};
  assign T895 = {T901, T896};
  assign T896 = T897 != 8'h0;
  assign T897 = pageReplEn & T1668;
  assign T1668 = {2'h0, T898};
  assign T898 = idxPagesOH_35 | tgtPagesOH_35;
  assign tgtPagesOH_35 = T899[3'h5:1'h0];
  assign T899 = 1'h1 << T900;
  assign T900 = tgtPages[6'h23];
  assign T901 = T902 != 8'h0;
  assign T902 = pageReplEn & T1669;
  assign T1669 = {2'h0, T903};
  assign T903 = idxPagesOH_36 | tgtPagesOH_36;
  assign tgtPagesOH_36 = T904[3'h5:1'h0];
  assign T904 = 1'h1 << T905;
  assign T905 = tgtPages[6'h24];
  assign T906 = {T912, T907};
  assign T907 = T908 != 8'h0;
  assign T908 = pageReplEn & T1670;
  assign T1670 = {2'h0, T909};
  assign T909 = idxPagesOH_37 | tgtPagesOH_37;
  assign tgtPagesOH_37 = T910[3'h5:1'h0];
  assign T910 = 1'h1 << T911;
  assign T911 = tgtPages[6'h25];
  assign T912 = T913 != 8'h0;
  assign T913 = pageReplEn & T1671;
  assign T1671 = {2'h0, T914};
  assign T914 = idxPagesOH_38 | tgtPagesOH_38;
  assign tgtPagesOH_38 = T915[3'h5:1'h0];
  assign T915 = 1'h1 << T916;
  assign T916 = tgtPages[6'h26];
  assign T917 = {T941, T918};
  assign T918 = {T930, T919};
  assign T919 = {T925, T920};
  assign T920 = T921 != 8'h0;
  assign T921 = pageReplEn & T1672;
  assign T1672 = {2'h0, T922};
  assign T922 = idxPagesOH_39 | tgtPagesOH_39;
  assign tgtPagesOH_39 = T923[3'h5:1'h0];
  assign T923 = 1'h1 << T924;
  assign T924 = tgtPages[6'h27];
  assign T925 = T926 != 8'h0;
  assign T926 = pageReplEn & T1673;
  assign T1673 = {2'h0, T927};
  assign T927 = idxPagesOH_40 | tgtPagesOH_40;
  assign tgtPagesOH_40 = T928[3'h5:1'h0];
  assign T928 = 1'h1 << T929;
  assign T929 = tgtPages[6'h28];
  assign T930 = {T936, T931};
  assign T931 = T932 != 8'h0;
  assign T932 = pageReplEn & T1674;
  assign T1674 = {2'h0, T933};
  assign T933 = idxPagesOH_41 | tgtPagesOH_41;
  assign tgtPagesOH_41 = T934[3'h5:1'h0];
  assign T934 = 1'h1 << T935;
  assign T935 = tgtPages[6'h29];
  assign T936 = T937 != 8'h0;
  assign T937 = pageReplEn & T1675;
  assign T1675 = {2'h0, T938};
  assign T938 = idxPagesOH_42 | tgtPagesOH_42;
  assign tgtPagesOH_42 = T939[3'h5:1'h0];
  assign T939 = 1'h1 << T940;
  assign T940 = tgtPages[6'h2a];
  assign T941 = {T953, T942};
  assign T942 = {T948, T943};
  assign T943 = T944 != 8'h0;
  assign T944 = pageReplEn & T1676;
  assign T1676 = {2'h0, T945};
  assign T945 = idxPagesOH_43 | tgtPagesOH_43;
  assign tgtPagesOH_43 = T946[3'h5:1'h0];
  assign T946 = 1'h1 << T947;
  assign T947 = tgtPages[6'h2b];
  assign T948 = T949 != 8'h0;
  assign T949 = pageReplEn & T1677;
  assign T1677 = {2'h0, T950};
  assign T950 = idxPagesOH_44 | tgtPagesOH_44;
  assign tgtPagesOH_44 = T951[3'h5:1'h0];
  assign T951 = 1'h1 << T952;
  assign T952 = tgtPages[6'h2c];
  assign T953 = {T959, T954};
  assign T954 = T955 != 8'h0;
  assign T955 = pageReplEn & T1678;
  assign T1678 = {2'h0, T956};
  assign T956 = idxPagesOH_45 | tgtPagesOH_45;
  assign tgtPagesOH_45 = T957[3'h5:1'h0];
  assign T957 = 1'h1 << T958;
  assign T958 = tgtPages[6'h2d];
  assign T959 = T960 != 8'h0;
  assign T960 = pageReplEn & T1679;
  assign T1679 = {2'h0, T961};
  assign T961 = idxPagesOH_46 | tgtPagesOH_46;
  assign tgtPagesOH_46 = T962[3'h5:1'h0];
  assign T962 = 1'h1 << T963;
  assign T963 = tgtPages[6'h2e];
  assign T964 = {T1012, T965};
  assign T965 = {T989, T966};
  assign T966 = {T978, T967};
  assign T967 = {T973, T968};
  assign T968 = T969 != 8'h0;
  assign T969 = pageReplEn & T1680;
  assign T1680 = {2'h0, T970};
  assign T970 = idxPagesOH_47 | tgtPagesOH_47;
  assign tgtPagesOH_47 = T971[3'h5:1'h0];
  assign T971 = 1'h1 << T972;
  assign T972 = tgtPages[6'h2f];
  assign T973 = T974 != 8'h0;
  assign T974 = pageReplEn & T1681;
  assign T1681 = {2'h0, T975};
  assign T975 = idxPagesOH_48 | tgtPagesOH_48;
  assign tgtPagesOH_48 = T976[3'h5:1'h0];
  assign T976 = 1'h1 << T977;
  assign T977 = tgtPages[6'h30];
  assign T978 = {T984, T979};
  assign T979 = T980 != 8'h0;
  assign T980 = pageReplEn & T1682;
  assign T1682 = {2'h0, T981};
  assign T981 = idxPagesOH_49 | tgtPagesOH_49;
  assign tgtPagesOH_49 = T982[3'h5:1'h0];
  assign T982 = 1'h1 << T983;
  assign T983 = tgtPages[6'h31];
  assign T984 = T985 != 8'h0;
  assign T985 = pageReplEn & T1683;
  assign T1683 = {2'h0, T986};
  assign T986 = idxPagesOH_50 | tgtPagesOH_50;
  assign tgtPagesOH_50 = T987[3'h5:1'h0];
  assign T987 = 1'h1 << T988;
  assign T988 = tgtPages[6'h32];
  assign T989 = {T1001, T990};
  assign T990 = {T996, T991};
  assign T991 = T992 != 8'h0;
  assign T992 = pageReplEn & T1684;
  assign T1684 = {2'h0, T993};
  assign T993 = idxPagesOH_51 | tgtPagesOH_51;
  assign tgtPagesOH_51 = T994[3'h5:1'h0];
  assign T994 = 1'h1 << T995;
  assign T995 = tgtPages[6'h33];
  assign T996 = T997 != 8'h0;
  assign T997 = pageReplEn & T1685;
  assign T1685 = {2'h0, T998};
  assign T998 = idxPagesOH_52 | tgtPagesOH_52;
  assign tgtPagesOH_52 = T999[3'h5:1'h0];
  assign T999 = 1'h1 << T1000;
  assign T1000 = tgtPages[6'h34];
  assign T1001 = {T1007, T1002};
  assign T1002 = T1003 != 8'h0;
  assign T1003 = pageReplEn & T1686;
  assign T1686 = {2'h0, T1004};
  assign T1004 = idxPagesOH_53 | tgtPagesOH_53;
  assign tgtPagesOH_53 = T1005[3'h5:1'h0];
  assign T1005 = 1'h1 << T1006;
  assign T1006 = tgtPages[6'h35];
  assign T1007 = T1008 != 8'h0;
  assign T1008 = pageReplEn & T1687;
  assign T1687 = {2'h0, T1009};
  assign T1009 = idxPagesOH_54 | tgtPagesOH_54;
  assign tgtPagesOH_54 = T1010[3'h5:1'h0];
  assign T1010 = 1'h1 << T1011;
  assign T1011 = tgtPages[6'h36];
  assign T1012 = {T1036, T1013};
  assign T1013 = {T1025, T1014};
  assign T1014 = {T1020, T1015};
  assign T1015 = T1016 != 8'h0;
  assign T1016 = pageReplEn & T1688;
  assign T1688 = {2'h0, T1017};
  assign T1017 = idxPagesOH_55 | tgtPagesOH_55;
  assign tgtPagesOH_55 = T1018[3'h5:1'h0];
  assign T1018 = 1'h1 << T1019;
  assign T1019 = tgtPages[6'h37];
  assign T1020 = T1021 != 8'h0;
  assign T1021 = pageReplEn & T1689;
  assign T1689 = {2'h0, T1022};
  assign T1022 = idxPagesOH_56 | tgtPagesOH_56;
  assign tgtPagesOH_56 = T1023[3'h5:1'h0];
  assign T1023 = 1'h1 << T1024;
  assign T1024 = tgtPages[6'h38];
  assign T1025 = {T1031, T1026};
  assign T1026 = T1027 != 8'h0;
  assign T1027 = pageReplEn & T1690;
  assign T1690 = {2'h0, T1028};
  assign T1028 = idxPagesOH_57 | tgtPagesOH_57;
  assign tgtPagesOH_57 = T1029[3'h5:1'h0];
  assign T1029 = 1'h1 << T1030;
  assign T1030 = tgtPages[6'h39];
  assign T1031 = T1032 != 8'h0;
  assign T1032 = pageReplEn & T1691;
  assign T1691 = {2'h0, T1033};
  assign T1033 = idxPagesOH_58 | tgtPagesOH_58;
  assign tgtPagesOH_58 = T1034[3'h5:1'h0];
  assign T1034 = 1'h1 << T1035;
  assign T1035 = tgtPages[6'h3a];
  assign T1036 = {T1048, T1037};
  assign T1037 = {T1043, T1038};
  assign T1038 = T1039 != 8'h0;
  assign T1039 = pageReplEn & T1692;
  assign T1692 = {2'h0, T1040};
  assign T1040 = idxPagesOH_59 | tgtPagesOH_59;
  assign tgtPagesOH_59 = T1041[3'h5:1'h0];
  assign T1041 = 1'h1 << T1042;
  assign T1042 = tgtPages[6'h3b];
  assign T1043 = T1044 != 8'h0;
  assign T1044 = pageReplEn & T1693;
  assign T1693 = {2'h0, T1045};
  assign T1045 = idxPagesOH_60 | tgtPagesOH_60;
  assign tgtPagesOH_60 = T1046[3'h5:1'h0];
  assign T1046 = 1'h1 << T1047;
  assign T1047 = tgtPages[6'h3c];
  assign T1048 = T1049 != 8'h0;
  assign T1049 = pageReplEn & T1694;
  assign T1694 = {2'h0, T1050};
  assign T1050 = idxPagesOH_61 | tgtPagesOH_61;
  assign tgtPagesOH_61 = T1051[3'h5:1'h0];
  assign T1051 = 1'h1 << T1052;
  assign T1052 = tgtPages[6'h3d];
  assign T1053 = T1060 | T1054;
  assign T1054 = T1696 & T1055;
  assign T1055 = T1057 | T1695;
  assign T1695 = {2'h0, T1056};
  assign T1056 = idxValid ^ idxValid;
  assign T1057 = 1'h1 << T54;
  assign T1696 = T1058 ? 64'hffffffffffffffff : 64'h0;
  assign T1058 = T1059;
  assign T1059 = updateValid;
  assign T1060 = T1697 & T1061;
  assign T1061 = ~ T1055;
  assign T1697 = {2'h0, T674};
  assign T1062 = io_req_valid & T1063;
  assign T1063 = hits != 62'h0;
  assign T1064 = {io_update_bits_taken, T1065};
  assign T1065 = io_update_bits_prediction_bits_bht_history[3'h6:1'h1];
  assign T1066 = T32 & io_update_bits_mispredict;
  assign T1067 = io_req_bits_addr[4'h8:2'h2];
  assign io_resp_bits_bht_history = T1068;
  assign T1068 = R38;
  assign io_resp_bits_entry = T1698;
  assign T1698 = {T1723, T1699};
  assign T1699 = {T1722, T1700};
  assign T1700 = {T1721, T1701};
  assign T1701 = {T1720, T1702};
  assign T1702 = {T1719, T1703};
  assign T1703 = T1704[1'h1:1'h1];
  assign T1704 = T1718 | T1705;
  assign T1705 = T1706[1'h1:1'h0];
  assign T1706 = T1717 | T1707;
  assign T1707 = T1708[2'h3:1'h0];
  assign T1708 = T1716 | T1709;
  assign T1709 = T1710[3'h7:1'h0];
  assign T1710 = T1715 | T1711;
  assign T1711 = T1712[4'hf:1'h0];
  assign T1712 = T1714 | T1713;
  assign T1713 = hits[5'h1f:1'h0];
  assign T1714 = hits[6'h3d:6'h20];
  assign T1715 = T1712[5'h1f:5'h10];
  assign T1716 = T1710[4'hf:4'h8];
  assign T1717 = T1708[3'h7:3'h4];
  assign T1718 = T1706[2'h3:2'h2];
  assign T1719 = T1718 != 2'h0;
  assign T1720 = T1717 != 4'h0;
  assign T1721 = T1716 != 8'h0;
  assign T1722 = T1715 != 16'h0;
  assign T1723 = T1714 != 30'h0;
  assign io_resp_bits_target = T1070;
  assign T1070 = T1581 ? io_update_bits_returnAddr : T1071;
  assign T1071 = T1564 ? T1531 : T1072;
  assign T1072 = {T1323, T1073};
  assign T1073 = T1080 | T1074;
  assign T1074 = T1079 ? T1075 : 13'h0;
  assign T1075 = tgts[6'h3d];
  assign T1724 = io_req_bits_addr[4'hc:1'h0];
  assign T1077 = T7 & T1078;
  assign T1078 = T54 < 6'h3e;
  assign T1079 = hits[6'h3d:6'h3d];
  assign T1080 = T1084 | T1081;
  assign T1081 = T1083 ? T1082 : 13'h0;
  assign T1082 = tgts[6'h3c];
  assign T1083 = hits[6'h3c:6'h3c];
  assign T1084 = T1088 | T1085;
  assign T1085 = T1087 ? T1086 : 13'h0;
  assign T1086 = tgts[6'h3b];
  assign T1087 = hits[6'h3b:6'h3b];
  assign T1088 = T1092 | T1089;
  assign T1089 = T1091 ? T1090 : 13'h0;
  assign T1090 = tgts[6'h3a];
  assign T1091 = hits[6'h3a:6'h3a];
  assign T1092 = T1096 | T1093;
  assign T1093 = T1095 ? T1094 : 13'h0;
  assign T1094 = tgts[6'h39];
  assign T1095 = hits[6'h39:6'h39];
  assign T1096 = T1100 | T1097;
  assign T1097 = T1099 ? T1098 : 13'h0;
  assign T1098 = tgts[6'h38];
  assign T1099 = hits[6'h38:6'h38];
  assign T1100 = T1104 | T1101;
  assign T1101 = T1103 ? T1102 : 13'h0;
  assign T1102 = tgts[6'h37];
  assign T1103 = hits[6'h37:6'h37];
  assign T1104 = T1108 | T1105;
  assign T1105 = T1107 ? T1106 : 13'h0;
  assign T1106 = tgts[6'h36];
  assign T1107 = hits[6'h36:6'h36];
  assign T1108 = T1112 | T1109;
  assign T1109 = T1111 ? T1110 : 13'h0;
  assign T1110 = tgts[6'h35];
  assign T1111 = hits[6'h35:6'h35];
  assign T1112 = T1116 | T1113;
  assign T1113 = T1115 ? T1114 : 13'h0;
  assign T1114 = tgts[6'h34];
  assign T1115 = hits[6'h34:6'h34];
  assign T1116 = T1120 | T1117;
  assign T1117 = T1119 ? T1118 : 13'h0;
  assign T1118 = tgts[6'h33];
  assign T1119 = hits[6'h33:6'h33];
  assign T1120 = T1124 | T1121;
  assign T1121 = T1123 ? T1122 : 13'h0;
  assign T1122 = tgts[6'h32];
  assign T1123 = hits[6'h32:6'h32];
  assign T1124 = T1128 | T1125;
  assign T1125 = T1127 ? T1126 : 13'h0;
  assign T1126 = tgts[6'h31];
  assign T1127 = hits[6'h31:6'h31];
  assign T1128 = T1132 | T1129;
  assign T1129 = T1131 ? T1130 : 13'h0;
  assign T1130 = tgts[6'h30];
  assign T1131 = hits[6'h30:6'h30];
  assign T1132 = T1136 | T1133;
  assign T1133 = T1135 ? T1134 : 13'h0;
  assign T1134 = tgts[6'h2f];
  assign T1135 = hits[6'h2f:6'h2f];
  assign T1136 = T1140 | T1137;
  assign T1137 = T1139 ? T1138 : 13'h0;
  assign T1138 = tgts[6'h2e];
  assign T1139 = hits[6'h2e:6'h2e];
  assign T1140 = T1144 | T1141;
  assign T1141 = T1143 ? T1142 : 13'h0;
  assign T1142 = tgts[6'h2d];
  assign T1143 = hits[6'h2d:6'h2d];
  assign T1144 = T1148 | T1145;
  assign T1145 = T1147 ? T1146 : 13'h0;
  assign T1146 = tgts[6'h2c];
  assign T1147 = hits[6'h2c:6'h2c];
  assign T1148 = T1152 | T1149;
  assign T1149 = T1151 ? T1150 : 13'h0;
  assign T1150 = tgts[6'h2b];
  assign T1151 = hits[6'h2b:6'h2b];
  assign T1152 = T1156 | T1153;
  assign T1153 = T1155 ? T1154 : 13'h0;
  assign T1154 = tgts[6'h2a];
  assign T1155 = hits[6'h2a:6'h2a];
  assign T1156 = T1160 | T1157;
  assign T1157 = T1159 ? T1158 : 13'h0;
  assign T1158 = tgts[6'h29];
  assign T1159 = hits[6'h29:6'h29];
  assign T1160 = T1164 | T1161;
  assign T1161 = T1163 ? T1162 : 13'h0;
  assign T1162 = tgts[6'h28];
  assign T1163 = hits[6'h28:6'h28];
  assign T1164 = T1168 | T1165;
  assign T1165 = T1167 ? T1166 : 13'h0;
  assign T1166 = tgts[6'h27];
  assign T1167 = hits[6'h27:6'h27];
  assign T1168 = T1172 | T1169;
  assign T1169 = T1171 ? T1170 : 13'h0;
  assign T1170 = tgts[6'h26];
  assign T1171 = hits[6'h26:6'h26];
  assign T1172 = T1176 | T1173;
  assign T1173 = T1175 ? T1174 : 13'h0;
  assign T1174 = tgts[6'h25];
  assign T1175 = hits[6'h25:6'h25];
  assign T1176 = T1180 | T1177;
  assign T1177 = T1179 ? T1178 : 13'h0;
  assign T1178 = tgts[6'h24];
  assign T1179 = hits[6'h24:6'h24];
  assign T1180 = T1184 | T1181;
  assign T1181 = T1183 ? T1182 : 13'h0;
  assign T1182 = tgts[6'h23];
  assign T1183 = hits[6'h23:6'h23];
  assign T1184 = T1188 | T1185;
  assign T1185 = T1187 ? T1186 : 13'h0;
  assign T1186 = tgts[6'h22];
  assign T1187 = hits[6'h22:6'h22];
  assign T1188 = T1192 | T1189;
  assign T1189 = T1191 ? T1190 : 13'h0;
  assign T1190 = tgts[6'h21];
  assign T1191 = hits[6'h21:6'h21];
  assign T1192 = T1196 | T1193;
  assign T1193 = T1195 ? T1194 : 13'h0;
  assign T1194 = tgts[6'h20];
  assign T1195 = hits[6'h20:6'h20];
  assign T1196 = T1200 | T1197;
  assign T1197 = T1199 ? T1198 : 13'h0;
  assign T1198 = tgts[6'h1f];
  assign T1199 = hits[5'h1f:5'h1f];
  assign T1200 = T1204 | T1201;
  assign T1201 = T1203 ? T1202 : 13'h0;
  assign T1202 = tgts[6'h1e];
  assign T1203 = hits[5'h1e:5'h1e];
  assign T1204 = T1208 | T1205;
  assign T1205 = T1207 ? T1206 : 13'h0;
  assign T1206 = tgts[6'h1d];
  assign T1207 = hits[5'h1d:5'h1d];
  assign T1208 = T1212 | T1209;
  assign T1209 = T1211 ? T1210 : 13'h0;
  assign T1210 = tgts[6'h1c];
  assign T1211 = hits[5'h1c:5'h1c];
  assign T1212 = T1216 | T1213;
  assign T1213 = T1215 ? T1214 : 13'h0;
  assign T1214 = tgts[6'h1b];
  assign T1215 = hits[5'h1b:5'h1b];
  assign T1216 = T1220 | T1217;
  assign T1217 = T1219 ? T1218 : 13'h0;
  assign T1218 = tgts[6'h1a];
  assign T1219 = hits[5'h1a:5'h1a];
  assign T1220 = T1224 | T1221;
  assign T1221 = T1223 ? T1222 : 13'h0;
  assign T1222 = tgts[6'h19];
  assign T1223 = hits[5'h19:5'h19];
  assign T1224 = T1228 | T1225;
  assign T1225 = T1227 ? T1226 : 13'h0;
  assign T1226 = tgts[6'h18];
  assign T1227 = hits[5'h18:5'h18];
  assign T1228 = T1232 | T1229;
  assign T1229 = T1231 ? T1230 : 13'h0;
  assign T1230 = tgts[6'h17];
  assign T1231 = hits[5'h17:5'h17];
  assign T1232 = T1236 | T1233;
  assign T1233 = T1235 ? T1234 : 13'h0;
  assign T1234 = tgts[6'h16];
  assign T1235 = hits[5'h16:5'h16];
  assign T1236 = T1240 | T1237;
  assign T1237 = T1239 ? T1238 : 13'h0;
  assign T1238 = tgts[6'h15];
  assign T1239 = hits[5'h15:5'h15];
  assign T1240 = T1244 | T1241;
  assign T1241 = T1243 ? T1242 : 13'h0;
  assign T1242 = tgts[6'h14];
  assign T1243 = hits[5'h14:5'h14];
  assign T1244 = T1248 | T1245;
  assign T1245 = T1247 ? T1246 : 13'h0;
  assign T1246 = tgts[6'h13];
  assign T1247 = hits[5'h13:5'h13];
  assign T1248 = T1252 | T1249;
  assign T1249 = T1251 ? T1250 : 13'h0;
  assign T1250 = tgts[6'h12];
  assign T1251 = hits[5'h12:5'h12];
  assign T1252 = T1256 | T1253;
  assign T1253 = T1255 ? T1254 : 13'h0;
  assign T1254 = tgts[6'h11];
  assign T1255 = hits[5'h11:5'h11];
  assign T1256 = T1260 | T1257;
  assign T1257 = T1259 ? T1258 : 13'h0;
  assign T1258 = tgts[6'h10];
  assign T1259 = hits[5'h10:5'h10];
  assign T1260 = T1264 | T1261;
  assign T1261 = T1263 ? T1262 : 13'h0;
  assign T1262 = tgts[6'hf];
  assign T1263 = hits[4'hf:4'hf];
  assign T1264 = T1268 | T1265;
  assign T1265 = T1267 ? T1266 : 13'h0;
  assign T1266 = tgts[6'he];
  assign T1267 = hits[4'he:4'he];
  assign T1268 = T1272 | T1269;
  assign T1269 = T1271 ? T1270 : 13'h0;
  assign T1270 = tgts[6'hd];
  assign T1271 = hits[4'hd:4'hd];
  assign T1272 = T1276 | T1273;
  assign T1273 = T1275 ? T1274 : 13'h0;
  assign T1274 = tgts[6'hc];
  assign T1275 = hits[4'hc:4'hc];
  assign T1276 = T1280 | T1277;
  assign T1277 = T1279 ? T1278 : 13'h0;
  assign T1278 = tgts[6'hb];
  assign T1279 = hits[4'hb:4'hb];
  assign T1280 = T1284 | T1281;
  assign T1281 = T1283 ? T1282 : 13'h0;
  assign T1282 = tgts[6'ha];
  assign T1283 = hits[4'ha:4'ha];
  assign T1284 = T1288 | T1285;
  assign T1285 = T1287 ? T1286 : 13'h0;
  assign T1286 = tgts[6'h9];
  assign T1287 = hits[4'h9:4'h9];
  assign T1288 = T1292 | T1289;
  assign T1289 = T1291 ? T1290 : 13'h0;
  assign T1290 = tgts[6'h8];
  assign T1291 = hits[4'h8:4'h8];
  assign T1292 = T1296 | T1293;
  assign T1293 = T1295 ? T1294 : 13'h0;
  assign T1294 = tgts[6'h7];
  assign T1295 = hits[3'h7:3'h7];
  assign T1296 = T1300 | T1297;
  assign T1297 = T1299 ? T1298 : 13'h0;
  assign T1298 = tgts[6'h6];
  assign T1299 = hits[3'h6:3'h6];
  assign T1300 = T1304 | T1301;
  assign T1301 = T1303 ? T1302 : 13'h0;
  assign T1302 = tgts[6'h5];
  assign T1303 = hits[3'h5:3'h5];
  assign T1304 = T1308 | T1305;
  assign T1305 = T1307 ? T1306 : 13'h0;
  assign T1306 = tgts[6'h4];
  assign T1307 = hits[3'h4:3'h4];
  assign T1308 = T1312 | T1309;
  assign T1309 = T1311 ? T1310 : 13'h0;
  assign T1310 = tgts[6'h3];
  assign T1311 = hits[2'h3:2'h3];
  assign T1312 = T1316 | T1313;
  assign T1313 = T1315 ? T1314 : 13'h0;
  assign T1314 = tgts[6'h2];
  assign T1315 = hits[2'h2:2'h2];
  assign T1316 = T1320 | T1317;
  assign T1317 = T1319 ? T1318 : 13'h0;
  assign T1318 = tgts[6'h1];
  assign T1319 = hits[1'h1:1'h1];
  assign T1320 = T1322 ? T1321 : 13'h0;
  assign T1321 = tgts[6'h0];
  assign T1322 = hits[1'h0:1'h0];
  assign T1323 = T1512 | T1324;
  assign T1324 = T1326 ? T1325 : 30'h0;
  assign T1325 = pages[3'h5];
  assign T1326 = T1327[3'h5:3'h5];
  assign T1327 = T1330 | T1328;
  assign T1328 = T1329 ? tgtPagesOH_61 : 6'h0;
  assign T1329 = hits[6'h3d:6'h3d];
  assign T1330 = T1333 | T1331;
  assign T1331 = T1332 ? tgtPagesOH_60 : 6'h0;
  assign T1332 = hits[6'h3c:6'h3c];
  assign T1333 = T1336 | T1334;
  assign T1334 = T1335 ? tgtPagesOH_59 : 6'h0;
  assign T1335 = hits[6'h3b:6'h3b];
  assign T1336 = T1339 | T1337;
  assign T1337 = T1338 ? tgtPagesOH_58 : 6'h0;
  assign T1338 = hits[6'h3a:6'h3a];
  assign T1339 = T1342 | T1340;
  assign T1340 = T1341 ? tgtPagesOH_57 : 6'h0;
  assign T1341 = hits[6'h39:6'h39];
  assign T1342 = T1345 | T1343;
  assign T1343 = T1344 ? tgtPagesOH_56 : 6'h0;
  assign T1344 = hits[6'h38:6'h38];
  assign T1345 = T1348 | T1346;
  assign T1346 = T1347 ? tgtPagesOH_55 : 6'h0;
  assign T1347 = hits[6'h37:6'h37];
  assign T1348 = T1351 | T1349;
  assign T1349 = T1350 ? tgtPagesOH_54 : 6'h0;
  assign T1350 = hits[6'h36:6'h36];
  assign T1351 = T1354 | T1352;
  assign T1352 = T1353 ? tgtPagesOH_53 : 6'h0;
  assign T1353 = hits[6'h35:6'h35];
  assign T1354 = T1357 | T1355;
  assign T1355 = T1356 ? tgtPagesOH_52 : 6'h0;
  assign T1356 = hits[6'h34:6'h34];
  assign T1357 = T1360 | T1358;
  assign T1358 = T1359 ? tgtPagesOH_51 : 6'h0;
  assign T1359 = hits[6'h33:6'h33];
  assign T1360 = T1363 | T1361;
  assign T1361 = T1362 ? tgtPagesOH_50 : 6'h0;
  assign T1362 = hits[6'h32:6'h32];
  assign T1363 = T1366 | T1364;
  assign T1364 = T1365 ? tgtPagesOH_49 : 6'h0;
  assign T1365 = hits[6'h31:6'h31];
  assign T1366 = T1369 | T1367;
  assign T1367 = T1368 ? tgtPagesOH_48 : 6'h0;
  assign T1368 = hits[6'h30:6'h30];
  assign T1369 = T1372 | T1370;
  assign T1370 = T1371 ? tgtPagesOH_47 : 6'h0;
  assign T1371 = hits[6'h2f:6'h2f];
  assign T1372 = T1375 | T1373;
  assign T1373 = T1374 ? tgtPagesOH_46 : 6'h0;
  assign T1374 = hits[6'h2e:6'h2e];
  assign T1375 = T1378 | T1376;
  assign T1376 = T1377 ? tgtPagesOH_45 : 6'h0;
  assign T1377 = hits[6'h2d:6'h2d];
  assign T1378 = T1381 | T1379;
  assign T1379 = T1380 ? tgtPagesOH_44 : 6'h0;
  assign T1380 = hits[6'h2c:6'h2c];
  assign T1381 = T1384 | T1382;
  assign T1382 = T1383 ? tgtPagesOH_43 : 6'h0;
  assign T1383 = hits[6'h2b:6'h2b];
  assign T1384 = T1387 | T1385;
  assign T1385 = T1386 ? tgtPagesOH_42 : 6'h0;
  assign T1386 = hits[6'h2a:6'h2a];
  assign T1387 = T1390 | T1388;
  assign T1388 = T1389 ? tgtPagesOH_41 : 6'h0;
  assign T1389 = hits[6'h29:6'h29];
  assign T1390 = T1393 | T1391;
  assign T1391 = T1392 ? tgtPagesOH_40 : 6'h0;
  assign T1392 = hits[6'h28:6'h28];
  assign T1393 = T1396 | T1394;
  assign T1394 = T1395 ? tgtPagesOH_39 : 6'h0;
  assign T1395 = hits[6'h27:6'h27];
  assign T1396 = T1399 | T1397;
  assign T1397 = T1398 ? tgtPagesOH_38 : 6'h0;
  assign T1398 = hits[6'h26:6'h26];
  assign T1399 = T1402 | T1400;
  assign T1400 = T1401 ? tgtPagesOH_37 : 6'h0;
  assign T1401 = hits[6'h25:6'h25];
  assign T1402 = T1405 | T1403;
  assign T1403 = T1404 ? tgtPagesOH_36 : 6'h0;
  assign T1404 = hits[6'h24:6'h24];
  assign T1405 = T1408 | T1406;
  assign T1406 = T1407 ? tgtPagesOH_35 : 6'h0;
  assign T1407 = hits[6'h23:6'h23];
  assign T1408 = T1411 | T1409;
  assign T1409 = T1410 ? tgtPagesOH_34 : 6'h0;
  assign T1410 = hits[6'h22:6'h22];
  assign T1411 = T1414 | T1412;
  assign T1412 = T1413 ? tgtPagesOH_33 : 6'h0;
  assign T1413 = hits[6'h21:6'h21];
  assign T1414 = T1417 | T1415;
  assign T1415 = T1416 ? tgtPagesOH_32 : 6'h0;
  assign T1416 = hits[6'h20:6'h20];
  assign T1417 = T1420 | T1418;
  assign T1418 = T1419 ? tgtPagesOH_31 : 6'h0;
  assign T1419 = hits[5'h1f:5'h1f];
  assign T1420 = T1423 | T1421;
  assign T1421 = T1422 ? tgtPagesOH_30 : 6'h0;
  assign T1422 = hits[5'h1e:5'h1e];
  assign T1423 = T1426 | T1424;
  assign T1424 = T1425 ? tgtPagesOH_29 : 6'h0;
  assign T1425 = hits[5'h1d:5'h1d];
  assign T1426 = T1429 | T1427;
  assign T1427 = T1428 ? tgtPagesOH_28 : 6'h0;
  assign T1428 = hits[5'h1c:5'h1c];
  assign T1429 = T1432 | T1430;
  assign T1430 = T1431 ? tgtPagesOH_27 : 6'h0;
  assign T1431 = hits[5'h1b:5'h1b];
  assign T1432 = T1435 | T1433;
  assign T1433 = T1434 ? tgtPagesOH_26 : 6'h0;
  assign T1434 = hits[5'h1a:5'h1a];
  assign T1435 = T1438 | T1436;
  assign T1436 = T1437 ? tgtPagesOH_25 : 6'h0;
  assign T1437 = hits[5'h19:5'h19];
  assign T1438 = T1441 | T1439;
  assign T1439 = T1440 ? tgtPagesOH_24 : 6'h0;
  assign T1440 = hits[5'h18:5'h18];
  assign T1441 = T1444 | T1442;
  assign T1442 = T1443 ? tgtPagesOH_23 : 6'h0;
  assign T1443 = hits[5'h17:5'h17];
  assign T1444 = T1447 | T1445;
  assign T1445 = T1446 ? tgtPagesOH_22 : 6'h0;
  assign T1446 = hits[5'h16:5'h16];
  assign T1447 = T1450 | T1448;
  assign T1448 = T1449 ? tgtPagesOH_21 : 6'h0;
  assign T1449 = hits[5'h15:5'h15];
  assign T1450 = T1453 | T1451;
  assign T1451 = T1452 ? tgtPagesOH_20 : 6'h0;
  assign T1452 = hits[5'h14:5'h14];
  assign T1453 = T1456 | T1454;
  assign T1454 = T1455 ? tgtPagesOH_19 : 6'h0;
  assign T1455 = hits[5'h13:5'h13];
  assign T1456 = T1459 | T1457;
  assign T1457 = T1458 ? tgtPagesOH_18 : 6'h0;
  assign T1458 = hits[5'h12:5'h12];
  assign T1459 = T1462 | T1460;
  assign T1460 = T1461 ? tgtPagesOH_17 : 6'h0;
  assign T1461 = hits[5'h11:5'h11];
  assign T1462 = T1465 | T1463;
  assign T1463 = T1464 ? tgtPagesOH_16 : 6'h0;
  assign T1464 = hits[5'h10:5'h10];
  assign T1465 = T1468 | T1466;
  assign T1466 = T1467 ? tgtPagesOH_15 : 6'h0;
  assign T1467 = hits[4'hf:4'hf];
  assign T1468 = T1471 | T1469;
  assign T1469 = T1470 ? tgtPagesOH_14 : 6'h0;
  assign T1470 = hits[4'he:4'he];
  assign T1471 = T1474 | T1472;
  assign T1472 = T1473 ? tgtPagesOH_13 : 6'h0;
  assign T1473 = hits[4'hd:4'hd];
  assign T1474 = T1477 | T1475;
  assign T1475 = T1476 ? tgtPagesOH_12 : 6'h0;
  assign T1476 = hits[4'hc:4'hc];
  assign T1477 = T1480 | T1478;
  assign T1478 = T1479 ? tgtPagesOH_11 : 6'h0;
  assign T1479 = hits[4'hb:4'hb];
  assign T1480 = T1483 | T1481;
  assign T1481 = T1482 ? tgtPagesOH_10 : 6'h0;
  assign T1482 = hits[4'ha:4'ha];
  assign T1483 = T1486 | T1484;
  assign T1484 = T1485 ? tgtPagesOH_9 : 6'h0;
  assign T1485 = hits[4'h9:4'h9];
  assign T1486 = T1489 | T1487;
  assign T1487 = T1488 ? tgtPagesOH_8 : 6'h0;
  assign T1488 = hits[4'h8:4'h8];
  assign T1489 = T1492 | T1490;
  assign T1490 = T1491 ? tgtPagesOH_7 : 6'h0;
  assign T1491 = hits[3'h7:3'h7];
  assign T1492 = T1495 | T1493;
  assign T1493 = T1494 ? tgtPagesOH_6 : 6'h0;
  assign T1494 = hits[3'h6:3'h6];
  assign T1495 = T1498 | T1496;
  assign T1496 = T1497 ? tgtPagesOH_5 : 6'h0;
  assign T1497 = hits[3'h5:3'h5];
  assign T1498 = T1501 | T1499;
  assign T1499 = T1500 ? tgtPagesOH_4 : 6'h0;
  assign T1500 = hits[3'h4:3'h4];
  assign T1501 = T1504 | T1502;
  assign T1502 = T1503 ? tgtPagesOH_3 : 6'h0;
  assign T1503 = hits[2'h3:2'h3];
  assign T1504 = T1507 | T1505;
  assign T1505 = T1506 ? tgtPagesOH_2 : 6'h0;
  assign T1506 = hits[2'h2:2'h2];
  assign T1507 = T1510 | T1508;
  assign T1508 = T1509 ? tgtPagesOH_1 : 6'h0;
  assign T1509 = hits[1'h1:1'h1];
  assign T1510 = T1511 ? tgtPagesOH_0 : 6'h0;
  assign T1511 = hits[1'h0:1'h0];
  assign T1512 = T1516 | T1513;
  assign T1513 = T1515 ? T1514 : 30'h0;
  assign T1514 = pages[3'h4];
  assign T1515 = T1327[3'h4:3'h4];
  assign T1516 = T1520 | T1517;
  assign T1517 = T1519 ? T1518 : 30'h0;
  assign T1518 = pages[3'h3];
  assign T1519 = T1327[2'h3:2'h3];
  assign T1520 = T1524 | T1521;
  assign T1521 = T1523 ? T1522 : 30'h0;
  assign T1522 = pages[3'h2];
  assign T1523 = T1327[2'h2:2'h2];
  assign T1524 = T1528 | T1525;
  assign T1525 = T1527 ? T1526 : 30'h0;
  assign T1526 = pages[3'h1];
  assign T1527 = T1327[1'h1:1'h1];
  assign T1528 = T1530 ? T1529 : 30'h0;
  assign T1529 = pages[3'h0];
  assign T1530 = T1327[1'h0:1'h0];
  assign T1531 = T1563 ? R1559 : R1532;
  assign T1533 = T1534 ? io_update_bits_returnAddr : R1532;
  assign T1534 = T1558 & T1535;
  assign T1535 = T1536[1'h0:1'h0];
  assign T1536 = 1'h1 << T1537;
  assign T1537 = T1538;
  assign T1538 = R1539 + 1'h1;
  assign T1725 = reset ? 1'h0 : T1540;
  assign T1540 = T1543 ? T1542 : T1541;
  assign T1541 = T1558 ? T1538 : R1539;
  assign T1542 = R1539 - 1'h1;
  assign T1543 = T1554 & T1544;
  assign T1544 = T1545 ^ 1'h1;
  assign T1545 = R1546 == 2'h0;
  assign T1726 = reset ? 2'h0 : T1547;
  assign T1547 = io_invalidate ? 2'h0 : T1548;
  assign T1548 = T1543 ? T1553 : T1549;
  assign T1549 = T1551 ? T1550 : R1546;
  assign T1550 = R1546 + 2'h1;
  assign T1551 = T1558 & T1552;
  assign T1552 = R1546 < 2'h2;
  assign T1553 = R1546 - 2'h1;
  assign T1554 = io_update_valid & T1555;
  assign T1555 = T1557 & T1556;
  assign T1556 = io_update_bits_isReturn & io_update_bits_prediction_valid;
  assign T1557 = io_update_bits_isCall ^ 1'h1;
  assign T1558 = io_update_valid & io_update_bits_isCall;
  assign T1560 = T1561 ? io_update_bits_returnAddr : R1559;
  assign T1561 = T1558 & T1562;
  assign T1562 = T1536[1'h1:1'h1];
  assign T1563 = R1539;
  assign T1564 = T1579 & T1565;
  assign T1565 = T1566 != 62'h0;
  assign T1566 = hits & useRAS;
  assign T1727 = T1567[6'h3d:1'h0];
  assign T1567 = T7 ? T1568 : T1728;
  assign T1728 = {2'h0, useRAS};
  assign T1568 = T1577 | T1569;
  assign T1569 = T1730 & T1570;
  assign T1570 = T1572 | T1729;
  assign T1729 = {2'h0, T1571};
  assign T1571 = useRAS ^ useRAS;
  assign T1572 = 1'h1 << T54;
  assign T1730 = T1573 ? 64'hffffffffffffffff : 64'h0;
  assign T1573 = T1574;
  assign T1574 = R1575;
  assign T1576 = io_update_valid ? io_update_bits_isReturn : R1575;
  assign T1577 = T1731 & T1578;
  assign T1578 = ~ T1570;
  assign T1731 = {2'h0, useRAS};
  assign T1579 = T1580 ^ 1'h1;
  assign T1580 = R1546 == 2'h0;
  assign T1581 = T1558 & T1565;
  assign io_resp_bits_taken = T1582;
  assign T1582 = T1583 ? 1'h0 : io_resp_valid;
  assign T1583 = T1587 & T1584;
  assign T1584 = T1585 ^ 1'h1;
  assign T1585 = T1586 != 62'h0;
  assign T1586 = hits & isJump;
  assign T1587 = T1588 ^ 1'h1;
  assign T1588 = T19[1'h0:1'h0];
  assign io_resp_valid = T1589;
  assign T1589 = hits != 62'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
`endif
    if(io_update_valid) begin
      R4 <= io_update_bits_target;
    end
    if(io_update_valid) begin
      R8 <= io_update_bits_taken;
    end
    if(io_update_valid) begin
      R11 <= io_update_bits_mispredict;
    end
    if(io_update_valid) begin
      updateHit <= io_update_bits_prediction_valid;
    end
    if(reset) begin
      R18 <= 1'h0;
    end else begin
      R18 <= io_update_valid;
    end
    if (T32)
      T21[T35] <= T23;
    if(T1066) begin
      R38 <= T1064;
    end else if(T44) begin
      R38 <= T41;
    end
    isJump <= T1591;
    if(reset) begin
      R55 <= 6'h0;
    end else if(T60) begin
      R55 <= T57;
    end
    if(io_update_valid) begin
      R63 <= io_update_bits_prediction_bits_entry;
    end
    if(io_update_valid) begin
      R67 <= io_update_bits_isJump;
    end
    pageValid <= T1597;
    if(reset) begin
      R88 <= 3'h0;
    end else if(T93) begin
      R88 <= T90;
    end
    if(io_update_valid) begin
      R101 <= io_update_bits_pc;
    end
    if (T110)
      pages[3'h5] <= T105;
    if (T115)
      pages[3'h3] <= T105;
    if (T119)
      pages[3'h1] <= T105;
    if (T126)
      pages[3'h4] <= T123;
    if (T131)
      pages[3'h2] <= T123;
    if (T135)
      pages[3'h0] <= T123;
    if (T180)
      idxPages[T54] <= T1606;
    if (T493)
      idxs[T54] <= T1617;
    idxValid <= T1618;
    if (T691)
      tgtPages[T54] <= T1622;
    if (T1077)
      tgts[T54] <= T1724;
    if(T1534) begin
      R1532 <= io_update_bits_returnAddr;
    end
    if(reset) begin
      R1539 <= 1'h0;
    end else if(T1543) begin
      R1539 <= T1542;
    end else if(T1558) begin
      R1539 <= T1538;
    end
    if(reset) begin
      R1546 <= 2'h0;
    end else if(io_invalidate) begin
      R1546 <= 2'h0;
    end else if(T1543) begin
      R1546 <= T1553;
    end else if(T1551) begin
      R1546 <= T1550;
    end
    if(T1561) begin
      R1559 <= io_update_bits_returnAddr;
    end
    useRAS <= T1727;
    if(io_update_valid) begin
      R1575 <= io_update_bits_isReturn;
    end
  end
endmodule

module FlowThroughSerializer_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [2:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input  io_in_bits_payload_uncached,
    input [1:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T38;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T39;
  wire T4;
  wire T5;
  reg  active;
  wire T40;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire T9;
  wire[1:0] T10;
  reg [1:0] rbits_payload_g_type;
  wire[1:0] T41;
  wire[1:0] T11;
  wire T12;
  reg  rbits_payload_uncached;
  wire T42;
  wire T13;
  wire[2:0] T14;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T43;
  wire[2:0] T15;
  wire[2:0] T16;
  reg [2:0] rbits_payload_client_xact_id;
  wire[2:0] T44;
  wire[2:0] T17;
  wire[511:0] T18;
  wire[511:0] T19;
  reg [511:0] rbits_payload_data;
  wire[511:0] T45;
  wire[511:0] T20;
  wire[511:0] T46;
  wire[127:0] T21;
  wire[127:0] T22;
  wire[127:0] shifter_0;
  wire[127:0] T23;
  wire[127:0] shifter_1;
  wire[127:0] T24;
  wire T25;
  wire[1:0] T26;
  wire[127:0] T27;
  wire[127:0] shifter_2;
  wire[127:0] T28;
  wire[127:0] shifter_3;
  wire[127:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  reg [1:0] rbits_header_dst;
  wire[1:0] T47;
  wire[1:0] T33;
  wire[1:0] T34;
  reg [1:0] rbits_header_src;
  wire[1:0] T48;
  wire[1:0] T35;
  wire T36;
  wire T37;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cnt = {1{$random}};
    active = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_uncached = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T9 & wrap;
  assign wrap = cnt == 2'h3;
  assign T38 = reset ? 2'h0 : T1;
  assign T1 = T0 ? 2'h0 : T2;
  assign T2 = T9 ? T8 : T3;
  assign T3 = T4 ? T39 : cnt;
  assign T39 = {1'h0, io_out_ready};
  assign T4 = T5 & io_in_valid;
  assign T5 = active ^ 1'h1;
  assign T40 = reset ? 1'h0 : T6;
  assign T6 = T0 ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : active;
  assign T8 = cnt + 2'h1;
  assign T9 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T10;
  assign T10 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T41 = reset ? io_in_bits_payload_g_type : T11;
  assign T11 = T4 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_uncached = T12;
  assign T12 = active ? rbits_payload_uncached : io_in_bits_payload_uncached;
  assign T42 = reset ? io_in_bits_payload_uncached : T13;
  assign T13 = T4 ? io_in_bits_payload_uncached : rbits_payload_uncached;
  assign io_out_bits_payload_master_xact_id = T14;
  assign T14 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T43 = reset ? io_in_bits_payload_master_xact_id : T15;
  assign T15 = T4 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T16;
  assign T16 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T44 = reset ? io_in_bits_payload_client_xact_id : T17;
  assign T17 = T4 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T18;
  assign T18 = active ? T46 : T19;
  assign T19 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T45 = reset ? io_in_bits_payload_data : T20;
  assign T20 = T4 ? io_in_bits_payload_data : rbits_payload_data;
  assign T46 = {384'h0, T21};
  assign T21 = T31 ? T27 : T22;
  assign T22 = T25 ? shifter_1 : shifter_0;
  assign shifter_0 = T23;
  assign T23 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T24;
  assign T24 = rbits_payload_data[8'hff:8'h80];
  assign T25 = T26[1'h0:1'h0];
  assign T26 = cnt;
  assign T27 = T30 ? shifter_3 : shifter_2;
  assign shifter_2 = T28;
  assign T28 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T29;
  assign T29 = rbits_payload_data[9'h1ff:9'h180];
  assign T30 = T26[1'h0:1'h0];
  assign T31 = T26[1'h1:1'h1];
  assign io_out_bits_header_dst = T32;
  assign T32 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T47 = reset ? io_in_bits_header_dst : T33;
  assign T33 = T4 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T34;
  assign T34 = active ? rbits_header_src : io_in_bits_header_src;
  assign T48 = reset ? io_in_bits_header_src : T35;
  assign T35 = T4 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T36;
  assign T36 = active | io_in_valid;
  assign io_in_ready = T37;
  assign T37 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      cnt <= 2'h0;
    end else if(T0) begin
      cnt <= 2'h0;
    end else if(T9) begin
      cnt <= T8;
    end else if(T4) begin
      cnt <= T39;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T0) begin
      active <= 1'h0;
    end else if(T4) begin
      active <= 1'h1;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T4) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_uncached <= io_in_bits_payload_uncached;
    end else if(T4) begin
      rbits_payload_uncached <= io_in_bits_payload_uncached;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T4) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T4) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T4) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T4) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T4) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output io_count
);

  wire T13;
  wire[1:0] T0;
  reg  full;
  wire T14;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[2:0] T3;
  wire[6:0] T4;
  reg [6:0] ram [0:0];
  wire[6:0] T5;
  wire[6:0] T6;
  wire[6:0] T7;
  wire[4:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire empty;
  wire T12;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T13;
  assign T13 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T14 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T3;
  assign T3 = T4[2'h2:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign io_deq_bits_header_dst = T9;
  assign T9 = T4[3'h4:2'h3];
  assign io_deq_bits_header_src = T10;
  assign T10 = T4[3'h6:3'h5];
  assign io_deq_valid = T11;
  assign T11 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [12:0] io_req_bits_idx,
    input [18:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[2:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[511:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire T208;
  wire T209;
  wire T210;
  wire[511:0] T0;
  wire[1:0] T1;
  wire T2;
  wire[511:0] T3;
  wire[2:0] T4;
  wire[25:0] T5;
  wire[25:0] T6;
  reg [31:0] s2_addr;
  wire[31:0] T7;
  wire[31:0] s1_addr;
  wire[31:0] T8;
  reg [12:0] s1_pgoff;
  wire[12:0] T9;
  wire T10;
  wire rdy;
  wire T11;
  wire T12;
  wire s2_miss;
  wire T13;
  wire s2_any_tag_hit;
  wire T14;
  wire T15;
  wire T16;
  wire s2_disparity_1;
  wire T17;
  reg  R18;
  wire T19;
  wire T20;
  wire T21;
  wire stall;
  wire T22;
  reg  s1_valid;
  wire T196;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  reg  R28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[6:0] T37;
  wire T38;
  reg [255:0] vb_array;
  wire[255:0] T197;
  wire[255:0] T39;
  wire[255:0] T40;
  wire[255:0] T41;
  wire[255:0] T42;
  wire[255:0] T43;
  wire[255:0] T44;
  wire[255:0] T45;
  wire[7:0] T46;
  wire[6:0] s2_idx;
  wire repl_way;
  reg [15:0] R47;
  wire[15:0] T198;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[14:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[255:0] T199;
  wire T58;
  wire[255:0] T59;
  wire[255:0] T60;
  wire T61;
  wire T62;
  reg  invalidated;
  wire T63;
  wire T64;
  wire T65;
  reg [1:0] state;
  wire[1:0] T200;
  wire[1:0] T66;
  wire[1:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[255:0] T78;
  wire[255:0] T79;
  wire[255:0] T80;
  wire[7:0] T81;
  wire[255:0] T201;
  wire T82;
  wire[255:0] T83;
  wire[255:0] T84;
  wire T85;
  wire[255:0] T86;
  wire[255:0] T87;
  wire[255:0] T88;
  wire[7:0] T89;
  wire[255:0] T202;
  wire T90;
  wire[255:0] T91;
  wire[255:0] T92;
  wire T93;
  wire s2_disparity_0;
  wire T94;
  reg  R95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  reg  R100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[6:0] T109;
  wire T110;
  wire T111;
  wire s2_tag_hit_1;
  wire T112;
  reg  R113;
  wire T114;
  wire s1_tag_match_1;
  wire T115;
  wire[18:0] s1_tag;
  wire[18:0] T116;
  wire[18:0] T117;
  wire[37:0] T118;
  wire T132;
  wire s0_valid;
  wire T133;
  wire T134;
  wire[6:0] T130;
  wire[12:0] s0_pgoff;
  wire T131;
  wire[37:0] T119;
  wire[37:0] T120;
  wire[37:0] T121;
  wire[18:0] T122;
  wire[18:0] T203;
  wire T123;
  wire[1:0] T124;
  wire[18:0] T125;
  wire[18:0] T204;
  wire T126;
  wire[37:0] T127;
  wire[18:0] T128;
  wire[18:0] s2_tag;
  reg [6:0] tag_raddr;
  wire[6:0] T129;
  wire s2_tag_hit_0;
  wire T135;
  reg  R136;
  wire T137;
  wire s1_tag_match_0;
  wire T138;
  wire[18:0] T139;
  wire[18:0] T140;
  reg  s2_valid;
  wire T205;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[127:0] T152;
  wire[127:0] T153;
  reg [127:0] s2_dout_1;
  wire[127:0] T154;
  wire[127:0] T155;
  wire T164;
  wire T165;
  wire T158;
  wire T159;
  wire[8:0] T163;
  wire[127:0] T157;
  wire[127:0] T206;
  wire[8:0] T160;
  reg [8:0] R161;
  wire[8:0] T162;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[127:0] T170;
  reg [127:0] s2_dout_0;
  wire[127:0] T171;
  wire[127:0] T172;
  wire T181;
  wire T182;
  wire T175;
  wire T176;
  wire[8:0] T180;
  wire[127:0] T174;
  wire[127:0] T207;
  wire[8:0] T177;
  reg [8:0] R178;
  wire[8:0] T179;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[31:0] T187;
  wire[31:0] T188;
  wire[31:0] s2_dout_word_1;
  wire[127:0] T189;
  wire[6:0] T190;
  wire[1:0] T191;
  wire[5:0] s2_offset;
  wire[31:0] T192;
  wire[31:0] s2_dout_word_0;
  wire[127:0] T193;
  wire[6:0] T194;
  wire[1:0] T195;
  wire s2_hit;
  wire FlowThroughSerializer_1_io_in_ready;
  wire FlowThroughSerializer_1_io_out_valid;
  wire[1:0] FlowThroughSerializer_1_io_out_bits_header_src;
  wire[511:0] FlowThroughSerializer_1_io_out_bits_payload_data;
  wire[2:0] FlowThroughSerializer_1_io_out_bits_payload_master_xact_id;
  wire FlowThroughSerializer_1_io_out_bits_payload_uncached;
  wire[1:0] FlowThroughSerializer_1_io_out_bits_payload_g_type;
  wire[1:0] FlowThroughSerializer_1_io_cnt;
  wire FlowThroughSerializer_1_io_done;
  wire ack_q_io_enq_ready;
  wire ack_q_io_deq_valid;
  wire[1:0] ack_q_io_deq_bits_header_src;
  wire[1:0] ack_q_io_deq_bits_header_dst;
  wire[2:0] ack_q_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R18 = {1{$random}};
    s1_valid = {1{$random}};
    R28 = {1{$random}};
    vb_array = {8{$random}};
    R47 = {1{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    R95 = {1{$random}};
    R100 = {1{$random}};
    R113 = {1{$random}};
    tag_raddr = {1{$random}};
    R136 = {1{$random}};
    s2_valid = {1{$random}};
    s2_dout_1 = {4{$random}};
    R161 = {1{$random}};
    s2_dout_0 = {4{$random}};
    R178 = {1{$random}};
  end
`endif

  assign T208 = FlowThroughSerializer_1_io_done & T209;
  assign T209 = FlowThroughSerializer_1_io_out_bits_payload_uncached | T210;
  assign T210 = FlowThroughSerializer_1_io_out_bits_payload_g_type != 2'h0;
  assign io_mem_finish_bits_payload_master_xact_id = ack_q_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ack_q_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ack_q_io_deq_bits_header_src;
  assign io_mem_finish_valid = ack_q_io_deq_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign io_mem_acquire_bits_payload_subblock = T0;
  assign T0 = 512'h7;
  assign io_mem_acquire_bits_payload_a_type = T1;
  assign T1 = 2'h0;
  assign io_mem_acquire_bits_payload_uncached = T2;
  assign T2 = 1'h1;
  assign io_mem_acquire_bits_payload_data = T3;
  assign T3 = 512'h0;
  assign io_mem_acquire_bits_payload_client_xact_id = T4;
  assign T4 = 3'h0;
  assign io_mem_acquire_bits_payload_addr = T5;
  assign T5 = T6;
  assign T6 = s2_addr >> 3'h6;
  assign T7 = T147 ? s1_addr : s2_addr;
  assign s1_addr = T8;
  assign T8 = {io_req_bits_ppn, s1_pgoff};
  assign T9 = T10 ? io_req_bits_idx : s1_pgoff;
  assign T10 = io_req_valid & rdy;
  assign rdy = T11;
  assign T11 = T146 & T12;
  assign T12 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T13;
  assign T13 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T14;
  assign T14 = T111 & T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = s2_disparity_0 | s2_disparity_1;
  assign s2_disparity_1 = T17;
  assign T17 = R28 & R18;
  assign T19 = T20 ? 1'h0 : R18;
  assign T20 = T22 & T21;
  assign T21 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T22 = s1_valid & rdy;
  assign T196 = reset ? 1'h0 : T23;
  assign T23 = T27 | T24;
  assign T24 = T26 & T25;
  assign T25 = io_req_bits_kill ^ 1'h1;
  assign T26 = s1_valid & stall;
  assign T27 = io_req_valid & rdy;
  assign T29 = T20 ? T30 : R28;
  assign T30 = T31;
  assign T31 = T38 & T32;
  assign T32 = T33 - 1'h1;
  assign T33 = 1'h1 << T34;
  assign T34 = T35 + 8'h1;
  assign T35 = T36 - T36;
  assign T36 = {1'h1, T37};
  assign T37 = s1_pgoff[4'hc:3'h6];
  assign T38 = vb_array >> T36;
  assign T197 = reset ? 256'h0 : T39;
  assign T39 = T93 ? T86 : T40;
  assign T40 = T85 ? T78 : T41;
  assign T41 = io_invalidate ? 256'h0 : T42;
  assign T42 = T61 ? T43 : vb_array;
  assign T43 = T59 | T44;
  assign T44 = T199 & T45;
  assign T45 = 1'h1 << T46;
  assign T46 = {repl_way, s2_idx};
  assign s2_idx = s2_addr[4'hc:3'h6];
  assign repl_way = R47[1'h0:1'h0];
  assign T198 = reset ? 16'h1 : T48;
  assign T48 = s2_miss ? T49 : R47;
  assign T49 = {T51, T50};
  assign T50 = R47[4'hf:1'h1];
  assign T51 = T53 ^ T52;
  assign T52 = R47[3'h5:3'h5];
  assign T53 = T55 ^ T54;
  assign T54 = R47[2'h3:2'h3];
  assign T55 = T57 ^ T56;
  assign T56 = R47[2'h2:2'h2];
  assign T57 = R47[1'h0:1'h0];
  assign T199 = T58 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T58 = 1'h1;
  assign T59 = vb_array & T60;
  assign T60 = ~ T45;
  assign T61 = FlowThroughSerializer_1_io_done & T62;
  assign T62 = invalidated ^ 1'h1;
  assign T63 = T65 ? 1'h0 : T64;
  assign T64 = io_invalidate ? 1'h1 : invalidated;
  assign T65 = 2'h0 == state;
  assign T200 = reset ? 2'h0 : T66;
  assign T66 = T76 ? 2'h0 : T67;
  assign T67 = T74 ? 2'h3 : T68;
  assign T68 = T71 ? 2'h2 : T69;
  assign T69 = T70 ? 2'h1 : state;
  assign T70 = T65 & s2_miss;
  assign T71 = T73 & T72;
  assign T72 = io_mem_acquire_ready & ack_q_io_enq_ready;
  assign T73 = 2'h1 == state;
  assign T74 = T75 & io_mem_grant_valid;
  assign T75 = 2'h2 == state;
  assign T76 = T77 & FlowThroughSerializer_1_io_done;
  assign T77 = 2'h3 == state;
  assign T78 = T83 | T79;
  assign T79 = T201 & T80;
  assign T80 = 1'h1 << T81;
  assign T81 = {1'h0, s2_idx};
  assign T201 = T82 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T82 = 1'h0;
  assign T83 = vb_array & T84;
  assign T84 = ~ T80;
  assign T85 = s2_valid & s2_disparity_0;
  assign T86 = T91 | T87;
  assign T87 = T202 & T88;
  assign T88 = 1'h1 << T89;
  assign T89 = {1'h1, s2_idx};
  assign T202 = T90 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T90 = 1'h0;
  assign T91 = vb_array & T92;
  assign T92 = ~ T88;
  assign T93 = s2_valid & s2_disparity_1;
  assign s2_disparity_0 = T94;
  assign T94 = R100 & R95;
  assign T96 = T97 ? 1'h0 : R95;
  assign T97 = T99 & T98;
  assign T98 = stall ^ 1'h1;
  assign T99 = s1_valid & rdy;
  assign T101 = T97 ? T102 : R100;
  assign T102 = T103;
  assign T103 = T110 & T104;
  assign T104 = T105 - 1'h1;
  assign T105 = 1'h1 << T106;
  assign T106 = T107 + 8'h1;
  assign T107 = T108 - T108;
  assign T108 = {1'h0, T109};
  assign T109 = s1_pgoff[4'hc:3'h6];
  assign T110 = vb_array >> T108;
  assign T111 = s2_tag_hit_0 | s2_tag_hit_1;
  assign s2_tag_hit_1 = T112;
  assign T112 = R28 & R113;
  assign T114 = T20 ? s1_tag_match_1 : R113;
  assign s1_tag_match_1 = T115;
  assign T115 = T116 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hd];
  assign T116 = T117[5'h12:1'h0];
  assign T117 = T118[6'h25:5'h13];
  assign T132 = T134 & s0_valid;
  assign s0_valid = io_req_valid | T133;
  assign T133 = s1_valid & stall;
  assign T134 = FlowThroughSerializer_1_io_done ^ 1'h1;
  assign T130 = s0_pgoff[4'hc:3'h6];
  assign s0_pgoff = T131 ? s1_pgoff : io_req_bits_idx;
  assign T131 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_1_io_done ? s2_idx : T130),
    .RW0E(T132 || FlowThroughSerializer_1_io_done),
    .RW0W(FlowThroughSerializer_1_io_done),
    .RW0I(T127),
    .RW0M(T120),
    .RW0O(T118)
  );
  assign T120 = T121;
  assign T121 = {T125, T122};
  assign T122 = 19'h0 - T203;
  assign T203 = {18'h0, T123};
  assign T123 = T124[1'h0:1'h0];
  assign T124 = 1'h1 << repl_way;
  assign T125 = 19'h0 - T204;
  assign T204 = {18'h0, T126};
  assign T126 = T124[1'h1:1'h1];
  assign T127 = {T128, T128};
  assign T128 = s2_tag;
  assign s2_tag = s2_addr[5'h1f:4'hd];
  assign T129 = T132 ? T130 : tag_raddr;
  assign s2_tag_hit_0 = T135;
  assign T135 = R100 & R136;
  assign T137 = T97 ? s1_tag_match_0 : R136;
  assign s1_tag_match_0 = T138;
  assign T138 = T139 == s1_tag;
  assign T139 = T140[5'h12:1'h0];
  assign T140 = T118[5'h12:1'h0];
  assign T205 = reset ? 1'h0 : T141;
  assign T141 = T143 | T142;
  assign T142 = io_resp_valid & stall;
  assign T143 = T145 & T144;
  assign T144 = io_req_bits_kill ^ 1'h1;
  assign T145 = s1_valid & rdy;
  assign T146 = state == 2'h0;
  assign T147 = T149 & T148;
  assign T148 = stall ^ 1'h1;
  assign T149 = s1_valid & rdy;
  assign io_mem_acquire_valid = T150;
  assign T150 = T151 & ack_q_io_enq_ready;
  assign T151 = state == 2'h1;
  assign io_resp_bits_datablock = T152;
  assign T152 = T170 | T153;
  assign T153 = s2_tag_hit_1 ? s2_dout_1 : 128'h0;
  assign T154 = T166 ? T155 : s2_dout_1;
  assign T164 = T165 & s0_valid;
  assign T165 = T158 ^ 1'h1;
  assign T158 = FlowThroughSerializer_1_io_out_valid & T159;
  assign T159 = repl_way == 1'h1;
  assign T163 = s0_pgoff[4'hc:3'h4];
  ICache_T156 T156 (
    .CLK(clk),
    .RW0A(T158 ? T160 : T163),
    .RW0E(T164 || T158),
    .RW0W(T158),
    .RW0I(T206),
    .RW0O(T155)
  );
  assign T206 = FlowThroughSerializer_1_io_out_bits_payload_data[7'h7f:1'h0];
  assign T160 = {s2_idx, FlowThroughSerializer_1_io_cnt};
  assign T162 = T164 ? T163 : R161;
  assign T166 = T167 & s1_tag_match_1;
  assign T167 = T169 & T168;
  assign T168 = stall ^ 1'h1;
  assign T169 = s1_valid & rdy;
  assign T170 = s2_tag_hit_0 ? s2_dout_0 : 128'h0;
  assign T171 = T183 ? T172 : s2_dout_0;
  assign T181 = T182 & s0_valid;
  assign T182 = T175 ^ 1'h1;
  assign T175 = FlowThroughSerializer_1_io_out_valid & T176;
  assign T176 = repl_way == 1'h0;
  assign T180 = s0_pgoff[4'hc:3'h4];
  ICache_T156 T173 (
    .CLK(clk),
    .RW0A(T175 ? T177 : T180),
    .RW0E(T181 || T175),
    .RW0W(T175),
    .RW0I(T207),
    .RW0O(T172)
  );
  assign T207 = FlowThroughSerializer_1_io_out_bits_payload_data[7'h7f:1'h0];
  assign T177 = {s2_idx, FlowThroughSerializer_1_io_cnt};
  assign T179 = T181 ? T180 : R178;
  assign T183 = T184 & s1_tag_match_0;
  assign T184 = T186 & T185;
  assign T185 = stall ^ 1'h1;
  assign T186 = s1_valid & rdy;
  assign io_resp_bits_data = T187;
  assign T187 = T192 | T188;
  assign T188 = s2_tag_hit_1 ? s2_dout_word_1 : 32'h0;
  assign s2_dout_word_1 = T189[5'h1f:1'h0];
  assign T189 = s2_dout_1 >> T190;
  assign T190 = T191 << 3'h5;
  assign T191 = s2_offset[2'h3:2'h2];
  assign s2_offset = s2_addr[3'h5:1'h0];
  assign T192 = s2_tag_hit_0 ? s2_dout_word_0 : 32'h0;
  assign s2_dout_word_0 = T193[5'h1f:1'h0];
  assign T193 = s2_dout_0 >> T194;
  assign T194 = T195 << 3'h5;
  assign T195 = s2_offset[2'h3:2'h2];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer_1 FlowThroughSerializer_1(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_1_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_1_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_1_io_out_bits_header_src ),
       //.io_out_bits_header_dst(  )
       .io_out_bits_payload_data( FlowThroughSerializer_1_io_out_bits_payload_data ),
       //.io_out_bits_payload_client_xact_id(  )
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_uncached( FlowThroughSerializer_1_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_1_io_out_bits_payload_g_type ),
       .io_cnt( FlowThroughSerializer_1_io_cnt ),
       .io_done( FlowThroughSerializer_1_io_done )
  );
  Queue_14 ack_q(.clk(clk), .reset(reset),
       .io_enq_ready( ack_q_io_enq_ready ),
       .io_enq_valid( T208 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( FlowThroughSerializer_1_io_out_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( FlowThroughSerializer_1_io_out_bits_payload_master_xact_id ),
       .io_deq_ready( io_mem_finish_ready ),
       .io_deq_valid( ack_q_io_deq_valid ),
       .io_deq_bits_header_src( ack_q_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ack_q_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ack_q_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ack_q.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(T147) begin
      s2_addr <= s1_addr;
    end
    if(T10) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T20) begin
      R18 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T23;
    end
    if(T20) begin
      R28 <= T30;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else if(T93) begin
      vb_array <= T86;
    end else if(T85) begin
      vb_array <= T78;
    end else if(io_invalidate) begin
      vb_array <= 256'h0;
    end else if(T61) begin
      vb_array <= T43;
    end
    if(reset) begin
      R47 <= 16'h1;
    end else if(s2_miss) begin
      R47 <= T49;
    end
    if(T65) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T76) begin
      state <= 2'h0;
    end else if(T74) begin
      state <= 2'h3;
    end else if(T71) begin
      state <= 2'h2;
    end else if(T70) begin
      state <= 2'h1;
    end
    if(T97) begin
      R95 <= 1'h0;
    end
    if(T97) begin
      R100 <= T102;
    end
    if(T20) begin
      R113 <= s1_tag_match_1;
    end
    if(T132) begin
      tag_raddr <= T130;
    end
    if(T97) begin
      R136 <= s1_tag_match_0;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T141;
    end
    if(T166) begin
      s2_dout_1 <= T155;
    end
    if(T164) begin
      R161 <= T163;
    end
    if(T183) begin
      s2_dout_0 <= T172;
    end
    if(T181) begin
      R178 <= T180;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input  io_clear_hit,
    input [36:0] io_tag,
    output io_hit,
    output[7:0] io_hits,
    output[7:0] io_valid_bits,
    input  io_write,
    input [36:0] io_write_tag,
    input [2:0] io_write_addr
);

  reg [7:0] vb_array;
  wire[7:0] T47;
  wire[7:0] T0;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[7:0] T4;
  wire[7:0] T5;
  wire[7:0] T48;
  wire T6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire T11;
  wire T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[3:0] T15;
  wire[1:0] T16;
  wire hits_0;
  wire T17;
  wire[36:0] T18;
  reg [36:0] cam_tags [7:0];
  wire[36:0] T19;
  wire T20;
  wire hits_1;
  wire T21;
  wire[36:0] T22;
  wire T23;
  wire[1:0] T24;
  wire hits_2;
  wire T25;
  wire[36:0] T26;
  wire T27;
  wire hits_3;
  wire T28;
  wire[36:0] T29;
  wire T30;
  wire[3:0] T31;
  wire[1:0] T32;
  wire hits_4;
  wire T33;
  wire[36:0] T34;
  wire T35;
  wire hits_5;
  wire T36;
  wire[36:0] T37;
  wire T38;
  wire[1:0] T39;
  wire hits_6;
  wire T40;
  wire[36:0] T41;
  wire T42;
  wire hits_7;
  wire T43;
  wire[36:0] T44;
  wire T45;
  wire T46;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
`endif

  assign io_valid_bits = vb_array;
  assign T47 = reset ? 8'h0 : T0;
  assign T0 = T11 ? T9 : T1;
  assign T1 = io_clear ? 8'h0 : T2;
  assign T2 = io_write ? T3 : vb_array;
  assign T3 = T7 | T4;
  assign T4 = T48 & T5;
  assign T5 = 1'h1 << io_write_addr;
  assign T48 = T6 ? 8'hff : 8'h0;
  assign T6 = 1'h1;
  assign T7 = vb_array & T8;
  assign T8 = ~ T5;
  assign T9 = vb_array & T10;
  assign T10 = ~ io_hits;
  assign T11 = T12 & io_clear_hit;
  assign T12 = io_clear ^ 1'h1;
  assign io_hits = T13;
  assign T13 = T14;
  assign T14 = {T31, T15};
  assign T15 = {T24, T16};
  assign T16 = {hits_1, hits_0};
  assign hits_0 = T20 & T17;
  assign T17 = T18 == io_tag;
  assign T18 = cam_tags[3'h0];
  assign T20 = vb_array[1'h0:1'h0];
  assign hits_1 = T23 & T21;
  assign T21 = T22 == io_tag;
  assign T22 = cam_tags[3'h1];
  assign T23 = vb_array[1'h1:1'h1];
  assign T24 = {hits_3, hits_2};
  assign hits_2 = T27 & T25;
  assign T25 = T26 == io_tag;
  assign T26 = cam_tags[3'h2];
  assign T27 = vb_array[2'h2:2'h2];
  assign hits_3 = T30 & T28;
  assign T28 = T29 == io_tag;
  assign T29 = cam_tags[3'h3];
  assign T30 = vb_array[2'h3:2'h3];
  assign T31 = {T39, T32};
  assign T32 = {hits_5, hits_4};
  assign hits_4 = T35 & T33;
  assign T33 = T34 == io_tag;
  assign T34 = cam_tags[3'h4];
  assign T35 = vb_array[3'h4:3'h4];
  assign hits_5 = T38 & T36;
  assign T36 = T37 == io_tag;
  assign T37 = cam_tags[3'h5];
  assign T38 = vb_array[3'h5:3'h5];
  assign T39 = {hits_7, hits_6};
  assign hits_6 = T42 & T40;
  assign T40 = T41 == io_tag;
  assign T41 = cam_tags[3'h6];
  assign T42 = vb_array[3'h6:3'h6];
  assign hits_7 = T45 & T43;
  assign T43 = T44 == io_tag;
  assign T44 = cam_tags[3'h7];
  assign T45 = vb_array[3'h7:3'h7];
  assign io_hit = T46;
  assign T46 = io_hits != 8'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 8'h0;
    end else if(T11) begin
      vb_array <= T9;
    end else if(io_clear) begin
      vb_array <= 8'h0;
    end else if(io_write) begin
      vb_array <= T3;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [30:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    output io_resp_miss,
    output[7:0] io_resp_hit_idx,
    output[18:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[29:0] io_ptw_req_bits,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [18:0] io_ptw_resp_bits_ppn,
    input [5:0] io_ptw_resp_bits_perm,
    input [7:0] io_ptw_status_ip,
    input [7:0] io_ptw_status_im,
    input [6:0] io_ptw_status_zero,
    input  io_ptw_status_er,
    input  io_ptw_status_vm,
    input  io_ptw_status_s64,
    input  io_ptw_status_u64,
    input  io_ptw_status_ef,
    input  io_ptw_status_pei,
    input  io_ptw_status_ei,
    input  io_ptw_status_ps,
    input  io_ptw_status_s,
    input  io_ptw_invalidate,
    input  io_ptw_sret
);

  reg [2:0] r_refill_waddr;
  wire[2:0] T32;
  wire[2:0] repl_waddr;
  wire[2:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[2:0] T38;
  wire[2:0] T39;
  wire T40;
  reg [7:0] R41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[14:0] T46;
  wire[2:0] T47;
  wire T48;
  wire[2:0] T180;
  wire[1:0] T181;
  wire T182;
  wire[1:0] T183;
  wire[1:0] T184;
  wire[3:0] T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[1:0] T188;
  wire T189;
  wire T190;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[10:0] T58;
  wire[7:0] T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire T64;
  wire tlb_hit;
  wire[2:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[1:0] T72;
  wire T73;
  wire[2:0] T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[2:0] T196;
  wire[2:0] T197;
  wire T198;
  wire[7:0] T74;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire has_invalid_entry;
  wire T75;
  wire T2;
  wire tlb_miss;
  wire T3;
  wire bad_va;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[36:0] T212;
  reg [37:0] r_refill_tag;
  wire[37:0] T0;
  wire[37:0] lookup_tag;
  wire[37:0] T1;
  wire T213;
  wire T214;
  reg [1:0] state;
  wire[1:0] T179;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[36:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[29:0] T178;
  wire T9;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[7:0] T27;
  reg [7:0] ux_array;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T205;
  wire T76;
  wire T77;
  wire[5:0] T78;
  wire[5:0] T206;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire T83;
  wire[7:0] T84;
  reg [7:0] sx_array;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T207;
  wire T89;
  wire T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[7:0] T98;
  reg [7:0] uw_array;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T208;
  wire T103;
  wire T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire T107;
  wire[7:0] T108;
  reg [7:0] sw_array;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T209;
  wire T113;
  wire T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[7:0] T122;
  reg [7:0] ur_array;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire[7:0] T210;
  wire T127;
  wire T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire T131;
  wire[7:0] T132;
  reg [7:0] sr_array;
  wire[7:0] T133;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[7:0] T211;
  wire T137;
  wire T138;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[18:0] T141;
  wire[18:0] T142;
  wire[18:0] T143;
  wire[18:0] T144;
  wire[18:0] T145;
  reg [18:0] tag_ram [7:0];
  wire[18:0] T146;
  wire T147;
  wire[18:0] T148;
  wire[18:0] T149;
  wire[18:0] T150;
  wire T151;
  wire[18:0] T152;
  wire[18:0] T153;
  wire[18:0] T154;
  wire T155;
  wire[18:0] T156;
  wire[18:0] T157;
  wire[18:0] T158;
  wire T159;
  wire[18:0] T160;
  wire[18:0] T161;
  wire[18:0] T162;
  wire T163;
  wire[18:0] T164;
  wire[18:0] T165;
  wire[18:0] T166;
  wire T167;
  wire[18:0] T168;
  wire[18:0] T169;
  wire[18:0] T170;
  wire T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire tag_cam_io_hit;
  wire[7:0] tag_cam_io_hits;
  wire[7:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R41 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    ux_array = {1{$random}};
    sx_array = {1{$random}};
    uw_array = {1{$random}};
    sw_array = {1{$random}};
    ur_array = {1{$random}};
    sr_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
`endif

  assign T32 = T2 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T191 : T33;
  assign T33 = T34[2'h2:1'h0];
  assign T34 = {T65, T35};
  assign T35 = T40 & T36;
  assign T36 = T37 - 1'h1;
  assign T37 = 1'h1 << T38;
  assign T38 = T39 + 3'h1;
  assign T39 = T65 - T65;
  assign T40 = R41 >> T65;
  assign T42 = T64 ? T43 : R41;
  assign T43 = T53 | T44;
  assign T44 = T52 ? 8'h0 : T45;
  assign T45 = T46[3'h7:1'h0];
  assign T46 = 8'h1 << T47;
  assign T47 = {T50, T48};
  assign T48 = T180[1'h1:1'h1];
  assign T180 = {T190, T181};
  assign T181 = {T189, T182};
  assign T182 = T183[1'h1:1'h1];
  assign T183 = T188 | T184;
  assign T184 = T185[1'h1:1'h0];
  assign T185 = T187 | T186;
  assign T186 = tag_cam_io_hits[2'h3:1'h0];
  assign T187 = tag_cam_io_hits[3'h7:3'h4];
  assign T188 = T185[2'h3:2'h2];
  assign T189 = T188 != 2'h0;
  assign T190 = T187 != 4'h0;
  assign T50 = {1'h1, T51};
  assign T51 = T180[2'h2:2'h2];
  assign T52 = T180[1'h0:1'h0];
  assign T53 = T55 & T54;
  assign T54 = ~ T45;
  assign T55 = T59 | T56;
  assign T56 = T48 ? 8'h0 : T57;
  assign T57 = T58[3'h7:1'h0];
  assign T58 = 8'h1 << T50;
  assign T59 = T61 & T60;
  assign T60 = ~ T57;
  assign T61 = T63 | T62;
  assign T62 = T51 ? 8'h0 : 8'h2;
  assign T63 = R41 & 8'hfd;
  assign T64 = io_req_valid & tlb_hit;
  assign tlb_hit = io_ptw_status_vm & tag_cam_io_hit;
  assign T65 = {T72, T66};
  assign T66 = T71 & T67;
  assign T67 = T68 - 1'h1;
  assign T68 = 1'h1 << T69;
  assign T69 = T70 + 2'h1;
  assign T70 = T72 - T72;
  assign T71 = R41 >> T72;
  assign T72 = {1'h1, T73};
  assign T73 = R41[1'h1:1'h1];
  assign T191 = T204 ? 1'h0 : T192;
  assign T192 = T203 ? 1'h1 : T193;
  assign T193 = T202 ? 2'h2 : T194;
  assign T194 = T201 ? 2'h3 : T195;
  assign T195 = T200 ? 3'h4 : T196;
  assign T196 = T199 ? 3'h5 : T197;
  assign T197 = T198 ? 3'h6 : 3'h7;
  assign T198 = T74[3'h6:3'h6];
  assign T74 = ~ tag_cam_io_valid_bits;
  assign T199 = T74[3'h5:3'h5];
  assign T200 = T74[3'h4:3'h4];
  assign T201 = T74[2'h3:2'h3];
  assign T202 = T74[2'h2:2'h2];
  assign T203 = T74[1'h1:1'h1];
  assign T204 = T74[1'h0:1'h0];
  assign has_invalid_entry = T75 ^ 1'h1;
  assign T75 = tag_cam_io_valid_bits == 8'hff;
  assign T2 = T8 & tlb_miss;
  assign tlb_miss = T6 & T3;
  assign T3 = bad_va ^ 1'h1;
  assign bad_va = T5 != T4;
  assign T4 = io_req_bits_vpn[5'h1d:5'h1d];
  assign T5 = io_req_bits_vpn[5'h1e:5'h1e];
  assign T6 = io_ptw_status_vm & T7;
  assign T7 = tag_cam_io_hit ^ 1'h1;
  assign T8 = io_req_ready & io_req_valid;
  assign T212 = r_refill_tag[6'h24:1'h0];
  assign T0 = T2 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T1;
  assign T1 = {io_req_bits_asid, io_req_bits_vpn};
  assign T213 = T214 & io_ptw_resp_valid;
  assign T214 = state == 2'h2;
  assign T179 = reset ? 2'h0 : T10;
  assign T10 = io_ptw_resp_valid ? 2'h0 : T11;
  assign T11 = T20 ? 2'h3 : T12;
  assign T12 = T19 ? 2'h3 : T13;
  assign T13 = T18 ? 2'h2 : T14;
  assign T14 = T16 ? 2'h0 : T15;
  assign T15 = T2 ? 2'h1 : state;
  assign T16 = T17 & io_ptw_invalidate;
  assign T17 = state == 2'h1;
  assign T18 = T17 & io_ptw_req_ready;
  assign T19 = T18 & io_ptw_invalidate;
  assign T20 = T21 & io_ptw_invalidate;
  assign T21 = state == 2'h2;
  assign T215 = lookup_tag[6'h24:1'h0];
  assign T216 = T219 & T217;
  assign T217 = io_req_bits_instruction ? io_resp_xcpt_if : T218;
  assign T218 = io_resp_xcpt_ld & io_resp_xcpt_st;
  assign T219 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits = T178;
  assign T178 = r_refill_tag[5'h1d:1'h0];
  assign io_ptw_req_valid = T9;
  assign T9 = state == 2'h1;
  assign io_resp_xcpt_if = T22;
  assign T22 = bad_va | T23;
  assign T23 = tlb_hit & T24;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_ptw_status_s ? T83 : T26;
  assign T26 = T27 != 8'h0;
  assign T27 = ux_array & tag_cam_io_hits;
  assign T28 = io_ptw_resp_valid ? T29 : ux_array;
  assign T29 = T81 | T30;
  assign T30 = T205 & T31;
  assign T31 = 1'h1 << r_refill_waddr;
  assign T205 = T76 ? 8'hff : 8'h0;
  assign T76 = T77;
  assign T77 = T78[2'h2:2'h2];
  assign T78 = T206 & io_ptw_resp_bits_perm;
  assign T206 = T79 ? 6'h3f : 6'h0;
  assign T79 = T80;
  assign T80 = io_ptw_resp_bits_error ^ 1'h1;
  assign T81 = ux_array & T82;
  assign T82 = ~ T31;
  assign T83 = T84 != 8'h0;
  assign T84 = sx_array & tag_cam_io_hits;
  assign T85 = io_ptw_resp_valid ? T86 : sx_array;
  assign T86 = T91 | T87;
  assign T87 = T207 & T88;
  assign T88 = 1'h1 << r_refill_waddr;
  assign T207 = T89 ? 8'hff : 8'h0;
  assign T89 = T90;
  assign T90 = T78[3'h5:3'h5];
  assign T91 = sx_array & T92;
  assign T92 = ~ T88;
  assign io_resp_xcpt_st = T93;
  assign T93 = bad_va | T94;
  assign T94 = tlb_hit & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = io_ptw_status_s ? T107 : T97;
  assign T97 = T98 != 8'h0;
  assign T98 = uw_array & tag_cam_io_hits;
  assign T99 = io_ptw_resp_valid ? T100 : uw_array;
  assign T100 = T105 | T101;
  assign T101 = T208 & T102;
  assign T102 = 1'h1 << r_refill_waddr;
  assign T208 = T103 ? 8'hff : 8'h0;
  assign T103 = T104;
  assign T104 = T78[1'h1:1'h1];
  assign T105 = uw_array & T106;
  assign T106 = ~ T102;
  assign T107 = T108 != 8'h0;
  assign T108 = sw_array & tag_cam_io_hits;
  assign T109 = io_ptw_resp_valid ? T110 : sw_array;
  assign T110 = T115 | T111;
  assign T111 = T209 & T112;
  assign T112 = 1'h1 << r_refill_waddr;
  assign T209 = T113 ? 8'hff : 8'h0;
  assign T113 = T114;
  assign T114 = T78[3'h4:3'h4];
  assign T115 = sw_array & T116;
  assign T116 = ~ T112;
  assign io_resp_xcpt_ld = T117;
  assign T117 = bad_va | T118;
  assign T118 = tlb_hit & T119;
  assign T119 = T120 ^ 1'h1;
  assign T120 = io_ptw_status_s ? T131 : T121;
  assign T121 = T122 != 8'h0;
  assign T122 = ur_array & tag_cam_io_hits;
  assign T123 = io_ptw_resp_valid ? T124 : ur_array;
  assign T124 = T129 | T125;
  assign T125 = T210 & T126;
  assign T126 = 1'h1 << r_refill_waddr;
  assign T210 = T127 ? 8'hff : 8'h0;
  assign T127 = T128;
  assign T128 = T78[1'h0:1'h0];
  assign T129 = ur_array & T130;
  assign T130 = ~ T126;
  assign T131 = T132 != 8'h0;
  assign T132 = sr_array & tag_cam_io_hits;
  assign T133 = io_ptw_resp_valid ? T134 : sr_array;
  assign T134 = T139 | T135;
  assign T135 = T211 & T136;
  assign T136 = 1'h1 << r_refill_waddr;
  assign T211 = T137 ? 8'hff : 8'h0;
  assign T137 = T138;
  assign T138 = T78[2'h3:2'h3];
  assign T139 = sr_array & T140;
  assign T140 = ~ T136;
  assign io_resp_ppn = T141;
  assign T141 = T175 ? T143 : T142;
  assign T142 = io_req_bits_vpn[5'h12:1'h0];
  assign T143 = T148 | T144;
  assign T144 = T147 ? T145 : 19'h0;
  assign T145 = tag_ram[3'h7];
  assign T147 = tag_cam_io_hits[3'h7:3'h7];
  assign T148 = T152 | T149;
  assign T149 = T151 ? T150 : 19'h0;
  assign T150 = tag_ram[3'h6];
  assign T151 = tag_cam_io_hits[3'h6:3'h6];
  assign T152 = T156 | T153;
  assign T153 = T155 ? T154 : 19'h0;
  assign T154 = tag_ram[3'h5];
  assign T155 = tag_cam_io_hits[3'h5:3'h5];
  assign T156 = T160 | T157;
  assign T157 = T159 ? T158 : 19'h0;
  assign T158 = tag_ram[3'h4];
  assign T159 = tag_cam_io_hits[3'h4:3'h4];
  assign T160 = T164 | T161;
  assign T161 = T163 ? T162 : 19'h0;
  assign T162 = tag_ram[3'h3];
  assign T163 = tag_cam_io_hits[2'h3:2'h3];
  assign T164 = T168 | T165;
  assign T165 = T167 ? T166 : 19'h0;
  assign T166 = tag_ram[3'h2];
  assign T167 = tag_cam_io_hits[2'h2:2'h2];
  assign T168 = T172 | T169;
  assign T169 = T171 ? T170 : 19'h0;
  assign T170 = tag_ram[3'h1];
  assign T171 = tag_cam_io_hits[1'h1:1'h1];
  assign T172 = T174 ? T173 : 19'h0;
  assign T173 = tag_ram[3'h0];
  assign T174 = tag_cam_io_hits[1'h0:1'h0];
  assign T175 = io_ptw_status_vm & T176;
  assign T176 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T177;
  assign T177 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( io_ptw_invalidate ),
       .io_clear_hit( T216 ),
       .io_tag( T215 ),
       .io_hit( tag_cam_io_hit ),
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T213 ),
       .io_write_tag( T212 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T2) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T64) begin
      R41 <= T43;
    end
    if(T2) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T20) begin
      state <= 2'h3;
    end else if(T19) begin
      state <= 2'h3;
    end else if(T18) begin
      state <= 2'h2;
    end else if(T16) begin
      state <= 2'h0;
    end else if(T2) begin
      state <= 2'h1;
    end
    if(io_ptw_resp_valid) begin
      ux_array <= T29;
    end
    if(io_ptw_resp_valid) begin
      sx_array <= T86;
    end
    if(io_ptw_resp_valid) begin
      uw_array <= T100;
    end
    if(io_ptw_resp_valid) begin
      sw_array <= T110;
    end
    if(io_ptw_resp_valid) begin
      ur_array <= T124;
    end
    if(io_ptw_resp_valid) begin
      sr_array <= T134;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [43:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[43:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_xcpt_ma,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output[42:0] io_cpu_btb_resp_bits_target,
    output[5:0] io_cpu_btb_resp_bits_entry,
    output[6:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input [42:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_btb_update_bits_pc,
    input [42:0] io_cpu_btb_update_bits_target,
    input [42:0] io_cpu_btb_update_bits_returnAddr,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isCall,
    input  io_cpu_btb_update_bits_isReturn,
    input  io_cpu_btb_update_bits_mispredict,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    input  io_cpu_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[2:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[511:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[30:0] T38;
  wire[43:0] s1_pc;
  reg [43:0] s1_pc_;
  wire[43:0] T19;
  wire[43:0] T20;
  wire[43:0] npc;
  wire[43:0] T21;
  wire[43:0] predicted_npc;
  wire[43:0] pcp4;
  wire[42:0] T22;
  wire[43:0] pcp4_0;
  wire T23;
  wire T24;
  wire T25;
  wire[43:0] btbTarget;
  wire T26;
  reg [43:0] s2_pc;
  wire[43:0] T36;
  wire[43:0] T18;
  wire T2;
  wire T3;
  wire icmiss;
  wire T4;
  reg  s2_valid;
  wire T33;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire stall;
  wire T9;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg  s1_same_block;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire s0_same_block;
  wire T48;
  wire[43:0] T49;
  wire[43:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[12:0] T59;
  wire[43:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[42:0] T65;
  wire[43:0] T66;
  wire T67;
  wire T68;
  wire T69;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T0;
  wire T1;
  reg [6:0] s2_btb_resp_bits_bht_history;
  wire[6:0] T10;
  reg [5:0] s2_btb_resp_bits_entry;
  wire[5:0] T11;
  reg [42:0] s2_btb_resp_bits_target;
  wire[42:0] T12;
  reg  s2_btb_resp_bits_taken;
  wire T13;
  reg  s2_btb_resp_valid;
  wire T34;
  wire T14;
  reg  s2_xcpt_if;
  wire T35;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire[31:0] T37;
  wire[127:0] T27;
  wire[6:0] T28;
  wire[1:0] T29;
  wire[43:0] T30;
  wire T31;
  wire T32;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire[42:0] btb_io_resp_bits_target;
  wire[5:0] btb_io_resp_bits_entry;
  wire[6:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[2:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire icache_io_mem_acquire_bits_payload_uncached;
  wire[1:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] icache_io_mem_acquire_bits_payload_subblock;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire tlb_io_resp_miss;
  wire[18:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[29:0] tlb_io_ptw_req_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
`endif

  assign T38 = s1_pc >> 4'hd;
  assign s1_pc = s1_pc_ & 44'hffffffffffe;
  assign T19 = io_cpu_req_valid ? io_cpu_req_bits_pc : T20;
  assign T20 = T8 ? npc : s1_pc_;
  assign npc = T21;
  assign T21 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : pcp4;
  assign pcp4 = {T23, T22};
  assign T22 = pcp4_0[6'h2a:1'h0];
  assign pcp4_0 = s1_pc + 44'h4;
  assign T23 = T25 & T24;
  assign T24 = pcp4_0[6'h2a:6'h2a];
  assign T25 = s1_pc[6'h2a:6'h2a];
  assign btbTarget = {T26, btb_io_resp_bits_target};
  assign T26 = btb_io_resp_bits_target[6'h2a:6'h2a];
  assign T36 = reset ? 44'h2000 : T18;
  assign T18 = T2 ? s1_pc : s2_pc;
  assign T2 = T8 & T3;
  assign T3 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T4;
  assign T4 = icache_io_resp_valid ^ 1'h1;
  assign T33 = reset ? 1'h1 : T5;
  assign T5 = io_cpu_req_valid ? 1'h0 : T6;
  assign T6 = T8 ? T7 : s2_valid;
  assign T7 = icmiss ^ 1'h1;
  assign T8 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T9;
  assign T9 = io_cpu_resp_ready ^ 1'h1;
  assign T39 = T41 & T40;
  assign T40 = icmiss ^ 1'h1;
  assign T41 = stall ^ 1'h1;
  assign T42 = T56 & T43;
  assign T43 = s1_same_block ^ 1'h1;
  assign T44 = io_cpu_req_valid ? 1'h0 : T45;
  assign T45 = T8 ? T46 : s1_same_block;
  assign T46 = s0_same_block & T47;
  assign T47 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T51 & T48;
  assign T48 = T50 == T49;
  assign T49 = s1_pc & 44'h10;
  assign T50 = pcp4 & 44'h10;
  assign T51 = T53 & T52;
  assign T52 = btb_io_resp_bits_taken ^ 1'h1;
  assign T53 = T55 & T54;
  assign T54 = io_cpu_req_valid ^ 1'h1;
  assign T55 = icmiss ^ 1'h1;
  assign T56 = stall ^ 1'h1;
  assign T57 = T58 | icmiss;
  assign T58 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T59 = T60[4'hc:1'h0];
  assign T60 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T61 = T63 & T62;
  assign T62 = s0_same_block ^ 1'h1;
  assign T63 = stall ^ 1'h1;
  assign T64 = io_cpu_invalidate | io_cpu_ptw_invalidate;
  assign T65 = T66[6'h2a:1'h0];
  assign T66 = s1_pc & 44'hffffffffffc;
  assign T67 = T69 & T68;
  assign T68 = icmiss ^ 1'h1;
  assign T69 = stall ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = icache_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = icache_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = icache_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = icache_io_mem_finish_valid;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_payload_subblock = icache_io_mem_acquire_bits_payload_subblock;
  assign io_mem_acquire_bits_payload_a_type = icache_io_mem_acquire_bits_payload_a_type;
  assign io_mem_acquire_bits_payload_uncached = icache_io_mem_acquire_bits_payload_uncached;
  assign io_mem_acquire_bits_payload_data = icache_io_mem_acquire_bits_payload_data;
  assign io_mem_acquire_bits_payload_client_xact_id = icache_io_mem_acquire_bits_payload_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = icache_io_mem_acquire_bits_payload_addr;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cpu_ptw_req_bits = tlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T0 = T1 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T1 = T2 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T10 = T1 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T11 = T1 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T12 = T1 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T13 = T1 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T34 = reset ? 1'h0 : T14;
  assign T14 = T2 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T35 = reset ? 1'h0 : T15;
  assign T15 = T2 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_xcpt_ma = T16;
  assign T16 = T17 != 2'h0;
  assign T17 = s2_pc[1'h1:1'h0];
  assign io_cpu_resp_bits_data = T37;
  assign T37 = T27[5'h1f:1'h0];
  assign T27 = icache_io_resp_bits_datablock >> T28;
  assign T28 = T29 << 3'h5;
  assign T29 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = T30;
  assign T30 = s2_pc & 44'hffffffffffc;
  assign io_cpu_resp_valid = T31;
  assign T31 = s2_valid & T32;
  assign T32 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T67 ),
       .io_req_bits_addr( T65 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_update_valid( io_cpu_btb_update_valid ),
       .io_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_update_bits_returnAddr( io_cpu_btb_update_bits_returnAddr ),
       .io_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_update_bits_isCall( io_cpu_btb_update_bits_isCall ),
       .io_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_update_bits_mispredict( io_cpu_btb_update_bits_mispredict ),
       .io_invalidate( T64 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T61 ),
       .io_req_bits_idx( T59 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T57 ),
       .io_resp_ready( T42 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( icache_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( icache_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T39 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T38 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_resp_miss( tlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits( tlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T8) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 44'h2000;
    end else if(T2) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T8) begin
      s2_valid <= T7;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T8) begin
      s1_same_block <= T46;
    end
    if(T1) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T1) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T1) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T1) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T1) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T2) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T2) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [18:0] io_req_bits_tag,
    input [6:0] io_req_bits_idx,
    input [3:0] io_req_bits_way_en,
    input [2:0] io_req_bits_client_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output[3:0] io_data_req_bits_way_en,
    output[12:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr,
    output[2:0] io_release_bits_client_xact_id,
    output[511:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg [511:0] R2;
  wire[511:0] T3;
  wire[511:0] T4;
  wire[383:0] T5;
  wire T6;
  reg  r2_data_req_fired;
  wire T37;
  wire T7;
  reg  r1_data_req_fired;
  wire T38;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  reg  active;
  wire T39;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [2:0] cnt;
  wire[2:0] T40;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  reg [2:0] req_client_xact_id;
  wire[2:0] T26;
  wire[25:0] T27;
  wire[25:0] T28;
  reg [6:0] req_idx;
  wire[6:0] T29;
  reg [18:0] req_tag;
  wire[18:0] T30;
  wire[12:0] T31;
  wire[8:0] T32;
  wire[1:0] T33;
  reg [3:0] req_way_en;
  wire[3:0] T34;
  wire fire;
  wire T35;
  wire T36;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    R2 = {16{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    cnt = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_idx = {1{$random}};
    req_tag = {1{$random}};
    req_way_en = {1{$random}};
  end
`endif

  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_data = R2;
  assign T3 = T6 ? T4 : R2;
  assign T4 = {io_data_resp, T5};
  assign T5 = R2[9'h1ff:8'h80];
  assign T6 = active & r2_data_req_fired;
  assign T37 = reset ? 1'h0 : T7;
  assign T7 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T38 = reset ? 1'h0 : T8;
  assign T8 = T10 ? 1'h1 : T9;
  assign T9 = active ? 1'h0 : r1_data_req_fired;
  assign T10 = active & T11;
  assign T11 = T13 & T12;
  assign T12 = io_meta_read_ready & io_meta_read_valid;
  assign T13 = io_data_req_ready & io_data_req_valid;
  assign T39 = reset ? 1'h0 : T14;
  assign T14 = T1 ? 1'h1 : T15;
  assign T15 = T17 ? T16 : active;
  assign T16 = io_release_ready ^ 1'h1;
  assign T17 = active & T18;
  assign T18 = T23 & T19;
  assign T19 = cnt == 3'h4;
  assign T40 = reset ? 3'h0 : T20;
  assign T20 = T1 ? 3'h0 : T21;
  assign T21 = T10 ? T22 : cnt;
  assign T22 = cnt + 3'h1;
  assign T23 = T25 & T24;
  assign T24 = r2_data_req_fired ^ 1'h1;
  assign T25 = r1_data_req_fired ^ 1'h1;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T26 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr = T27;
  assign T27 = T28;
  assign T28 = {req_tag, req_idx};
  assign T29 = T1 ? io_req_bits_idx : req_idx;
  assign T30 = T1 ? io_req_bits_tag : req_tag;
  assign io_release_valid = T17;
  assign io_data_req_bits_addr = T31;
  assign T31 = T32 << 3'h4;
  assign T32 = {req_idx, T33};
  assign T33 = cnt[1'h1:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T34 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T35;
  assign T35 = cnt < 3'h4;
  assign io_meta_read_bits_tag = req_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T36;
  assign T36 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T6) begin
      R2 <= T4;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T10) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T17) begin
      active <= T16;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else if(T1) begin
      cnt <= 3'h0;
    end else if(T10) begin
      cnt <= T22;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_idx <= io_req_bits_idx;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr,
    input [1:0] io_req_bits_p_type,
    input [2:0] io_req_bits_client_xact_id,
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr,
    output[2:0] io_rep_bits_client_xact_id,
    output[511:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[2:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    input [3:0] io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_line_state_state
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  reg [1:0] req_p_type;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [3:0] state;
  wire[3:0] T91;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  reg [1:0] line_state_state;
  wire[1:0] T29;
  wire T30;
  wire hit;
  reg [3:0] way_en;
  wire[3:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  reg [2:0] req_client_xact_id;
  wire[2:0] T50;
  wire[6:0] T92;
  reg [25:0] req_addr;
  wire[25:0] T51;
  wire[18:0] T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[18:0] T61;
  wire[6:0] T93;
  wire T62;
  wire[18:0] T63;
  wire[6:0] T94;
  wire T64;
  wire[2:0] T65;
  wire[2:0] T66;
  wire[2:0] T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire[511:0] T82;
  wire[2:0] T83;
  wire[25:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_p_type = {1{$random}};
    state = {1{$random}};
    line_state_state = {1{$random}};
    way_en = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr = {1{$random}};
  end
`endif

  assign io_wb_req_bits_r_type = T0;
  assign T0 = T47 ? T41 : T1;
  assign T1 = T40 ? 3'h4 : T2;
  assign T2 = T39 ? 3'h5 : T3;
  assign T3 = T4 ? 3'h6 : 3'h4;
  assign T4 = req_p_type == 2'h2;
  assign T5 = T6 ? io_req_bits_p_type : req_p_type;
  assign T6 = T7 & io_req_valid;
  assign T7 = state == 4'h1;
  assign T91 = reset ? 4'h1 : T8;
  assign T8 = T38 ? 4'h1 : T9;
  assign T9 = T6 ? 4'h2 : T10;
  assign T10 = T36 ? 4'h3 : T11;
  assign T11 = T35 ? 4'h4 : T12;
  assign T12 = T33 ? 4'h2 : T13;
  assign T13 = T32 ? 4'h5 : T14;
  assign T14 = T30 ? T27 : T15;
  assign T15 = T25 ? 4'h1 : T16;
  assign T16 = T23 ? 4'h7 : T17;
  assign T17 = T21 ? 4'h8 : T18;
  assign T18 = T19 ? 4'h1 : state;
  assign T19 = T20 & io_meta_write_ready;
  assign T20 = state == 4'h8;
  assign T21 = T22 & io_wb_req_ready;
  assign T22 = state == 4'h7;
  assign T23 = T24 & io_wb_req_ready;
  assign T24 = state == 4'h6;
  assign T25 = T26 & io_rep_ready;
  assign T26 = state == 4'h5;
  assign T27 = T28 ? 4'h6 : 4'h8;
  assign T28 = line_state_state == 2'h2;
  assign T29 = T32 ? io_line_state_state : line_state_state;
  assign T30 = T25 & hit;
  assign hit = way_en != 4'h0;
  assign T31 = T32 ? io_way_en : way_en;
  assign T32 = state == 4'h4;
  assign T33 = T32 & T34;
  assign T34 = io_mshr_rdy ^ 1'h1;
  assign T35 = state == 4'h3;
  assign T36 = T37 & io_meta_read_ready;
  assign T37 = state == 4'h2;
  assign T38 = state == 4'h0;
  assign T39 = req_p_type == 2'h1;
  assign T40 = req_p_type == 2'h0;
  assign T41 = T46 ? 3'h1 : T42;
  assign T42 = T45 ? 3'h2 : T43;
  assign T43 = T44 ? 3'h3 : 3'h1;
  assign T44 = req_p_type == 2'h2;
  assign T45 = req_p_type == 2'h1;
  assign T46 = req_p_type == 2'h0;
  assign T47 = T48 == 2'h2;
  assign T48 = hit ? line_state_state : T49;
  assign T49 = 2'h0;
  assign io_wb_req_bits_client_xact_id = req_client_xact_id;
  assign T50 = T6 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_wb_req_bits_way_en = way_en;
  assign io_wb_req_bits_idx = T92;
  assign T92 = req_addr[3'h6:1'h0];
  assign T51 = T6 ? io_req_bits_addr : req_addr;
  assign io_wb_req_bits_tag = T52;
  assign T52 = req_addr >> 3'h7;
  assign io_wb_req_valid = T53;
  assign T53 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T54;
  assign T54 = T55;
  assign T55 = T60 ? 2'h0 : T56;
  assign T56 = T59 ? 2'h1 : T57;
  assign T57 = T58 ? line_state_state : line_state_state;
  assign T58 = req_p_type == 2'h2;
  assign T59 = req_p_type == 2'h1;
  assign T60 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T61;
  assign T61 = req_addr >> 3'h7;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T93;
  assign T93 = req_addr[3'h6:1'h0];
  assign io_meta_write_valid = T62;
  assign T62 = state == 4'h8;
  assign io_meta_read_bits_tag = T63;
  assign T63 = req_addr >> 3'h7;
  assign io_meta_read_bits_idx = T94;
  assign T94 = req_addr[3'h6:1'h0];
  assign io_meta_read_valid = T64;
  assign T64 = state == 4'h2;
  assign io_rep_bits_r_type = T65;
  assign T65 = T66;
  assign T66 = T79 ? T73 : T67;
  assign T67 = T72 ? 3'h4 : T68;
  assign T68 = T71 ? 3'h5 : T69;
  assign T69 = T70 ? 3'h6 : 3'h4;
  assign T70 = req_p_type == 2'h2;
  assign T71 = req_p_type == 2'h1;
  assign T72 = req_p_type == 2'h0;
  assign T73 = T78 ? 3'h1 : T74;
  assign T74 = T77 ? 3'h2 : T75;
  assign T75 = T76 ? 3'h3 : 3'h1;
  assign T76 = req_p_type == 2'h2;
  assign T77 = req_p_type == 2'h1;
  assign T78 = req_p_type == 2'h0;
  assign T79 = T80 == 2'h2;
  assign T80 = hit ? line_state_state : T81;
  assign T81 = 2'h0;
  assign io_rep_bits_data = T82;
  assign T82 = 512'h0;
  assign io_rep_bits_client_xact_id = T83;
  assign T83 = req_client_xact_id;
  assign io_rep_bits_addr = T84;
  assign T84 = req_addr;
  assign io_rep_valid = T85;
  assign T85 = T89 & T86;
  assign T86 = T87 ^ 1'h1;
  assign T87 = hit & T88;
  assign T88 = line_state_state == 2'h2;
  assign T89 = state == 4'h5;
  assign io_req_ready = T90;
  assign T90 = state == 4'h1;

  always @(posedge clk) begin
    if(T6) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(reset) begin
      state <= 4'h1;
    end else if(T38) begin
      state <= 4'h1;
    end else if(T6) begin
      state <= 4'h2;
    end else if(T36) begin
      state <= 4'h3;
    end else if(T35) begin
      state <= 4'h4;
    end else if(T33) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T30) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T23) begin
      state <= 4'h7;
    end else if(T21) begin
      state <= 4'h8;
    end else if(T19) begin
      state <= 4'h1;
    end
    if(T32) begin
      line_state_state <= io_line_state_state;
    end
    if(T32) begin
      way_en <= io_way_en;
    end
    if(T6) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T6) begin
      req_addr <= io_req_bits_addr;
    end
  end
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    input [18:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input [18:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[18:0] io_out_bits_tag,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[18:0] T2;
  wire T3;
  wire[6:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T2;
  assign T2 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T3 = T0;
  assign io_out_bits_idx = T4;
  assign T4 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [18:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [18:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[18:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[1:0] T2;
  wire T3;
  wire[18:0] T4;
  wire[3:0] T5;
  wire[6:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T2;
  assign T2 = T3 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T3 = T0;
  assign io_out_bits_data_tag = T4;
  assign T4 = T3 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T5;
  assign T5 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T6;
  assign T6 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [2:0] io_in_1_bits_client_xact_id,
    input [511:0] io_in_1_bits_data,
    input  io_in_1_bits_uncached,
    input [1:0] io_in_1_bits_a_type,
    input [511:0] io_in_1_bits_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [2:0] io_in_0_bits_client_xact_id,
    input [511:0] io_in_0_bits_data,
    input  io_in_0_bits_uncached,
    input [1:0] io_in_0_bits_a_type,
    input [511:0] io_in_0_bits_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[2:0] io_out_bits_client_xact_id,
    output[511:0] io_out_bits_data,
    output io_out_bits_uncached,
    output[1:0] io_out_bits_a_type,
    output[511:0] io_out_bits_subblock,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[511:0] T2;
  wire T3;
  wire[1:0] T4;
  wire T5;
  wire[511:0] T6;
  wire[2:0] T7;
  wire[25:0] T8;
  wire T9;
  wire T10;
  wire T11;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_subblock = T2;
  assign T2 = T3 ? io_in_1_bits_subblock : io_in_0_bits_subblock;
  assign T3 = T0;
  assign io_out_bits_a_type = T4;
  assign T4 = T3 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_uncached = T5;
  assign T5 = T3 ? io_in_1_bits_uncached : io_in_0_bits_uncached;
  assign io_out_bits_data = T6;
  assign T6 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T7;
  assign T7 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T8;
  assign T8 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T9;
  assign T9 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_9(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_payload_master_xact_id = T2;
  assign T2 = T3 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T3 = T0;
  assign io_out_bits_header_dst = T4;
  assign T4 = T3 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T5;
  assign T5 = T3 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T6;
  assign T6 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [18:0] io_in_1_bits_tag,
    input [6:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [2:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [18:0] io_in_0_bits_tag,
    input [6:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [2:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[18:0] io_out_bits_tag,
    output[6:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[2:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[3:0] T5;
  wire[6:0] T6;
  wire[18:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_client_xact_id = T4;
  assign T4 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_way_en = T5;
  assign T5 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T6;
  assign T6 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_bits_tag = T7;
  assign T7 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_valid = T8;
  assign T8 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_10(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [8:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [8:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[2:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[8:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[4:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[8:0] T5;
  wire[43:0] T6;
  wire T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T2;
  assign T2 = T3 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T3 = T0;
  assign io_out_bits_cmd = T4;
  assign T4 = T3 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T5;
  assign T5 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T6;
  assign T6 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T7;
  assign T7 = T3 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T8;
  assign T8 = T3 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T9;
  assign T9 = T3 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T10;
  assign T10 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_11(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits = T2;
  assign T2 = T3 ? io_in_1_bits : io_in_0_bits;
  assign T3 = T0;
  assign io_out_valid = T4;
  assign T4 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_17(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [8:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[8:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T29;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T30;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T31;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[67:0] T11;
  reg [67:0] ram [15:0];
  wire[67:0] T12;
  wire[67:0] T13;
  wire[67:0] T14;
  wire[62:0] T15;
  wire[9:0] T16;
  wire[52:0] T17;
  wire[4:0] T18;
  wire[3:0] T19;
  wire[4:0] T20;
  wire[8:0] T21;
  wire[43:0] T22;
  wire T23;
  wire[2:0] T24;
  wire T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T29 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T30 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T31 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_cmd, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_addr, io_enq_bits_tag};
  assign T18 = {io_enq_bits_kill, T19};
  assign T19 = {io_enq_bits_typ, io_enq_bits_phys};
  assign io_deq_bits_cmd = T20;
  assign T20 = T11[4'h9:3'h5];
  assign io_deq_bits_tag = T21;
  assign T21 = T11[5'h12:4'ha];
  assign io_deq_bits_addr = T22;
  assign T22 = T11[6'h3e:5'h13];
  assign io_deq_bits_phys = T23;
  assign T23 = T11[6'h3f:6'h3f];
  assign io_deq_bits_typ = T24;
  assign T24 = T11[7'h42:7'h40];
  assign io_deq_bits_kill = T25;
  assign T25 = T11[7'h43:7'h43];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input [4:0] io_req_bits_sdq_id,
    output io_idx_match,
    output[18:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[2:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output io_mem_req_bits_uncached,
    output[1:0] io_mem_req_bits_a_type,
    output[511:0] io_mem_req_bits_subblock,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[2:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T190;
  wire can_finish;
  wire T77;
  reg [3:0] state;
  wire[3:0] T186;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire refill_done;
  wire T28;
  reg [1:0] refill_count;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire reply;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T78;
  wire T79;
  wire T80;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire wb_done;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T82;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire sec_rdy;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire idx_match;
  wire[6:0] T70;
  wire[6:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T71;
  wire T208;
  wire T0;
  wire T1;
  wire T2;
  reg [1:0] meta_hazard;
  wire[1:0] T185;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg [3:0] req_way_en;
  wire[3:0] T72;
  reg [18:0] req_old_meta_tag;
  wire[18:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire[4:0] T81;
  wire[43:0] T187;
  wire[31:0] T83;
  wire[31:0] T84;
  wire[12:0] T85;
  wire[5:0] T86;
  wire T87;
  wire T88;
  wire[1:0] T89;
  reg [1:0] line_state_state;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T93;
  wire[1:0] T94;
  wire T95;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[1:0] meta_on_flush_state;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[12:0] T109;
  wire[8:0] T110;
  wire[511:0] T111;
  wire[1:0] T112;
  reg [1:0] acquire_type;
  wire[1:0] T113;
  wire[1:0] T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire[1:0] T188;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[511:0] T140;
  wire[2:0] T141;
  wire[25:0] T142;
  wire[25:0] T143;
  wire[25:0] T144;
  wire T145;
  wire T146;
  wire[18:0] T189;
  wire[30:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire T184;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[2:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[8:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T190 = io_mem_finish_ready & can_finish;
  assign can_finish = T78 | T77;
  assign T77 = state == 4'h5;
  assign T186 = reset ? 4'h0 : T10;
  assign T10 = T64 ? T62 : T11;
  assign T11 = T60 ? 4'h4 : T12;
  assign T12 = T42 ? 4'h6 : T13;
  assign T13 = T41 ? 4'h2 : T14;
  assign T14 = T39 ? 4'h3 : T15;
  assign T15 = T37 ? 4'h4 : T16;
  assign T16 = T36 ? 4'h5 : T17;
  assign T17 = T27 ? 4'h6 : T18;
  assign T18 = T25 ? 4'h7 : T19;
  assign T19 = T24 ? 4'h8 : T20;
  assign T20 = T21 ? 4'h0 : state;
  assign T21 = T23 & T22;
  assign T22 = rpq_io_deq_valid ^ 1'h1;
  assign T23 = state == 4'h8;
  assign T24 = state == 4'h7;
  assign T25 = T26 & io_meta_write_ready;
  assign T26 = state == 4'h6;
  assign T27 = T35 & refill_done;
  assign refill_done = reply & T28;
  assign T28 = refill_count == 2'h3;
  assign T29 = T33 ? 2'h0 : T30;
  assign T30 = T32 ? T31 : refill_count;
  assign T31 = refill_count + 2'h1;
  assign T32 = T35 & reply;
  assign T33 = io_req_pri_val & io_req_pri_rdy;
  assign reply = io_mem_grant_valid & T34;
  assign T34 = io_mem_grant_bits_payload_client_xact_id == 3'h0;
  assign T35 = state == 4'h5;
  assign T36 = io_mem_req_ready & io_mem_req_valid;
  assign T37 = T38 & io_meta_write_ready;
  assign T38 = state == 4'h3;
  assign T39 = T40 & reply;
  assign T40 = state == 4'h2;
  assign T41 = io_wb_req_ready & io_wb_req_valid;
  assign T42 = T59 & T43;
  assign T43 = T48 ? T47 : T44;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T46 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T47 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T33 & io_req_bits_tag_match;
  assign T60 = T59 & T61;
  assign T61 = T43 ^ 1'h1;
  assign T62 = T63 ? 4'h1 : 4'h3;
  assign T63 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T64 = T33 & T65;
  assign T65 = io_req_bits_tag_match ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = state == 4'h4;
  assign T80 = state == 4'h0;
  assign T191 = T194 & T192;
  assign T192 = io_mem_grant_bits_payload_uncached | T193;
  assign T193 = io_mem_grant_bits_payload_g_type != 2'h0;
  assign T194 = wb_done | refill_done;
  assign wb_done = reply & T195;
  assign T195 = state == 4'h2;
  assign T196 = T82 ? 1'h0 : T197;
  assign T197 = T199 | T198;
  assign T198 = state == 4'h0;
  assign T199 = io_replay_ready & T200;
  assign T200 = state == 4'h8;
  assign T82 = io_meta_read_ready ^ 1'h1;
  assign T201 = T206 & T202;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T205 | T204;
  assign T204 = io_req_bits_cmd == 5'h3;
  assign T205 = io_req_bits_cmd == 5'h2;
  assign T206 = T208 | T207;
  assign T207 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T151;
  assign T151 = T179 | T152;
  assign T152 = T176 & T153;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T168 | T155;
  assign T155 = T157 & T156;
  assign T156 = io_mem_req_bits_a_type != 2'h1;
  assign T157 = T159 | T158;
  assign T158 = io_req_bits_cmd == 5'h6;
  assign T159 = T161 | T160;
  assign T160 = io_req_bits_cmd == 5'h3;
  assign T161 = T165 | T162;
  assign T162 = T164 | T163;
  assign T163 = io_req_bits_cmd == 5'h4;
  assign T164 = io_req_bits_cmd[2'h3:2'h3];
  assign T165 = T167 | T166;
  assign T166 = io_req_bits_cmd == 5'h7;
  assign T167 = io_req_bits_cmd == 5'h1;
  assign T168 = T169 & io_mem_req_bits_uncached;
  assign T169 = T173 | T170;
  assign T170 = T172 | T171;
  assign T171 = io_req_bits_cmd == 5'h4;
  assign T172 = io_req_bits_cmd[2'h3:2'h3];
  assign T173 = T175 | T174;
  assign T174 = io_req_bits_cmd == 5'h6;
  assign T175 = io_req_bits_cmd == 5'h0;
  assign T176 = T178 | T177;
  assign T177 = state == 4'h5;
  assign T178 = state == 4'h4;
  assign T179 = T181 | T180;
  assign T180 = state == 4'h3;
  assign T181 = T183 | T182;
  assign T182 = state == 4'h2;
  assign T183 = state == 4'h1;
  assign idx_match = req_idx == T70;
  assign T70 = io_req_bits_addr[4'hc:3'h6];
  assign req_idx = req_addr[4'hc:3'h6];
  assign T71 = T33 ? io_req_bits_addr : req_addr;
  assign T208 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T0;
  assign T0 = T69 | T1;
  assign T1 = T8 & T2;
  assign T2 = meta_hazard == 2'h0;
  assign T185 = reset ? 2'h0 : T3;
  assign T3 = T7 ? 2'h1 : T4;
  assign T4 = T6 ? T5 : meta_hazard;
  assign T5 = meta_hazard + 2'h1;
  assign T6 = meta_hazard != 2'h0;
  assign T7 = io_meta_write_ready & io_meta_write_valid;
  assign T8 = T66 & T9;
  assign T9 = state != 4'h3;
  assign T66 = T68 & T67;
  assign T67 = state != 4'h2;
  assign T68 = state != 4'h1;
  assign T69 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_client_xact_id = 3'h0;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T72 = T33 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T73 = T33 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T74;
  assign T74 = T75 & ackq_io_enq_ready;
  assign T75 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T76;
  assign T76 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T81;
  assign T81 = T82 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T187;
  assign T187 = {12'h0, T83};
  assign T83 = T84;
  assign T84 = {io_tag, T85};
  assign T85 = {req_idx, T86};
  assign T86 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T87;
  assign T87 = T88 & rpq_io_deq_valid;
  assign T88 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T89;
  assign T89 = T104 ? meta_on_flush_state : line_state_state;
  assign T90 = T42 ? meta_on_hit_state : T91;
  assign T91 = T33 ? meta_on_flush_state : T92;
  assign T92 = T32 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T93;
  assign T93 = io_mem_grant_bits_payload_uncached ? 2'h0 : T94;
  assign T94 = T95 ? 2'h1 : 2'h2;
  assign T95 = io_mem_grant_bits_payload_g_type == 2'h1;
  assign meta_on_hit_state = T96;
  assign T96 = T97 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign T97 = T101 | T98;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h4;
  assign T100 = io_req_bits_cmd[2'h3:2'h3];
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h7;
  assign T103 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T104 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T105;
  assign T105 = T107 | T106;
  assign T106 = state == 4'h3;
  assign T107 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T108;
  assign T108 = state == 4'h8;
  assign io_mem_resp_addr = T109;
  assign T109 = T110 << 3'h4;
  assign T110 = {req_idx, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_subblock = T111;
  assign T111 = 512'h0;
  assign io_mem_req_bits_a_type = T112;
  assign T112 = acquire_type;
  assign T113 = T33 ? T188 : T114;
  assign T114 = T127 ? T115 : acquire_type;
  assign T115 = T116 ? 2'h1 : io_mem_req_bits_a_type;
  assign T116 = T118 | T117;
  assign T117 = io_req_bits_cmd == 5'h6;
  assign T118 = T120 | T119;
  assign T119 = io_req_bits_cmd == 5'h3;
  assign T120 = T124 | T121;
  assign T121 = T123 | T122;
  assign T122 = io_req_bits_cmd == 5'h4;
  assign T123 = io_req_bits_cmd[2'h3:2'h3];
  assign T124 = T126 | T125;
  assign T125 = io_req_bits_cmd == 5'h7;
  assign T126 = io_req_bits_cmd == 5'h1;
  assign T127 = io_req_sec_val & io_req_sec_rdy;
  assign T188 = {1'h0, T128};
  assign T128 = T130 | T129;
  assign T129 = io_req_bits_cmd == 5'h6;
  assign T130 = T132 | T131;
  assign T131 = io_req_bits_cmd == 5'h3;
  assign T132 = T136 | T133;
  assign T133 = T135 | T134;
  assign T134 = io_req_bits_cmd == 5'h4;
  assign T135 = io_req_bits_cmd[2'h3:2'h3];
  assign T136 = T138 | T137;
  assign T137 = io_req_bits_cmd == 5'h7;
  assign T138 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_uncached = T139;
  assign T139 = 1'h0;
  assign io_mem_req_bits_data = T140;
  assign T140 = 512'h0;
  assign io_mem_req_bits_client_xact_id = T141;
  assign T141 = 3'h0;
  assign io_mem_req_bits_addr = T142;
  assign T142 = T143;
  assign T143 = T144;
  assign T144 = {io_tag, req_idx};
  assign io_mem_req_valid = T145;
  assign T145 = T146 & ackq_io_enq_ready;
  assign T146 = state == 4'h4;
  assign io_tag = T189;
  assign T189 = T147[5'h12:1'h0];
  assign T147 = req_addr >> 4'hd;
  assign io_idx_match = T148;
  assign T148 = T149 & idx_match;
  assign T149 = state != 4'h0;
  assign io_req_sec_rdy = T150;
  assign T150 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T184;
  assign T184 = state == 4'h0;
  Queue_17 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T201 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T196 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_14 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T191 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T190 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T64) begin
      state <= T62;
    end else if(T60) begin
      state <= 4'h4;
    end else if(T42) begin
      state <= 4'h6;
    end else if(T41) begin
      state <= 4'h2;
    end else if(T39) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= 4'h5;
    end else if(T27) begin
      state <= 4'h6;
    end else if(T25) begin
      state <= 4'h7;
    end else if(T24) begin
      state <= 4'h8;
    end else if(T21) begin
      state <= 4'h0;
    end
    if(T33) begin
      refill_count <= 2'h0;
    end else if(T32) begin
      refill_count <= T31;
    end
    if(T33) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T7) begin
      meta_hazard <= 2'h1;
    end else if(T6) begin
      meta_hazard <= T5;
    end
    if(T33) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T33) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T42) begin
      line_state_state <= meta_on_hit_state;
    end else if(T33) begin
      line_state_state <= meta_on_flush_state;
    end else if(T32) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T33) begin
      acquire_type <= T188;
    end else if(T127) begin
      acquire_type <= T115;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input [4:0] io_req_bits_sdq_id,
    output io_idx_match,
    output[18:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[2:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output io_mem_req_bits_uncached,
    output[1:0] io_mem_req_bits_a_type,
    output[511:0] io_mem_req_bits_subblock,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[2:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T190;
  wire can_finish;
  wire T77;
  reg [3:0] state;
  wire[3:0] T186;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire refill_done;
  wire T28;
  reg [1:0] refill_count;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire reply;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T78;
  wire T79;
  wire T80;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire wb_done;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T82;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire sec_rdy;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire idx_match;
  wire[6:0] T70;
  wire[6:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T71;
  wire T208;
  wire T0;
  wire T1;
  wire T2;
  reg [1:0] meta_hazard;
  wire[1:0] T185;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg [3:0] req_way_en;
  wire[3:0] T72;
  reg [18:0] req_old_meta_tag;
  wire[18:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire[4:0] T81;
  wire[43:0] T187;
  wire[31:0] T83;
  wire[31:0] T84;
  wire[12:0] T85;
  wire[5:0] T86;
  wire T87;
  wire T88;
  wire[1:0] T89;
  reg [1:0] line_state_state;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T93;
  wire[1:0] T94;
  wire T95;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[1:0] meta_on_flush_state;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[12:0] T109;
  wire[8:0] T110;
  wire[511:0] T111;
  wire[1:0] T112;
  reg [1:0] acquire_type;
  wire[1:0] T113;
  wire[1:0] T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire[1:0] T188;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[511:0] T140;
  wire[2:0] T141;
  wire[25:0] T142;
  wire[25:0] T143;
  wire[25:0] T144;
  wire T145;
  wire T146;
  wire[18:0] T189;
  wire[30:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire T184;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[2:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[8:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T190 = io_mem_finish_ready & can_finish;
  assign can_finish = T78 | T77;
  assign T77 = state == 4'h5;
  assign T186 = reset ? 4'h0 : T10;
  assign T10 = T64 ? T62 : T11;
  assign T11 = T60 ? 4'h4 : T12;
  assign T12 = T42 ? 4'h6 : T13;
  assign T13 = T41 ? 4'h2 : T14;
  assign T14 = T39 ? 4'h3 : T15;
  assign T15 = T37 ? 4'h4 : T16;
  assign T16 = T36 ? 4'h5 : T17;
  assign T17 = T27 ? 4'h6 : T18;
  assign T18 = T25 ? 4'h7 : T19;
  assign T19 = T24 ? 4'h8 : T20;
  assign T20 = T21 ? 4'h0 : state;
  assign T21 = T23 & T22;
  assign T22 = rpq_io_deq_valid ^ 1'h1;
  assign T23 = state == 4'h8;
  assign T24 = state == 4'h7;
  assign T25 = T26 & io_meta_write_ready;
  assign T26 = state == 4'h6;
  assign T27 = T35 & refill_done;
  assign refill_done = reply & T28;
  assign T28 = refill_count == 2'h3;
  assign T29 = T33 ? 2'h0 : T30;
  assign T30 = T32 ? T31 : refill_count;
  assign T31 = refill_count + 2'h1;
  assign T32 = T35 & reply;
  assign T33 = io_req_pri_val & io_req_pri_rdy;
  assign reply = io_mem_grant_valid & T34;
  assign T34 = io_mem_grant_bits_payload_client_xact_id == 3'h1;
  assign T35 = state == 4'h5;
  assign T36 = io_mem_req_ready & io_mem_req_valid;
  assign T37 = T38 & io_meta_write_ready;
  assign T38 = state == 4'h3;
  assign T39 = T40 & reply;
  assign T40 = state == 4'h2;
  assign T41 = io_wb_req_ready & io_wb_req_valid;
  assign T42 = T59 & T43;
  assign T43 = T48 ? T47 : T44;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T46 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T47 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T33 & io_req_bits_tag_match;
  assign T60 = T59 & T61;
  assign T61 = T43 ^ 1'h1;
  assign T62 = T63 ? 4'h1 : 4'h3;
  assign T63 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T64 = T33 & T65;
  assign T65 = io_req_bits_tag_match ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = state == 4'h4;
  assign T80 = state == 4'h0;
  assign T191 = T194 & T192;
  assign T192 = io_mem_grant_bits_payload_uncached | T193;
  assign T193 = io_mem_grant_bits_payload_g_type != 2'h0;
  assign T194 = wb_done | refill_done;
  assign wb_done = reply & T195;
  assign T195 = state == 4'h2;
  assign T196 = T82 ? 1'h0 : T197;
  assign T197 = T199 | T198;
  assign T198 = state == 4'h0;
  assign T199 = io_replay_ready & T200;
  assign T200 = state == 4'h8;
  assign T82 = io_meta_read_ready ^ 1'h1;
  assign T201 = T206 & T202;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T205 | T204;
  assign T204 = io_req_bits_cmd == 5'h3;
  assign T205 = io_req_bits_cmd == 5'h2;
  assign T206 = T208 | T207;
  assign T207 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T151;
  assign T151 = T179 | T152;
  assign T152 = T176 & T153;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T168 | T155;
  assign T155 = T157 & T156;
  assign T156 = io_mem_req_bits_a_type != 2'h1;
  assign T157 = T159 | T158;
  assign T158 = io_req_bits_cmd == 5'h6;
  assign T159 = T161 | T160;
  assign T160 = io_req_bits_cmd == 5'h3;
  assign T161 = T165 | T162;
  assign T162 = T164 | T163;
  assign T163 = io_req_bits_cmd == 5'h4;
  assign T164 = io_req_bits_cmd[2'h3:2'h3];
  assign T165 = T167 | T166;
  assign T166 = io_req_bits_cmd == 5'h7;
  assign T167 = io_req_bits_cmd == 5'h1;
  assign T168 = T169 & io_mem_req_bits_uncached;
  assign T169 = T173 | T170;
  assign T170 = T172 | T171;
  assign T171 = io_req_bits_cmd == 5'h4;
  assign T172 = io_req_bits_cmd[2'h3:2'h3];
  assign T173 = T175 | T174;
  assign T174 = io_req_bits_cmd == 5'h6;
  assign T175 = io_req_bits_cmd == 5'h0;
  assign T176 = T178 | T177;
  assign T177 = state == 4'h5;
  assign T178 = state == 4'h4;
  assign T179 = T181 | T180;
  assign T180 = state == 4'h3;
  assign T181 = T183 | T182;
  assign T182 = state == 4'h2;
  assign T183 = state == 4'h1;
  assign idx_match = req_idx == T70;
  assign T70 = io_req_bits_addr[4'hc:3'h6];
  assign req_idx = req_addr[4'hc:3'h6];
  assign T71 = T33 ? io_req_bits_addr : req_addr;
  assign T208 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T0;
  assign T0 = T69 | T1;
  assign T1 = T8 & T2;
  assign T2 = meta_hazard == 2'h0;
  assign T185 = reset ? 2'h0 : T3;
  assign T3 = T7 ? 2'h1 : T4;
  assign T4 = T6 ? T5 : meta_hazard;
  assign T5 = meta_hazard + 2'h1;
  assign T6 = meta_hazard != 2'h0;
  assign T7 = io_meta_write_ready & io_meta_write_valid;
  assign T8 = T66 & T9;
  assign T9 = state != 4'h3;
  assign T66 = T68 & T67;
  assign T67 = state != 4'h2;
  assign T68 = state != 4'h1;
  assign T69 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_client_xact_id = 3'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T72 = T33 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T73 = T33 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T74;
  assign T74 = T75 & ackq_io_enq_ready;
  assign T75 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T76;
  assign T76 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T81;
  assign T81 = T82 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T187;
  assign T187 = {12'h0, T83};
  assign T83 = T84;
  assign T84 = {io_tag, T85};
  assign T85 = {req_idx, T86};
  assign T86 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T87;
  assign T87 = T88 & rpq_io_deq_valid;
  assign T88 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T89;
  assign T89 = T104 ? meta_on_flush_state : line_state_state;
  assign T90 = T42 ? meta_on_hit_state : T91;
  assign T91 = T33 ? meta_on_flush_state : T92;
  assign T92 = T32 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T93;
  assign T93 = io_mem_grant_bits_payload_uncached ? 2'h0 : T94;
  assign T94 = T95 ? 2'h1 : 2'h2;
  assign T95 = io_mem_grant_bits_payload_g_type == 2'h1;
  assign meta_on_hit_state = T96;
  assign T96 = T97 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign T97 = T101 | T98;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h4;
  assign T100 = io_req_bits_cmd[2'h3:2'h3];
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h7;
  assign T103 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T104 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T105;
  assign T105 = T107 | T106;
  assign T106 = state == 4'h3;
  assign T107 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T108;
  assign T108 = state == 4'h8;
  assign io_mem_resp_addr = T109;
  assign T109 = T110 << 3'h4;
  assign T110 = {req_idx, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_subblock = T111;
  assign T111 = 512'h0;
  assign io_mem_req_bits_a_type = T112;
  assign T112 = acquire_type;
  assign T113 = T33 ? T188 : T114;
  assign T114 = T127 ? T115 : acquire_type;
  assign T115 = T116 ? 2'h1 : io_mem_req_bits_a_type;
  assign T116 = T118 | T117;
  assign T117 = io_req_bits_cmd == 5'h6;
  assign T118 = T120 | T119;
  assign T119 = io_req_bits_cmd == 5'h3;
  assign T120 = T124 | T121;
  assign T121 = T123 | T122;
  assign T122 = io_req_bits_cmd == 5'h4;
  assign T123 = io_req_bits_cmd[2'h3:2'h3];
  assign T124 = T126 | T125;
  assign T125 = io_req_bits_cmd == 5'h7;
  assign T126 = io_req_bits_cmd == 5'h1;
  assign T127 = io_req_sec_val & io_req_sec_rdy;
  assign T188 = {1'h0, T128};
  assign T128 = T130 | T129;
  assign T129 = io_req_bits_cmd == 5'h6;
  assign T130 = T132 | T131;
  assign T131 = io_req_bits_cmd == 5'h3;
  assign T132 = T136 | T133;
  assign T133 = T135 | T134;
  assign T134 = io_req_bits_cmd == 5'h4;
  assign T135 = io_req_bits_cmd[2'h3:2'h3];
  assign T136 = T138 | T137;
  assign T137 = io_req_bits_cmd == 5'h7;
  assign T138 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_uncached = T139;
  assign T139 = 1'h0;
  assign io_mem_req_bits_data = T140;
  assign T140 = 512'h0;
  assign io_mem_req_bits_client_xact_id = T141;
  assign T141 = 3'h1;
  assign io_mem_req_bits_addr = T142;
  assign T142 = T143;
  assign T143 = T144;
  assign T144 = {io_tag, req_idx};
  assign io_mem_req_valid = T145;
  assign T145 = T146 & ackq_io_enq_ready;
  assign T146 = state == 4'h4;
  assign io_tag = T189;
  assign T189 = T147[5'h12:1'h0];
  assign T147 = req_addr >> 4'hd;
  assign io_idx_match = T148;
  assign T148 = T149 & idx_match;
  assign T149 = state != 4'h0;
  assign io_req_sec_rdy = T150;
  assign T150 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T184;
  assign T184 = state == 4'h0;
  Queue_17 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T201 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T196 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_14 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T191 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T190 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T64) begin
      state <= T62;
    end else if(T60) begin
      state <= 4'h4;
    end else if(T42) begin
      state <= 4'h6;
    end else if(T41) begin
      state <= 4'h2;
    end else if(T39) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= 4'h5;
    end else if(T27) begin
      state <= 4'h6;
    end else if(T25) begin
      state <= 4'h7;
    end else if(T24) begin
      state <= 4'h8;
    end else if(T21) begin
      state <= 4'h0;
    end
    if(T33) begin
      refill_count <= 2'h0;
    end else if(T32) begin
      refill_count <= T31;
    end
    if(T33) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T7) begin
      meta_hazard <= 2'h1;
    end else if(T6) begin
      meta_hazard <= T5;
    end
    if(T33) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T33) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T42) begin
      line_state_state <= meta_on_hit_state;
    end else if(T33) begin
      line_state_state <= meta_on_flush_state;
    end else if(T32) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T33) begin
      acquire_type <= T188;
    end else if(T127) begin
      acquire_type <= T115;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input [63:0] io_req_bits_data,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[2:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output io_mem_req_bits_uncached,
    output[1:0] io_mem_req_bits_a_type,
    output[511:0] io_mem_req_bits_subblock,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[63:0] io_replay_bits_data,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[2:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire[4:0] T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire[4:0] T95;
  wire[4:0] T96;
  wire[4:0] T97;
  wire[4:0] T98;
  wire[4:0] T99;
  wire[4:0] T100;
  wire[4:0] T101;
  wire[4:0] T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire[4:0] T106;
  wire[4:0] T107;
  wire T108;
  wire[16:0] T21;
  wire[16:0] T22;
  reg [16:0] sdq_val;
  wire[16:0] T109;
  wire[31:0] T110;
  wire[31:0] T23;
  wire[31:0] T111;
  wire[31:0] T24;
  wire[31:0] T112;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T113;
  wire sdq_enq;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire[16:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire[16:0] T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire[16:0] T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire[16:0] T41;
  wire[16:0] T42;
  wire[16:0] T43;
  wire T44;
  wire[16:0] T45;
  wire[16:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[31:0] T114;
  wire[16:0] T66;
  wire[16:0] T115;
  wire free_sdq;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[31:0] T75;
  wire[31:0] T116;
  wire T76;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T134;
  wire tag_match;
  wire[30:0] T88;
  wire[30:0] T133;
  wire[18:0] T89;
  wire[18:0] T90;
  wire[18:0] tagList_1;
  wire idxMatch_1;
  wire[18:0] T91;
  wire[18:0] tagList_0;
  wire idxMatch_0;
  wire T135;
  wire sdq_rdy;
  wire T85;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire idx_match;
  wire T140;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[63:0] T8;
  reg [63:0] sdq [16:0];
  wire[63:0] T9;
  wire T10;
  wire T11;
  wire[4:0] T12;
  reg [4:0] R77;
  wire[4:0] T78;
  wire[127:0] T79;
  wire[127:0] memRespMux_0_data;
  wire[127:0] memRespMux_1_data;
  wire T80;
  wire T132;
  wire[1:0] T81;
  wire[1:0] memRespMux_0_wmask;
  wire[1:0] memRespMux_1_wmask;
  wire[12:0] T82;
  wire[12:0] memRespMux_0_addr;
  wire[12:0] memRespMux_1_addr;
  wire[3:0] T83;
  wire[3:0] memRespMux_0_way_en;
  wire[3:0] memRespMux_1_way_en;
  wire T84;
  wire T86;
  wire pri_rdy;
  wire T87;
  wire sec_rdy;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[6:0] meta_read_arb_io_out_bits_idx;
  wire[18:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[6:0] meta_write_arb_io_out_bits_idx;
  wire[3:0] meta_write_arb_io_out_bits_way_en;
  wire[18:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr;
  wire[2:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[511:0] mem_req_arb_io_out_bits_data;
  wire mem_req_arb_io_out_bits_uncached;
  wire[1:0] mem_req_arb_io_out_bits_a_type;
  wire[511:0] mem_req_arb_io_out_bits_subblock;
  wire mem_finish_arb_io_in_1_ready;
  wire mem_finish_arb_io_in_0_ready;
  wire mem_finish_arb_io_out_valid;
  wire[1:0] mem_finish_arb_io_out_bits_header_src;
  wire[1:0] mem_finish_arb_io_out_bits_header_dst;
  wire[2:0] mem_finish_arb_io_out_bits_payload_master_xact_id;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[18:0] wb_req_arb_io_out_bits_tag;
  wire[6:0] wb_req_arb_io_out_bits_idx;
  wire[3:0] wb_req_arb_io_out_bits_way_en;
  wire[2:0] wb_req_arb_io_out_bits_client_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire replay_arb_io_out_bits_kill;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_phys;
  wire[43:0] replay_arb_io_out_bits_addr;
  wire[8:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire MSHR_0_io_req_pri_rdy;
  wire MSHR_0_io_req_sec_rdy;
  wire MSHR_0_io_idx_match;
  wire[18:0] MSHR_0_io_tag;
  wire MSHR_0_io_mem_req_valid;
  wire[25:0] MSHR_0_io_mem_req_bits_addr;
  wire[2:0] MSHR_0_io_mem_req_bits_client_xact_id;
  wire[511:0] MSHR_0_io_mem_req_bits_data;
  wire MSHR_0_io_mem_req_bits_uncached;
  wire[1:0] MSHR_0_io_mem_req_bits_a_type;
  wire[511:0] MSHR_0_io_mem_req_bits_subblock;
  wire[3:0] MSHR_0_io_mem_resp_way_en;
  wire[12:0] MSHR_0_io_mem_resp_addr;
  wire[1:0] MSHR_0_io_mem_resp_wmask;
  wire[127:0] MSHR_0_io_mem_resp_data;
  wire MSHR_0_io_meta_read_valid;
  wire[6:0] MSHR_0_io_meta_read_bits_idx;
  wire[18:0] MSHR_0_io_meta_read_bits_tag;
  wire MSHR_0_io_meta_write_valid;
  wire[6:0] MSHR_0_io_meta_write_bits_idx;
  wire[3:0] MSHR_0_io_meta_write_bits_way_en;
  wire[18:0] MSHR_0_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_0_io_meta_write_bits_data_coh_state;
  wire MSHR_0_io_replay_valid;
  wire MSHR_0_io_replay_bits_kill;
  wire[2:0] MSHR_0_io_replay_bits_typ;
  wire MSHR_0_io_replay_bits_phys;
  wire[43:0] MSHR_0_io_replay_bits_addr;
  wire[8:0] MSHR_0_io_replay_bits_tag;
  wire[4:0] MSHR_0_io_replay_bits_cmd;
  wire[4:0] MSHR_0_io_replay_bits_sdq_id;
  wire MSHR_0_io_mem_finish_valid;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_dst;
  wire[2:0] MSHR_0_io_mem_finish_bits_payload_master_xact_id;
  wire MSHR_0_io_wb_req_valid;
  wire[18:0] MSHR_0_io_wb_req_bits_tag;
  wire[6:0] MSHR_0_io_wb_req_bits_idx;
  wire[3:0] MSHR_0_io_wb_req_bits_way_en;
  wire[2:0] MSHR_0_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_0_io_wb_req_bits_r_type;
  wire MSHR_0_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[18:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr;
  wire[2:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[511:0] MSHR_1_io_mem_req_bits_data;
  wire MSHR_1_io_mem_req_bits_uncached;
  wire[1:0] MSHR_1_io_mem_req_bits_a_type;
  wire[511:0] MSHR_1_io_mem_req_bits_subblock;
  wire[3:0] MSHR_1_io_mem_resp_way_en;
  wire[12:0] MSHR_1_io_mem_resp_addr;
  wire[1:0] MSHR_1_io_mem_resp_wmask;
  wire[127:0] MSHR_1_io_mem_resp_data;
  wire MSHR_1_io_meta_read_valid;
  wire[6:0] MSHR_1_io_meta_read_bits_idx;
  wire[18:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[6:0] MSHR_1_io_meta_write_bits_idx;
  wire[3:0] MSHR_1_io_meta_write_bits_way_en;
  wire[18:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire MSHR_1_io_replay_bits_kill;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_phys;
  wire[43:0] MSHR_1_io_replay_bits_addr;
  wire[8:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_mem_finish_valid;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_dst;
  wire[2:0] MSHR_1_io_mem_finish_bits_payload_master_xact_id;
  wire MSHR_1_io_wb_req_valid;
  wire[18:0] MSHR_1_io_wb_req_bits_tag;
  wire[6:0] MSHR_1_io_wb_req_bits_idx;
  wire[3:0] MSHR_1_io_wb_req_bits_way_en;
  wire[2:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R77 = {1{$random}};
  end
`endif

  assign T92 = T131 ? 1'h0 : T93;
  assign T93 = T130 ? 1'h1 : T94;
  assign T94 = T129 ? 2'h2 : T95;
  assign T95 = T128 ? 2'h3 : T96;
  assign T96 = T127 ? 3'h4 : T97;
  assign T97 = T126 ? 3'h5 : T98;
  assign T98 = T125 ? 3'h6 : T99;
  assign T99 = T124 ? 3'h7 : T100;
  assign T100 = T123 ? 4'h8 : T101;
  assign T101 = T122 ? 4'h9 : T102;
  assign T102 = T121 ? 4'ha : T103;
  assign T103 = T120 ? 4'hb : T104;
  assign T104 = T119 ? 4'hc : T105;
  assign T105 = T118 ? 4'hd : T106;
  assign T106 = T117 ? 4'he : T107;
  assign T107 = T108 ? 4'hf : 5'h10;
  assign T108 = T21[4'hf:4'hf];
  assign T21 = ~ T22;
  assign T22 = sdq_val[5'h10:1'h0];
  assign T109 = T110[5'h10:1'h0];
  assign T110 = reset ? 32'h0 : T23;
  assign T23 = T76 ? T24 : T111;
  assign T111 = {15'h0, sdq_val};
  assign T24 = T63 | T112;
  assign T112 = {15'h0, T25};
  assign T25 = T27 & T26;
  assign T26 = 17'h0 - T113;
  assign T113 = {16'h0, sdq_enq};
  assign sdq_enq = T20 & T13;
  assign T13 = T17 | T14;
  assign T14 = T16 | T15;
  assign T15 = io_req_bits_cmd == 5'h4;
  assign T16 = io_req_bits_cmd[2'h3:2'h3];
  assign T17 = T19 | T18;
  assign T18 = io_req_bits_cmd == 5'h7;
  assign T19 = io_req_bits_cmd == 5'h1;
  assign T20 = io_req_valid & io_req_ready;
  assign T27 = T62 ? 17'h1 : T28;
  assign T28 = T61 ? 17'h2 : T29;
  assign T29 = T60 ? 17'h4 : T30;
  assign T30 = T59 ? 17'h8 : T31;
  assign T31 = T58 ? 17'h10 : T32;
  assign T32 = T57 ? 17'h20 : T33;
  assign T33 = T56 ? 17'h40 : T34;
  assign T34 = T55 ? 17'h80 : T35;
  assign T35 = T54 ? 17'h100 : T36;
  assign T36 = T53 ? 17'h200 : T37;
  assign T37 = T52 ? 17'h400 : T38;
  assign T38 = T51 ? 17'h800 : T39;
  assign T39 = T50 ? 17'h1000 : T40;
  assign T40 = T49 ? 17'h2000 : T41;
  assign T41 = T48 ? 17'h4000 : T42;
  assign T42 = T47 ? 17'h8000 : T43;
  assign T43 = T44 ? 17'h10000 : 17'h0;
  assign T44 = T45[5'h10:5'h10];
  assign T45 = ~ T46;
  assign T46 = sdq_val[5'h10:1'h0];
  assign T47 = T45[4'hf:4'hf];
  assign T48 = T45[4'he:4'he];
  assign T49 = T45[4'hd:4'hd];
  assign T50 = T45[4'hc:4'hc];
  assign T51 = T45[4'hb:4'hb];
  assign T52 = T45[4'ha:4'ha];
  assign T53 = T45[4'h9:4'h9];
  assign T54 = T45[4'h8:4'h8];
  assign T55 = T45[3'h7:3'h7];
  assign T56 = T45[3'h6:3'h6];
  assign T57 = T45[3'h5:3'h5];
  assign T58 = T45[3'h4:3'h4];
  assign T59 = T45[2'h3:2'h3];
  assign T60 = T45[2'h2:2'h2];
  assign T61 = T45[1'h1:1'h1];
  assign T62 = T45[1'h0:1'h0];
  assign T63 = T116 & T64;
  assign T64 = ~ T65;
  assign T65 = T75 & T114;
  assign T114 = {15'h0, T66};
  assign T66 = 17'h0 - T115;
  assign T115 = {16'h0, free_sdq};
  assign free_sdq = T74 & T67;
  assign T67 = T71 | T68;
  assign T68 = T70 | T69;
  assign T69 = io_replay_bits_cmd == 5'h4;
  assign T70 = io_replay_bits_cmd[2'h3:2'h3];
  assign T71 = T73 | T72;
  assign T72 = io_replay_bits_cmd == 5'h7;
  assign T73 = io_replay_bits_cmd == 5'h1;
  assign T74 = io_replay_ready & io_replay_valid;
  assign T75 = 1'h1 << replay_arb_io_out_bits_sdq_id;
  assign T116 = {15'h0, sdq_val};
  assign T76 = io_replay_valid | sdq_enq;
  assign T117 = T21[4'he:4'he];
  assign T118 = T21[4'hd:4'hd];
  assign T119 = T21[4'hc:4'hc];
  assign T120 = T21[4'hb:4'hb];
  assign T121 = T21[4'ha:4'ha];
  assign T122 = T21[4'h9:4'h9];
  assign T123 = T21[4'h8:4'h8];
  assign T124 = T21[3'h7:3'h7];
  assign T125 = T21[3'h6:3'h6];
  assign T126 = T21[3'h5:3'h5];
  assign T127 = T21[3'h4:3'h4];
  assign T128 = T21[2'h3:2'h3];
  assign T129 = T21[2'h2:2'h2];
  assign T130 = T21[1'h1:1'h1];
  assign T131 = T21[1'h0:1'h0];
  assign T134 = T135 & tag_match;
  assign tag_match = T133 == T88;
  assign T88 = io_req_bits_addr >> 4'hd;
  assign T133 = {12'h0, T89};
  assign T89 = T91 | T90;
  assign T90 = idxMatch_1 ? tagList_1 : 19'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T91 = idxMatch_0 ? tagList_0 : 19'h0;
  assign tagList_0 = MSHR_0_io_tag;
  assign idxMatch_0 = MSHR_0_io_idx_match;
  assign T135 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T85 ^ 1'h1;
  assign T85 = sdq_val == 17'h1ffff;
  assign T136 = T137 & tag_match;
  assign T137 = io_req_valid & sdq_rdy;
  assign T138 = T140 & T139;
  assign T139 = idx_match ^ 1'h1;
  assign idx_match = MSHR_0_io_idx_match | MSHR_1_io_idx_match;
  assign T140 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T0;
  assign T0 = T3 ? 1'h0 : T1;
  assign T1 = T2 == 1'h0;
  assign T2 = MSHR_0_io_req_pri_rdy ^ 1'h1;
  assign T3 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T4;
  assign T4 = T7 ? 1'h0 : T5;
  assign T5 = T6 == 1'h0;
  assign T6 = MSHR_0_io_probe_rdy ^ 1'h1;
  assign T7 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_idx = wb_req_arb_io_out_bits_idx;
  assign io_wb_req_bits_tag = wb_req_arb_io_out_bits_tag;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_mem_finish_bits_payload_master_xact_id = mem_finish_arb_io_out_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mem_finish_arb_io_out_bits_header_dst;
  assign io_mem_finish_bits_header_src = mem_finish_arb_io_out_bits_header_src;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_replay_bits_data = T8;
  assign T8 = sdq[R77];
  assign T10 = sdq_enq & T11;
  assign T11 = T12 < 5'h11;
  assign T12 = T92[3'h4:1'h0];
  assign T78 = free_sdq ? replay_arb_io_out_bits_sdq_id : R77;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_mem_resp_data = T79;
  assign T79 = T80 ? memRespMux_1_data : memRespMux_0_data;
  assign memRespMux_0_data = MSHR_0_io_mem_resp_data;
  assign memRespMux_1_data = MSHR_1_io_mem_resp_data;
  assign T80 = T132;
  assign T132 = io_mem_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_mem_resp_wmask = T81;
  assign T81 = T80 ? memRespMux_1_wmask : memRespMux_0_wmask;
  assign memRespMux_0_wmask = MSHR_0_io_mem_resp_wmask;
  assign memRespMux_1_wmask = MSHR_1_io_mem_resp_wmask;
  assign io_mem_resp_addr = T82;
  assign T82 = T80 ? memRespMux_1_addr : memRespMux_0_addr;
  assign memRespMux_0_addr = MSHR_0_io_mem_resp_addr;
  assign memRespMux_1_addr = MSHR_1_io_mem_resp_addr;
  assign io_mem_resp_way_en = T83;
  assign T83 = T80 ? memRespMux_1_way_en : memRespMux_0_way_en;
  assign memRespMux_0_way_en = MSHR_0_io_mem_resp_way_en;
  assign memRespMux_1_way_en = MSHR_1_io_mem_resp_way_en;
  assign io_mem_req_bits_subblock = mem_req_arb_io_out_bits_subblock;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_uncached = mem_req_arb_io_out_bits_uncached;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr = mem_req_arb_io_out_bits_addr;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T84;
  assign T84 = T86 & sdq_rdy;
  assign T86 = idx_match ? T87 : pri_rdy;
  assign pri_rdy = MSHR_0_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T87 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_0_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_7 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  Arbiter_8 mem_req_arb(
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_in_1_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_in_1_bits_uncached( MSHR_1_io_mem_req_bits_uncached ),
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_in_1_bits_subblock( MSHR_1_io_mem_req_bits_subblock ),
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_req_valid ),
       .io_in_0_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       .io_in_0_bits_data( MSHR_0_io_mem_req_bits_data ),
       .io_in_0_bits_uncached( MSHR_0_io_mem_req_bits_uncached ),
       .io_in_0_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       .io_in_0_bits_subblock( MSHR_0_io_mem_req_bits_subblock ),
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr( mem_req_arb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_uncached( mem_req_arb_io_out_bits_uncached ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_subblock( mem_req_arb_io_out_bits_subblock )
       //.io_chosen(  )
  );
  Arbiter_9 mem_finish_arb(
       .io_in_1_ready( mem_finish_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_finish_valid ),
       .io_in_1_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_in_1_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( mem_finish_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_finish_valid ),
       .io_in_0_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_in_0_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_mem_finish_ready ),
       .io_out_valid( mem_finish_arb_io_out_valid ),
       .io_out_bits_header_src( mem_finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( mem_finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( mem_finish_arb_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  Arbiter_5 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_wb_req_valid ),
       .io_in_0_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_tag( wb_req_arb_io_out_bits_tag ),
       .io_out_bits_idx( wb_req_arb_io_out_bits_idx ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  Arbiter_10 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_replay_valid ),
       .io_in_0_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_in_0_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_in_0_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_in_0_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_in_0_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_in_0_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_11 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T138 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  MSHR_0 MSHR_0(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_0_io_req_pri_rdy ),
       .io_req_sec_val( T136 ),
       .io_req_sec_rdy( MSHR_0_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_bits_sdq_id( T92 ),
       .io_idx_match( MSHR_0_io_idx_match ),
       .io_tag( MSHR_0_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_0_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( MSHR_0_io_mem_req_bits_data ),
       .io_mem_req_bits_uncached( MSHR_0_io_mem_req_bits_uncached ),
       .io_mem_req_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       .io_mem_req_bits_subblock( MSHR_0_io_mem_req_bits_subblock ),
       .io_mem_resp_way_en( MSHR_0_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_0_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_0_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_0_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_0_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_0_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_0_io_replay_valid ),
       .io_replay_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_0_ready ),
       .io_mem_finish_valid( MSHR_0_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_0_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_0_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_0.io_mem_resp_wmask = {1{$random}};
    assign MSHR_0.io_mem_resp_data = {4{$random}};
  `endif
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T134 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_bits_sdq_id( T92 ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_mem_req_bits_uncached( MSHR_1_io_mem_req_bits_uncached ),
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_mem_req_bits_subblock( MSHR_1_io_mem_req_bits_subblock ),
       .io_mem_resp_way_en( MSHR_1_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_1_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_1_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_1_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_1_ready ),
       .io_mem_finish_valid( MSHR_1_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_1.io_mem_resp_wmask = {1{$random}};
    assign MSHR_1.io_mem_resp_data = {4{$random}};
  `endif

  always @(posedge clk) begin
    sdq_val <= T109;
    if (T10)
      sdq[T92] <= io_req_bits_data;
    if(free_sdq) begin
      R77 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [6:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [6:0] io_write_bits_idx,
    input [3:0] io_write_bits_way_en,
    input [18:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[18:0] io_resp_3_tag,
    output[1:0] io_resp_3_coh_state,
    output[18:0] io_resp_2_tag,
    output[1:0] io_resp_2_coh_state,
    output[18:0] io_resp_1_tag,
    output[1:0] io_resp_1_coh_state,
    output[18:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[20:0] T1;
  wire[83:0] tags;
  wire[83:0] T2;
  wire[83:0] T3;
  wire[83:0] T4;
  wire[41:0] T5;
  wire[20:0] T6;
  wire[20:0] T40;
  wire T7;
  wire[3:0] wmask;
  wire rst;
  reg [7:0] rst_cnt;
  wire[7:0] T41;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[20:0] T10;
  wire[20:0] T42;
  wire T11;
  wire[41:0] T12;
  wire[20:0] T13;
  wire[20:0] T43;
  wire T14;
  wire[20:0] T15;
  wire[20:0] T44;
  wire T16;
  wire[83:0] T17;
  wire[41:0] T18;
  wire[20:0] wdata;
  wire[20:0] T19;
  wire[1:0] T20;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T21;
  wire[18:0] T22;
  wire[18:0] rstVal_tag;
  wire T23;
  wire[6:0] T45;
  wire[7:0] waddr;
  wire[7:0] T46;
  reg [6:0] R24;
  wire[6:0] T25;
  wire[18:0] T26;
  wire[1:0] T27;
  wire[20:0] T28;
  wire[18:0] T29;
  wire[1:0] T30;
  wire[20:0] T31;
  wire[18:0] T32;
  wire[1:0] T33;
  wire[20:0] T34;
  wire[18:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R24 = {1{$random}};
  end
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = tags[5'h14:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T45),
    .W0E(T23),
    .W0I(T17),
    .W0M(T3),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(tags)
  );
  assign T3 = T4;
  assign T4 = {T12, T5};
  assign T5 = {T10, T6};
  assign T6 = 21'h0 - T40;
  assign T40 = {20'h0, T7};
  assign T7 = wmask[1'h0:1'h0];
  assign wmask = rst ? 4'hf : io_write_bits_way_en;
  assign rst = rst_cnt < 8'h80;
  assign T41 = reset ? 8'h0 : T8;
  assign T8 = rst ? T9 : rst_cnt;
  assign T9 = rst_cnt + 8'h1;
  assign T10 = 21'h0 - T42;
  assign T42 = {20'h0, T11};
  assign T11 = wmask[1'h1:1'h1];
  assign T12 = {T15, T13};
  assign T13 = 21'h0 - T43;
  assign T43 = {20'h0, T14};
  assign T14 = wmask[2'h2:2'h2];
  assign T15 = 21'h0 - T44;
  assign T44 = {20'h0, T16};
  assign T16 = wmask[2'h3:2'h3];
  assign T17 = {T18, T18};
  assign T18 = {wdata, wdata};
  assign wdata = T19;
  assign T19 = {T22, T20};
  assign T20 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T21;
  assign T21 = 2'h0;
  assign T22 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 19'h0;
  assign T23 = rst | io_write_valid;
  assign T45 = waddr[3'h6:1'h0];
  assign waddr = rst ? rst_cnt : T46;
  assign T46 = {1'h0, io_write_bits_idx};
  assign T25 = io_read_valid ? io_read_bits_idx : R24;
  assign io_resp_0_tag = T26;
  assign T26 = T1[5'h14:2'h2];
  assign io_resp_1_coh_state = T27;
  assign T27 = T28[1'h1:1'h0];
  assign T28 = tags[6'h29:5'h15];
  assign io_resp_1_tag = T29;
  assign T29 = T28[5'h14:2'h2];
  assign io_resp_2_coh_state = T30;
  assign T30 = T31[1'h1:1'h0];
  assign T31 = tags[6'h3e:6'h2a];
  assign io_resp_2_tag = T32;
  assign T32 = T31[5'h14:2'h2];
  assign io_resp_3_coh_state = T33;
  assign T33 = T34[1'h1:1'h0];
  assign T34 = tags[7'h53:6'h3f];
  assign io_resp_3_tag = T35;
  assign T35 = T34[5'h14:2'h2];
  assign io_write_ready = T36;
  assign T36 = rst ^ 1'h1;
  assign io_read_ready = T37;
  assign T37 = T39 & T38;
  assign T38 = io_write_valid ^ 1'h1;
  assign T39 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 8'h0;
    end else if(rst) begin
      rst_cnt <= T9;
    end
    if(io_read_valid) begin
      R24 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [6:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [6:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [6:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[6:0] T5;
  wire[6:0] T6;
  wire[6:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T5;
  assign T5 = T13 ? io_in_4_bits_idx : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_valid = T14;
  assign T14 = T21 ? io_in_4_valid : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26 ^ 1'h1;
  assign T26 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T30 | io_in_2_valid;
  assign T30 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T34 | io_in_3_valid;
  assign T34 = T35 | io_in_2_valid;
  assign T35 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input [3:0] io_read_bits_way_en,
    input [12:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input [3:0] io_write_bits_way_en,
    input [12:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_3,
    output[127:0] io_resp_2,
    output[127:0] io_resp_1,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[127:0] T4;
  wire[127:0] T5;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire[8:0] raddr;
  wire[127:0] T7;
  wire[127:0] T8;
  wire[127:0] T9;
  wire[63:0] T10;
  wire[63:0] T116;
  wire T11;
  wire[1:0] T12;
  wire[63:0] T13;
  wire[63:0] T117;
  wire T14;
  wire[127:0] T15;
  wire[63:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[8:0] waddr;
  reg [8:0] R21;
  wire[8:0] T22;
  wire T26;
  wire T27;
  reg [12:0] R28;
  wire[12:0] T29;
  wire[63:0] T30;
  wire[127:0] T31;
  wire[127:0] T32;
  wire T49;
  wire T50;
  wire[127:0] T34;
  wire[127:0] T35;
  wire[127:0] T36;
  wire[63:0] T37;
  wire[63:0] T118;
  wire T38;
  wire[63:0] T39;
  wire[63:0] T119;
  wire T40;
  wire[127:0] T41;
  wire[63:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg [8:0] R47;
  wire[8:0] T48;
  wire[127:0] T51;
  wire[127:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire T55;
  wire T56;
  wire[63:0] T57;
  wire[127:0] T58;
  wire[127:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[127:0] T62;
  wire[127:0] T63;
  wire T81;
  wire T82;
  wire[1:0] T83;
  wire[127:0] T65;
  wire[127:0] T66;
  wire[127:0] T67;
  wire[63:0] T68;
  wire[63:0] T120;
  wire T69;
  wire[1:0] T70;
  wire[63:0] T71;
  wire[63:0] T121;
  wire T72;
  wire[127:0] T73;
  wire[63:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [8:0] R79;
  wire[8:0] T80;
  wire T84;
  wire T85;
  reg [12:0] R86;
  wire[12:0] T87;
  wire[63:0] T88;
  wire[127:0] T89;
  wire[127:0] T90;
  wire T107;
  wire T108;
  wire[127:0] T92;
  wire[127:0] T93;
  wire[127:0] T94;
  wire[63:0] T95;
  wire[63:0] T122;
  wire T96;
  wire[63:0] T97;
  wire[63:0] T123;
  wire T98;
  wire[127:0] T99;
  wire[63:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg [8:0] R105;
  wire[8:0] T106;
  wire[127:0] T109;
  wire[127:0] T110;
  wire[63:0] T111;
  wire[63:0] T112;
  wire T113;
  wire T114;
  wire[63:0] T115;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R21 = {1{$random}};
    R28 = {1{$random}};
    R47 = {1{$random}};
    R79 = {1{$random}};
    R86 = {1{$random}};
    R105 = {1{$random}};
  end
`endif

  assign io_resp_0 = T0;
  assign T0 = T1;
  assign T1 = {T30, T2};
  assign T2 = T26 ? T30 : T3;
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = T5;
  assign T23 = T24 & io_read_valid;
  assign T24 = T25 != 2'h0;
  assign T25 = io_read_bits_way_en[1'h1:1'h0];
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T6 T6 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T17),
    .W0I(T15),
    .W0M(T8),
    .R1A(raddr),
    .R1E(T23),
    .R1O(T5)
  );
  assign T8 = T9;
  assign T9 = {T13, T10};
  assign T10 = 64'h0 - T116;
  assign T116 = {63'h0, T11};
  assign T11 = T12[1'h0:1'h0];
  assign T12 = io_write_bits_way_en[1'h1:1'h0];
  assign T13 = 64'h0 - T117;
  assign T117 = {63'h0, T14};
  assign T14 = T12[1'h1:1'h1];
  assign T15 = {T16, T16};
  assign T16 = io_write_bits_data[6'h3f:1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_write_bits_wmask[1'h0:1'h0];
  assign T19 = T20 & io_write_valid;
  assign T20 = T12 != 2'h0;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T22 = T23 ? raddr : R21;
  assign T26 = T27;
  assign T27 = R28[2'h3:2'h3];
  assign T29 = io_read_valid ? io_read_bits_addr : R28;
  assign T30 = T31[6'h3f:1'h0];
  assign T31 = T32;
  assign T49 = T50 & io_read_valid;
  assign T50 = T25 != 2'h0;
  DataArray_T6 T33 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T43),
    .W0I(T41),
    .W0M(T35),
    .R1A(raddr),
    .R1E(T49),
    .R1O(T32)
  );
  assign T35 = T36;
  assign T36 = {T39, T37};
  assign T37 = 64'h0 - T118;
  assign T118 = {63'h0, T38};
  assign T38 = T12[1'h0:1'h0];
  assign T39 = 64'h0 - T119;
  assign T119 = {63'h0, T40};
  assign T40 = T12[1'h1:1'h1];
  assign T41 = {T42, T42};
  assign T42 = io_write_bits_data[7'h7f:7'h40];
  assign T43 = T45 & T44;
  assign T44 = io_write_bits_wmask[1'h1:1'h1];
  assign T45 = T46 & io_write_valid;
  assign T46 = T12 != 2'h0;
  assign T48 = T49 ? raddr : R47;
  assign io_resp_1 = T51;
  assign T51 = T52;
  assign T52 = {T57, T53};
  assign T53 = T55 ? T57 : T54;
  assign T54 = T4[7'h7f:7'h40];
  assign T55 = T56;
  assign T56 = R28[2'h3:2'h3];
  assign T57 = T31[7'h7f:7'h40];
  assign io_resp_2 = T58;
  assign T58 = T59;
  assign T59 = {T88, T60};
  assign T60 = T84 ? T88 : T61;
  assign T61 = T62[6'h3f:1'h0];
  assign T62 = T63;
  assign T81 = T82 & io_read_valid;
  assign T82 = T83 != 2'h0;
  assign T83 = io_read_bits_way_en[2'h3:2'h2];
  DataArray_T6 T64 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T75),
    .W0I(T73),
    .W0M(T66),
    .R1A(raddr),
    .R1E(T81),
    .R1O(T63)
  );
  assign T66 = T67;
  assign T67 = {T71, T68};
  assign T68 = 64'h0 - T120;
  assign T120 = {63'h0, T69};
  assign T69 = T70[1'h0:1'h0];
  assign T70 = io_write_bits_way_en[2'h3:2'h2];
  assign T71 = 64'h0 - T121;
  assign T121 = {63'h0, T72};
  assign T72 = T70[1'h1:1'h1];
  assign T73 = {T74, T74};
  assign T74 = io_write_bits_data[6'h3f:1'h0];
  assign T75 = T77 & T76;
  assign T76 = io_write_bits_wmask[1'h0:1'h0];
  assign T77 = T78 & io_write_valid;
  assign T78 = T70 != 2'h0;
  assign T80 = T81 ? raddr : R79;
  assign T84 = T85;
  assign T85 = R86[2'h3:2'h3];
  assign T87 = io_read_valid ? io_read_bits_addr : R86;
  assign T88 = T89[6'h3f:1'h0];
  assign T89 = T90;
  assign T107 = T108 & io_read_valid;
  assign T108 = T83 != 2'h0;
  DataArray_T6 T91 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T101),
    .W0I(T99),
    .W0M(T93),
    .R1A(raddr),
    .R1E(T107),
    .R1O(T90)
  );
  assign T93 = T94;
  assign T94 = {T97, T95};
  assign T95 = 64'h0 - T122;
  assign T122 = {63'h0, T96};
  assign T96 = T70[1'h0:1'h0];
  assign T97 = 64'h0 - T123;
  assign T123 = {63'h0, T98};
  assign T98 = T70[1'h1:1'h1];
  assign T99 = {T100, T100};
  assign T100 = io_write_bits_data[7'h7f:7'h40];
  assign T101 = T103 & T102;
  assign T102 = io_write_bits_wmask[1'h1:1'h1];
  assign T103 = T104 & io_write_valid;
  assign T104 = T70 != 2'h0;
  assign T106 = T107 ? raddr : R105;
  assign io_resp_3 = T109;
  assign T109 = T110;
  assign T110 = {T115, T111};
  assign T111 = T113 ? T115 : T112;
  assign T112 = T62[7'h7f:7'h40];
  assign T113 = T114;
  assign T114 = R86[2'h3:2'h3];
  assign T115 = T89[7'h7f:7'h40];
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T23) begin
      R21 <= raddr;
    end
    if(io_read_valid) begin
      R28 <= io_read_bits_addr;
    end
    if(T49) begin
      R47 <= raddr;
    end
    if(T81) begin
      R79 <= raddr;
    end
    if(io_read_valid) begin
      R86 <= io_read_bits_addr;
    end
    if(T107) begin
      R105 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input [3:0] io_in_3_bits_way_en,
    input [12:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [3:0] io_in_2_bits_way_en,
    input [12:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [12:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [12:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[12:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[12:0] T4;
  wire[12:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[12:0] T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[3:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : T3;
  assign T3 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = T0;
  assign T8 = T9 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign io_out_bits_way_en = T11;
  assign T11 = T16 ? T14 : T12;
  assign T12 = T13 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T13 = T7[1'h0:1'h0];
  assign T14 = T15 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T7[1'h1:1'h1];
  assign io_out_valid = T17;
  assign T17 = T22 ? T20 : T18;
  assign T18 = T19 ? io_in_1_valid : io_in_0_valid;
  assign T19 = T7[1'h0:1'h0];
  assign T20 = T21 ? io_in_3_valid : io_in_2_valid;
  assign T21 = T7[1'h0:1'h0];
  assign T22 = T7[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_2_valid;
  assign T31 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [12:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [12:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[12:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[127:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[12:0] T5;
  wire[3:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T2;
  assign T2 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T3 = T0;
  assign io_out_bits_wmask = T4;
  assign T4 = T3 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T5;
  assign T5 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [3:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T118;
  wire[87:0] T0;
  wire[87:0] T1;
  wire[87:0] T119;
  wire[87:0] T2;
  wire[87:0] wmask;
  wire[87:0] T3;
  wire[47:0] T4;
  wire[23:0] T5;
  wire[15:0] T6;
  wire[7:0] T7;
  wire[7:0] T120;
  wire T8;
  wire[10:0] T9;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[10:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[10:0] T121;
  wire[8:0] T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[10:0] T122;
  wire[7:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T123;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T124;
  wire T32;
  wire[23:0] T33;
  wire[15:0] T34;
  wire[7:0] T35;
  wire[7:0] T125;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T126;
  wire T38;
  wire[7:0] T39;
  wire[7:0] T127;
  wire T40;
  wire[39:0] T41;
  wire[23:0] T42;
  wire[15:0] T43;
  wire[7:0] T44;
  wire[7:0] T128;
  wire T45;
  wire[7:0] T46;
  wire[7:0] T129;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T130;
  wire T49;
  wire[15:0] T50;
  wire[7:0] T51;
  wire[7:0] T131;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T132;
  wire T54;
  wire[87:0] T55;
  wire[87:0] T133;
  wire[63:0] out;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] rhs;
  wire[63:0] T62;
  wire[31:0] T63;
  wire[63:0] T64;
  wire[31:0] T65;
  wire[15:0] T66;
  wire[63:0] T67;
  wire[31:0] T68;
  wire[15:0] T69;
  wire[7:0] T70;
  wire T71;
  wire max;
  wire T72;
  wire[4:0] T134;
  wire T73;
  wire[4:0] T135;
  wire min;
  wire T74;
  wire[4:0] T136;
  wire T75;
  wire[4:0] T137;
  wire less;
  wire T76;
  wire cmp_rhs;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire word;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire cmp_lhs;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire sgned;
  wire T93;
  wire[4:0] T138;
  wire T94;
  wire[4:0] T139;
  wire lt;
  wire T95;
  wire T96;
  wire lt_lo;
  wire[31:0] T97;
  wire[31:0] T98;
  wire eq_hi;
  wire[31:0] T99;
  wire[31:0] T100;
  wire lt_hi;
  wire[31:0] T101;
  wire[31:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[63:0] T106;
  wire T107;
  wire[4:0] T140;
  wire[63:0] T108;
  wire T109;
  wire[4:0] T141;
  wire[63:0] T110;
  wire T111;
  wire[4:0] T142;
  wire[63:0] adder_out;
  wire[63:0] T112;
  wire[63:0] mask;
  wire[63:0] T143;
  wire[31:0] T113;
  wire T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire T117;
  wire[4:0] T144;


  assign io_out = T118;
  assign T118 = T0[6'h3f:1'h0];
  assign T0 = T55 | T1;
  assign T1 = T2 & T119;
  assign T119 = {24'h0, io_lhs};
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T41, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = {T29, T7};
  assign T7 = 8'h0 - T120;
  assign T120 = {7'h0, T8};
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T26 ? T122 : T10;
  assign T10 = T21 ? T121 : T11;
  assign T11 = T15 ? T12 : 11'hff;
  assign T12 = 4'hf << T13;
  assign T13 = {T14, 2'h0};
  assign T14 = io_addr[2'h2:2'h2];
  assign T15 = T17 | T16;
  assign T16 = io_typ == 3'h6;
  assign T17 = io_typ == 3'h2;
  assign T121 = {2'h0, T18};
  assign T18 = 2'h3 << T19;
  assign T19 = {T20, 1'h0};
  assign T20 = io_addr[2'h2:1'h1];
  assign T21 = T23 | T22;
  assign T22 = io_typ == 3'h5;
  assign T23 = io_typ == 3'h1;
  assign T122 = {3'h0, T24};
  assign T24 = 1'h1 << T25;
  assign T25 = io_addr[2'h2:1'h0];
  assign T26 = T28 | T27;
  assign T27 = io_typ == 3'h4;
  assign T28 = io_typ == 3'h0;
  assign T29 = 8'h0 - T123;
  assign T123 = {7'h0, T30};
  assign T30 = T9[1'h1:1'h1];
  assign T31 = 8'h0 - T124;
  assign T124 = {7'h0, T32};
  assign T32 = T9[2'h2:2'h2];
  assign T33 = {T39, T34};
  assign T34 = {T37, T35};
  assign T35 = 8'h0 - T125;
  assign T125 = {7'h0, T36};
  assign T36 = T9[2'h3:2'h3];
  assign T37 = 8'h0 - T126;
  assign T126 = {7'h0, T38};
  assign T38 = T9[3'h4:3'h4];
  assign T39 = 8'h0 - T127;
  assign T127 = {7'h0, T40};
  assign T40 = T9[3'h5:3'h5];
  assign T41 = {T50, T42};
  assign T42 = {T48, T43};
  assign T43 = {T46, T44};
  assign T44 = 8'h0 - T128;
  assign T128 = {7'h0, T45};
  assign T45 = T9[3'h6:3'h6];
  assign T46 = 8'h0 - T129;
  assign T129 = {7'h0, T47};
  assign T47 = T9[3'h7:3'h7];
  assign T48 = 8'h0 - T130;
  assign T130 = {7'h0, T49};
  assign T49 = T9[4'h8:4'h8];
  assign T50 = {T53, T51};
  assign T51 = 8'h0 - T131;
  assign T131 = {7'h0, T52};
  assign T52 = T9[4'h9:4'h9];
  assign T53 = 8'h0 - T132;
  assign T132 = {7'h0, T54};
  assign T54 = T9[4'ha:4'ha];
  assign T55 = wmask & T133;
  assign T133 = {24'h0, out};
  assign out = T117 ? adder_out : T56;
  assign T56 = T111 ? T110 : T57;
  assign T57 = T109 ? T108 : T58;
  assign T58 = T107 ? T106 : T59;
  assign T59 = T71 ? io_lhs : T60;
  assign T60 = T26 ? T67 : T61;
  assign T61 = T21 ? T64 : rhs;
  assign rhs = T15 ? T62 : io_rhs;
  assign T62 = {T63, T63};
  assign T63 = io_rhs[5'h1f:1'h0];
  assign T64 = {T65, T65};
  assign T65 = {T66, T66};
  assign T66 = io_rhs[4'hf:1'h0];
  assign T67 = {T68, T68};
  assign T68 = {T69, T69};
  assign T69 = {T70, T70};
  assign T70 = io_rhs[3'h7:1'h0];
  assign T71 = less ? min : max;
  assign max = T73 | T72;
  assign T72 = T134 == 5'hf;
  assign T134 = {1'h0, io_cmd};
  assign T73 = T135 == 5'hd;
  assign T135 = {1'h0, io_cmd};
  assign min = T75 | T74;
  assign T74 = T136 == 5'he;
  assign T136 = {1'h0, io_cmd};
  assign T75 = T137 == 5'hc;
  assign T137 = {1'h0, io_cmd};
  assign less = T105 ? lt : T76;
  assign T76 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T79 ? T78 : T77;
  assign T77 = rhs[6'h3f:6'h3f];
  assign T78 = rhs[5'h1f:5'h1f];
  assign T79 = word & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_addr[2'h2:2'h2];
  assign word = T83 | T82;
  assign T82 = io_typ == 3'h4;
  assign T83 = T85 | T84;
  assign T84 = io_typ == 3'h0;
  assign T85 = T87 | T86;
  assign T86 = io_typ == 3'h6;
  assign T87 = io_typ == 3'h2;
  assign cmp_lhs = T90 ? T89 : T88;
  assign T88 = io_lhs[6'h3f:6'h3f];
  assign T89 = io_lhs[5'h1f:5'h1f];
  assign T90 = word & T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = io_addr[2'h2:2'h2];
  assign sgned = T94 | T93;
  assign T93 = T138 == 5'hd;
  assign T138 = {1'h0, io_cmd};
  assign T94 = T139 == 5'hc;
  assign T139 = {1'h0, io_cmd};
  assign lt = word ? T103 : T95;
  assign T95 = lt_hi | T96;
  assign T96 = eq_hi & lt_lo;
  assign lt_lo = T98 < T97;
  assign T97 = rhs[5'h1f:1'h0];
  assign T98 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T100 == T99;
  assign T99 = rhs[6'h3f:6'h20];
  assign T100 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T102 < T101;
  assign T101 = rhs[6'h3f:6'h20];
  assign T102 = io_lhs[6'h3f:6'h20];
  assign T103 = T104 ? lt_hi : lt_lo;
  assign T104 = io_addr[2'h2:2'h2];
  assign T105 = cmp_lhs == cmp_rhs;
  assign T106 = io_lhs ^ rhs;
  assign T107 = T140 == 5'h9;
  assign T140 = {1'h0, io_cmd};
  assign T108 = io_lhs | rhs;
  assign T109 = T141 == 5'ha;
  assign T141 = {1'h0, io_cmd};
  assign T110 = io_lhs & rhs;
  assign T111 = T142 == 5'hb;
  assign T142 = {1'h0, io_cmd};
  assign adder_out = T115 + T112;
  assign T112 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T143;
  assign T143 = {32'h0, T113};
  assign T113 = T114 << 5'h1f;
  assign T114 = io_addr[2'h2:2'h2];
  assign T115 = T116;
  assign T116 = io_lhs & mask;
  assign T117 = T144 == 5'h8;
  assign T144 = {1'h0, io_cmd};
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [2:0] io_in_1_bits_client_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [2:0] io_in_0_bits_client_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[2:0] io_out_bits_client_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[511:0] T4;
  wire[2:0] T5;
  wire[25:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_data = T4;
  assign T4 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T6;
  assign T6 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module FlowThroughSerializer_0(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [2:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input  io_in_bits_payload_uncached,
    input [1:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg  active;
  wire T50;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T51;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T52;
  wire[1:0] T20;
  wire T21;
  wire[1:0] T22;
  reg [1:0] rbits_payload_g_type;
  wire[1:0] T53;
  wire[1:0] T23;
  wire T24;
  reg  rbits_payload_uncached;
  wire T54;
  wire T25;
  wire[2:0] T26;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T55;
  wire[2:0] T27;
  wire[2:0] T28;
  reg [2:0] rbits_payload_client_xact_id;
  wire[2:0] T56;
  wire[2:0] T29;
  wire[511:0] T30;
  wire[511:0] T31;
  reg [511:0] rbits_payload_data;
  wire[511:0] T57;
  wire[511:0] T32;
  wire[511:0] T58;
  wire[127:0] T33;
  wire[127:0] T34;
  wire[127:0] shifter_0;
  wire[127:0] T35;
  wire[127:0] shifter_1;
  wire[127:0] T36;
  wire T37;
  wire[1:0] T38;
  wire[127:0] T39;
  wire[127:0] shifter_2;
  wire[127:0] T40;
  wire[127:0] shifter_3;
  wire[127:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  reg [1:0] rbits_header_dst;
  wire[1:0] T59;
  wire[1:0] T45;
  wire[1:0] T46;
  reg [1:0] rbits_header_src;
  wire[1:0] T60;
  wire[1:0] T47;
  wire T48;
  wire T49;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    active = {1{$random}};
    cnt = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_uncached = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T16 ? 1'h1 : T1;
  assign T1 = T7 ? T2 : 1'h0;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_bits_payload_uncached ? 1'h0 : T4;
  assign T4 = T6 | T5;
  assign T5 = io_in_bits_payload_g_type == 2'h2;
  assign T6 = io_in_bits_payload_g_type == 2'h1;
  assign T7 = T8 & io_in_valid;
  assign T8 = active ^ 1'h1;
  assign T50 = reset ? 1'h0 : T9;
  assign T9 = T16 ? 1'h0 : T10;
  assign T10 = T11 ? 1'h1 : active;
  assign T11 = T7 & T12;
  assign T12 = io_in_bits_payload_uncached ? 1'h0 : T13;
  assign T13 = T15 | T14;
  assign T14 = io_in_bits_payload_g_type == 2'h2;
  assign T15 = io_in_bits_payload_g_type == 2'h1;
  assign T16 = T21 & wrap;
  assign wrap = cnt == 2'h3;
  assign T51 = reset ? 2'h0 : T17;
  assign T17 = T16 ? 2'h0 : T18;
  assign T18 = T21 ? T20 : T19;
  assign T19 = T11 ? T52 : cnt;
  assign T52 = {1'h0, io_out_ready};
  assign T20 = cnt + 2'h1;
  assign T21 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T22;
  assign T22 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T53 = reset ? io_in_bits_payload_g_type : T23;
  assign T23 = T11 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_uncached = T24;
  assign T24 = active ? rbits_payload_uncached : io_in_bits_payload_uncached;
  assign T54 = reset ? io_in_bits_payload_uncached : T25;
  assign T25 = T11 ? io_in_bits_payload_uncached : rbits_payload_uncached;
  assign io_out_bits_payload_master_xact_id = T26;
  assign T26 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T55 = reset ? io_in_bits_payload_master_xact_id : T27;
  assign T27 = T11 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T28;
  assign T28 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T56 = reset ? io_in_bits_payload_client_xact_id : T29;
  assign T29 = T11 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T30;
  assign T30 = active ? T58 : T31;
  assign T31 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T57 = reset ? io_in_bits_payload_data : T32;
  assign T32 = T11 ? io_in_bits_payload_data : rbits_payload_data;
  assign T58 = {384'h0, T33};
  assign T33 = T43 ? T39 : T34;
  assign T34 = T37 ? shifter_1 : shifter_0;
  assign shifter_0 = T35;
  assign T35 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T36;
  assign T36 = rbits_payload_data[8'hff:8'h80];
  assign T37 = T38[1'h0:1'h0];
  assign T38 = cnt;
  assign T39 = T42 ? shifter_3 : shifter_2;
  assign shifter_2 = T40;
  assign T40 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T41;
  assign T41 = rbits_payload_data[9'h1ff:9'h180];
  assign T42 = T38[1'h0:1'h0];
  assign T43 = T38[1'h1:1'h1];
  assign io_out_bits_header_dst = T44;
  assign T44 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T59 = reset ? io_in_bits_header_dst : T45;
  assign T45 = T11 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T46;
  assign T46 = active ? rbits_header_src : io_in_bits_header_src;
  assign T60 = reset ? io_in_bits_header_src : T47;
  assign T47 = T11 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T48;
  assign T48 = active | io_in_valid;
  assign io_in_ready = T49;
  assign T49 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else if(T16) begin
      active <= 1'h0;
    end else if(T11) begin
      active <= 1'h1;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T16) begin
      cnt <= 2'h0;
    end else if(T21) begin
      cnt <= T20;
    end else if(T11) begin
      cnt <= T52;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T11) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_uncached <= io_in_bits_payload_uncached;
    end else if(T11) begin
      rbits_payload_uncached <= io_in_bits_payload_uncached;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T11) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T11) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T11) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T11) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T11) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input  io_cpu_req_bits_kill,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_phys,
    input [43:0] io_cpu_req_bits_addr,
    input [8:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    input [63:0] io_cpu_req_bits_data,
    output io_cpu_resp_valid,
    output[63:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output[2:0] io_cpu_resp_bits_typ,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[8:0] io_cpu_resp_bits_tag,
    output[3:0] io_cpu_resp_bits_cmd,
    output[43:0] io_cpu_resp_bits_addr,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[8:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    output io_cpu_ordered,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[2:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[511:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_header_src,
    output[1:0] io_mem_release_bits_header_dst,
    output[25:0] io_mem_release_bits_payload_addr,
    output[2:0] io_mem_release_bits_payload_client_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type
);

  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  reg [63:0] s2_req_data;
  wire[63:0] T194;
  wire[63:0] T195;
  wire[63:0] T196;
  reg  s1_replay;
  wire T422;
  wire T25;
  wire T197;
  wire s1_write;
  wire T152;
  wire T153;
  reg [4:0] s1_req_cmd;
  wire[4:0] T18;
  wire[4:0] T19;
  wire[4:0] T20;
  reg [4:0] s2_req_cmd;
  wire[4:0] T17;
  wire s2_recycle;
  wire T21;
  reg  s2_recycle_next;
  wire T421;
  wire T22;
  wire T23;
  wire T24;
  reg  s1_valid;
  wire T423;
  wire T26;
  wire T27;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire[1:0] T28;
  wire T29;
  wire s2_hit;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  reg [1:0] R44;
  wire[1:0] T45;
  wire T46;
  reg [3:0] s2_tag_match_way;
  wire[3:0] T47;
  wire[3:0] s1_tag_match_way;
  wire[3:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] s1_tag_eq_way;
  wire[3:0] T53;
  wire[1:0] T54;
  wire T55;
  wire[18:0] T56;
  wire[31:0] s1_addr;
  wire[12:0] T57;
  reg [43:0] s1_req_addr;
  wire[43:0] T58;
  wire[43:0] T59;
  wire[43:0] T60;
  wire[43:0] T61;
  wire[43:0] T62;
  wire[43:0] T424;
  wire[31:0] T63;
  wire[25:0] T64;
  wire[43:0] T425;
  wire[31:0] T65;
  wire[25:0] T66;
  reg [43:0] s2_req_addr;
  wire[43:0] T67;
  wire[43:0] T426;
  wire T68;
  wire[18:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[18:0] T72;
  wire T73;
  wire[18:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] T87;
  reg [1:0] R88;
  wire[1:0] T89;
  wire T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire[1:0] T93;
  reg [1:0] R94;
  wire[1:0] T95;
  wire T96;
  wire[1:0] T97;
  wire[1:0] T98;
  reg [1:0] R99;
  wire[1:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire s2_tag_match;
  wire T119;
  wire s2_replay;
  wire T120;
  reg  R121;
  wire T427;
  reg  s2_valid;
  wire T428;
  wire s1_valid_masked;
  wire T122;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T198;
  wire[63:0] T199;
  wire[63:0] T200;
  wire T201;
  reg  s1_recycled;
  wire T202;
  wire[63:0] T459;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T219;
  wire[63:0] T220;
  wire[127:0] s2_data_muxed;
  wire[127:0] T221;
  wire[127:0] s2_data_3;
  wire[127:0] T222;
  wire[127:0] T223;
  reg [63:0] R224;
  wire[63:0] T431;
  wire[127:0] T225;
  wire[127:0] T432;
  wire[127:0] T226;
  wire T227;
  wire T228;
  reg [63:0] R229;
  wire[63:0] T230;
  wire[63:0] T231;
  wire T232;
  wire s1_writeback;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[127:0] T237;
  wire[127:0] T238;
  wire[127:0] s2_data_2;
  wire[127:0] T239;
  wire[127:0] T240;
  reg [63:0] R241;
  wire[63:0] T433;
  wire[127:0] T242;
  wire[127:0] T434;
  wire[127:0] T243;
  wire T244;
  wire T245;
  reg [63:0] R246;
  wire[63:0] T247;
  wire[63:0] T248;
  wire T249;
  wire T250;
  wire[127:0] T251;
  wire[127:0] T252;
  wire[127:0] s2_data_1;
  wire[127:0] T253;
  wire[127:0] T254;
  reg [63:0] R255;
  wire[63:0] T435;
  wire[127:0] T256;
  wire[127:0] T436;
  wire[127:0] T257;
  wire T258;
  wire T259;
  reg [63:0] R260;
  wire[63:0] T261;
  wire[63:0] T262;
  wire T263;
  wire T264;
  wire[127:0] T265;
  wire[127:0] s2_data_0;
  wire[127:0] T266;
  wire[127:0] T267;
  reg [63:0] R268;
  wire[63:0] T437;
  wire[127:0] T269;
  wire[127:0] T438;
  wire[127:0] T270;
  wire T271;
  wire T272;
  reg [63:0] R273;
  wire[63:0] T274;
  wire[63:0] T275;
  wire T276;
  wire T277;
  wire[63:0] T278;
  wire[127:0] T439;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T279;
  wire[63:0] T280;
  wire[63:0] T281;
  reg [63:0] s4_req_data;
  wire[63:0] T282;
  wire T283;
  reg  s3_valid;
  wire T440;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire s2_sc_fail;
  wire T204;
  wire s2_lrsc_addr_match;
  wire T205;
  wire[37:0] T206;
  reg [37:0] lrsc_addr;
  wire[37:0] T207;
  wire[37:0] T208;
  wire T16;
  wire s2_lr;
  wire T123;
  wire T124;
  wire s2_valid_masked;
  wire T125;
  wire T126;
  wire s2_nack;
  wire s2_nack_miss;
  wire T127;
  wire T128;
  wire T129;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T130;
  wire s1_nack;
  wire T131;
  wire T132;
  wire T133;
  wire[6:0] T134;
  wire T135;
  wire T136;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T420;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[4:0] T11;
  wire[4:0] T12;
  wire[4:0] T13;
  wire T14;
  wire T15;
  wire T137;
  wire s2_sc;
  wire T294;
  wire T295;
  reg [63:0] s3_req_data;
  wire[63:0] T441;
  wire[127:0] T296;
  wire[127:0] T442;
  wire[63:0] T297;
  wire[127:0] T298;
  wire[127:0] T443;
  wire[127:0] s2_data_corrected;
  wire[127:0] T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  reg [4:0] s3_req_cmd;
  wire[4:0] T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[40:0] T321;
  reg [43:0] s3_req_addr;
  wire[43:0] T322;
  wire[40:0] T444;
  wire[28:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[40:0] T334;
  wire[40:0] T445;
  wire[28:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  reg [4:0] s4_req_cmd;
  wire[4:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire[40:0] T352;
  reg [43:0] s4_req_addr;
  wire[43:0] T353;
  wire[40:0] T446;
  wire[28:0] T354;
  reg  s4_valid;
  wire T447;
  wire T355;
  reg  s2_store_bypass;
  wire T356;
  wire T357;
  reg [2:0] s2_req_typ;
  wire[2:0] T173;
  reg [2:0] s1_req_typ;
  wire[2:0] T170;
  wire[2:0] T171;
  wire[2:0] T172;
  wire[3:0] T460;
  wire[5:0] T461;
  wire[127:0] T462;
  wire[1:0] T463;
  wire T464;
  wire T465;
  wire[12:0] T466;
  reg [3:0] s3_way;
  wire[3:0] T467;
  wire[127:0] T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[12:0] T476;
  wire[12:0] T477;
  wire[12:0] T478;
  wire[127:0] T479;
  wire[127:0] T480;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[6:0] T481;
  wire[37:0] T482;
  wire[6:0] T483;
  wire[37:0] T484;
  reg  s1_req_phys;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  reg  s2_req_phys;
  wire T490;
  wire[30:0] T491;
  wire T492;
  wire T493;
  wire T494;
  wire s1_readwrite;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire s1_read;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T499;
  wire T500;
  wire[3:0] T501;
  wire[3:0] s2_replaced_way_en;
  reg [1:0] R502;
  wire[1:0] T503;
  wire[1:0] T504;
  reg [15:0] R505;
  wire[15:0] T506;
  wire[15:0] T507;
  wire[15:0] T508;
  wire[14:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire[1:0] T519;
  wire[1:0] T520;
  wire[20:0] T521;
  wire[20:0] T522;
  wire[20:0] T523;
  wire[20:0] T524;
  reg [1:0] R525;
  wire[1:0] T526;
  wire T527;
  wire T528;
  wire[3:0] s1_replaced_way_en;
  wire[1:0] T529;
  reg [18:0] R530;
  wire[18:0] T531;
  wire T532;
  wire[20:0] T533;
  wire[20:0] T534;
  wire[20:0] T535;
  wire[20:0] T536;
  reg [1:0] R537;
  wire[1:0] T538;
  wire T539;
  wire T540;
  reg [18:0] R541;
  wire[18:0] T542;
  wire T543;
  wire[20:0] T544;
  wire[20:0] T545;
  wire[20:0] T546;
  wire[20:0] T547;
  reg [1:0] R548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  reg [18:0] R552;
  wire[18:0] T553;
  wire T554;
  wire[20:0] T555;
  wire[20:0] T556;
  wire[20:0] T557;
  reg [1:0] R558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  reg [18:0] R562;
  wire[18:0] T563;
  wire T564;
  wire[1:0] T565;
  wire[18:0] T566;
  wire[18:0] T567;
  wire[18:0] T568;
  reg [8:0] s2_req_tag;
  wire[8:0] T191;
  reg [8:0] s1_req_tag;
  wire[8:0] T188;
  wire[8:0] T189;
  wire[8:0] T190;
  reg  s2_req_kill;
  wire T569;
  reg  s1_req_kill;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] probe_bits_p_type;
  wire[25:0] probe_bits_addr;
  wire T596;
  wire T597;
  wire probe_valid;
  wire[2:0] T0;
  wire[511:0] T1;
  wire[2:0] T2;
  wire[25:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire probe_ready;
  wire T7;
  wire T8;
  wire[511:0] T138;
  wire[1:0] T139;
  wire T140;
  wire[511:0] T141;
  wire[2:0] T142;
  wire[25:0] T143;
  wire[1:0] T144;
  wire[1:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T158;
  wire T165;
  wire misaligned;
  wire T166;
  wire T167;
  wire[2:0] T168;
  wire T169;
  wire T174;
  wire T175;
  wire T176;
  wire[1:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T192;
  wire T193;
  wire s1_sc;
  wire[3:0] T429;
  wire[63:0] T203;
  wire[63:0] T430;
  wire[63:0] T209;
  wire[7:0] T210;
  wire[7:0] T211;
  wire[7:0] T212;
  wire[63:0] T213;
  wire[15:0] T214;
  wire[15:0] T215;
  wire[63:0] T216;
  wire[31:0] T217;
  wire[31:0] T218;
  wire[31:0] T358;
  wire T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T448;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire[15:0] T375;
  wire T376;
  wire[47:0] T377;
  wire[47:0] T378;
  wire[47:0] T379;
  wire[47:0] T449;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire[7:0] T385;
  wire T386;
  wire[55:0] T387;
  wire[55:0] T388;
  wire[55:0] T389;
  wire[55:0] T450;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  reg  block_miss;
  wire T451;
  wire T418;
  wire T419;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[6:0] wb_io_meta_read_bits_idx;
  wire[18:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire[3:0] wb_io_data_req_bits_way_en;
  wire[12:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[25:0] wb_io_release_bits_addr;
  wire[2:0] wb_io_release_bits_client_xact_id;
  wire[511:0] wb_io_release_bits_data;
  wire[2:0] wb_io_release_bits_r_type;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[25:0] prober_io_rep_bits_addr;
  wire[2:0] prober_io_rep_bits_client_xact_id;
  wire[511:0] prober_io_rep_bits_data;
  wire[2:0] prober_io_rep_bits_r_type;
  wire prober_io_meta_read_valid;
  wire[6:0] prober_io_meta_read_bits_idx;
  wire[18:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[6:0] prober_io_meta_write_bits_idx;
  wire[3:0] prober_io_meta_write_bits_way_en;
  wire[18:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[18:0] prober_io_wb_req_bits_tag;
  wire[6:0] prober_io_wb_req_bits_idx;
  wire[3:0] prober_io_wb_req_bits_way_en;
  wire[2:0] prober_io_wb_req_bits_client_xact_id;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[18:0] meta_io_resp_3_tag;
  wire[1:0] meta_io_resp_3_coh_state;
  wire[18:0] meta_io_resp_2_tag;
  wire[1:0] meta_io_resp_2_coh_state;
  wire[18:0] meta_io_resp_1_tag;
  wire[1:0] meta_io_resp_1_coh_state;
  wire[18:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[6:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[6:0] metaWriteArb_io_out_bits_idx;
  wire[3:0] metaWriteArb_io_out_bits_way_en;
  wire[18:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_3;
  wire[127:0] data_io_resp_2;
  wire[127:0] data_io_resp_1;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire[3:0] readArb_io_out_bits_way_en;
  wire[12:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire[3:0] writeArb_io_out_bits_way_en;
  wire[12:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[25:0] releaseArb_io_out_bits_addr;
  wire[2:0] releaseArb_io_out_bits_client_xact_id;
  wire[511:0] releaseArb_io_out_bits_data;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire FlowThroughSerializer_0_io_in_ready;
  wire FlowThroughSerializer_0_io_out_valid;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_header_src;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_header_dst;
  wire[511:0] FlowThroughSerializer_0_io_out_bits_payload_data;
  wire[2:0] FlowThroughSerializer_0_io_out_bits_payload_client_xact_id;
  wire[2:0] FlowThroughSerializer_0_io_out_bits_payload_master_xact_id;
  wire FlowThroughSerializer_0_io_out_bits_payload_uncached;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_payload_g_type;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[18:0] wbArb_io_out_bits_tag;
  wire[6:0] wbArb_io_out_bits_idx;
  wire[3:0] wbArb_io_out_bits_way_en;
  wire[2:0] wbArb_io_out_bits_client_xact_id;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[18:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[29:0] dtlb_io_ptw_req_bits;
  wire mshrs_io_req_ready;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr;
  wire[2:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[511:0] mshrs_io_mem_req_bits_data;
  wire mshrs_io_mem_req_bits_uncached;
  wire[1:0] mshrs_io_mem_req_bits_a_type;
  wire[511:0] mshrs_io_mem_req_bits_subblock;
  wire[3:0] mshrs_io_mem_resp_way_en;
  wire[12:0] mshrs_io_mem_resp_addr;
  wire mshrs_io_meta_read_valid;
  wire[6:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[6:0] mshrs_io_meta_write_bits_idx;
  wire[3:0] mshrs_io_meta_write_bits_way_en;
  wire[18:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire mshrs_io_replay_bits_kill;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_phys;
  wire[43:0] mshrs_io_replay_bits_addr;
  wire[8:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire[63:0] mshrs_io_replay_bits_data;
  wire mshrs_io_mem_finish_valid;
  wire[1:0] mshrs_io_mem_finish_bits_header_src;
  wire[1:0] mshrs_io_mem_finish_bits_header_dst;
  wire[2:0] mshrs_io_mem_finish_bits_payload_master_xact_id;
  wire mshrs_io_wb_req_valid;
  wire[18:0] mshrs_io_wb_req_bits_tag;
  wire[6:0] mshrs_io_wb_req_bits_idx;
  wire[3:0] mshrs_io_wb_req_bits_way_en;
  wire[2:0] mshrs_io_wb_req_bits_client_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    R44 = {1{$random}};
    s2_tag_match_way = {1{$random}};
    s1_req_addr = {2{$random}};
    s2_req_addr = {2{$random}};
    R88 = {1{$random}};
    R94 = {1{$random}};
    R99 = {1{$random}};
    R121 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R224 = {2{$random}};
    R229 = {2{$random}};
    R241 = {2{$random}};
    R246 = {2{$random}};
    R255 = {2{$random}};
    R260 = {2{$random}};
    R268 = {2{$random}};
    R273 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R502 = {1{$random}};
    R505 = {1{$random}};
    R525 = {1{$random}};
    R530 = {1{$random}};
    R537 = {1{$random}};
    R541 = {1{$random}};
    R548 = {1{$random}};
    R552 = {1{$random}};
    R558 = {1{$random}};
    R562 = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    block_miss = {1{$random}};
  end
`endif

  assign T452 = writeArb_io_in_1_ready | T453;
  assign T453 = T454 ^ 1'h1;
  assign T454 = FlowThroughSerializer_0_io_out_bits_payload_uncached ? 1'h0 : T455;
  assign T455 = T457 | T456;
  assign T456 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 2'h2;
  assign T457 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 2'h1;
  assign T458 = io_mem_release_ready;
  assign T194 = T201 ? s1_req_data : T195;
  assign T195 = T197 ? T196 : s2_req_data;
  assign T196 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T422 = reset ? 1'h0 : T25;
  assign T25 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T197 = s1_clk_en & s1_write;
  assign s1_write = T155 | T152;
  assign T152 = T154 | T153;
  assign T153 = s1_req_cmd == 5'h4;
  assign T18 = s2_recycle ? s2_req_cmd : T19;
  assign T19 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T20;
  assign T20 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T17 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T21;
  assign T21 = s2_recycle_ecc | s2_recycle_next;
  assign T421 = reset ? 1'h0 : T22;
  assign T22 = T27 ? T23 : s2_recycle_next;
  assign T23 = T24 & s2_recycle_ecc;
  assign T24 = s1_valid | s1_replay;
  assign T423 = reset ? 1'h0 : T26;
  assign T26 = io_cpu_req_ready & io_cpu_req_valid;
  assign T27 = s1_valid | s1_replay;
  assign s2_recycle_ecc = T29 & s2_data_correctable;
  assign s2_data_correctable = T28[1'h0:1'h0];
  assign T28 = 2'h0;
  assign T29 = T119 & s2_hit;
  assign s2_hit = T102 & T30;
  assign T30 = T40 == T31;
  assign T31 = T32;
  assign T32 = T33 ? 2'h2 : T40;
  assign T33 = T37 | T34;
  assign T34 = T36 | T35;
  assign T35 = s2_req_cmd == 5'h4;
  assign T36 = s2_req_cmd[2'h3:2'h3];
  assign T37 = T39 | T38;
  assign T38 = s2_req_cmd == 5'h7;
  assign T39 = s2_req_cmd == 5'h1;
  assign T40 = T41[1'h1:1'h0];
  assign T41 = T85 | T42;
  assign T42 = T46 ? T43 : 2'h0;
  assign T43 = R44;
  assign T45 = s1_clk_en ? meta_io_resp_3_coh_state : R44;
  assign T46 = s2_tag_match_way[2'h3:2'h3];
  assign T47 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T48;
  assign T48 = {T78, T49};
  assign T49 = {T75, T50};
  assign T50 = T52 & T51;
  assign T51 = meta_io_resp_0_coh_state != 2'h0;
  assign T52 = s1_tag_eq_way[1'h0:1'h0];
  assign s1_tag_eq_way = T53;
  assign T53 = {T70, T54};
  assign T54 = {T68, T55};
  assign T55 = meta_io_resp_0_tag == T56;
  assign T56 = s1_addr >> 4'hd;
  assign s1_addr = {dtlb_io_resp_ppn, T57};
  assign T57 = s1_req_addr[4'hc:1'h0];
  assign T58 = s2_recycle ? s2_req_addr : T59;
  assign T59 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T60;
  assign T60 = prober_io_meta_read_valid ? T425 : T61;
  assign T61 = wb_io_meta_read_valid ? T424 : T62;
  assign T62 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T424 = {12'h0, T63};
  assign T63 = T64 << 3'h6;
  assign T64 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T425 = {12'h0, T65};
  assign T65 = T66 << 3'h6;
  assign T66 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T67 = s1_clk_en ? T426 : s2_req_addr;
  assign T426 = {12'h0, s1_addr};
  assign T68 = meta_io_resp_1_tag == T69;
  assign T69 = s1_addr >> 4'hd;
  assign T70 = {T73, T71};
  assign T71 = meta_io_resp_2_tag == T72;
  assign T72 = s1_addr >> 4'hd;
  assign T73 = meta_io_resp_3_tag == T74;
  assign T74 = s1_addr >> 4'hd;
  assign T75 = T77 & T76;
  assign T76 = meta_io_resp_1_coh_state != 2'h0;
  assign T77 = s1_tag_eq_way[1'h1:1'h1];
  assign T78 = {T82, T79};
  assign T79 = T81 & T80;
  assign T80 = meta_io_resp_2_coh_state != 2'h0;
  assign T81 = s1_tag_eq_way[2'h2:2'h2];
  assign T82 = T84 & T83;
  assign T83 = meta_io_resp_3_coh_state != 2'h0;
  assign T84 = s1_tag_eq_way[2'h3:2'h3];
  assign T85 = T91 | T86;
  assign T86 = T90 ? T87 : 2'h0;
  assign T87 = R88;
  assign T89 = s1_clk_en ? meta_io_resp_2_coh_state : R88;
  assign T90 = s2_tag_match_way[2'h2:2'h2];
  assign T91 = T97 | T92;
  assign T92 = T96 ? T93 : 2'h0;
  assign T93 = R94;
  assign T95 = s1_clk_en ? meta_io_resp_1_coh_state : R94;
  assign T96 = s2_tag_match_way[1'h1:1'h1];
  assign T97 = T101 ? T98 : 2'h0;
  assign T98 = R99;
  assign T100 = s1_clk_en ? meta_io_resp_0_coh_state : R99;
  assign T101 = s2_tag_match_way[1'h0:1'h0];
  assign T102 = s2_tag_match & T103;
  assign T103 = T108 ? T107 : T104;
  assign T104 = T106 | T105;
  assign T105 = T40 == 2'h2;
  assign T106 = T40 == 2'h1;
  assign T107 = T40 == 2'h2;
  assign T108 = T110 | T109;
  assign T109 = s2_req_cmd == 5'h6;
  assign T110 = T112 | T111;
  assign T111 = s2_req_cmd == 5'h3;
  assign T112 = T116 | T113;
  assign T113 = T115 | T114;
  assign T114 = s2_req_cmd == 5'h4;
  assign T115 = s2_req_cmd[2'h3:2'h3];
  assign T116 = T118 | T117;
  assign T117 = s2_req_cmd == 5'h7;
  assign T118 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 4'h0;
  assign T119 = s2_valid | s2_replay;
  assign s2_replay = R121 & T120;
  assign T120 = s2_req_cmd != 5'h5;
  assign T427 = reset ? 1'h0 : s1_replay;
  assign T428 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T122;
  assign T122 = io_cpu_req_bits_kill ^ 1'h1;
  assign T154 = s1_req_cmd[2'h3:2'h3];
  assign T155 = T157 | T156;
  assign T156 = s1_req_cmd == 5'h7;
  assign T157 = s1_req_cmd == 5'h1;
  assign T198 = s2_recycle ? s2_req_data : T199;
  assign T199 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T200;
  assign T200 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T201 = s1_clk_en & s1_recycled;
  assign T202 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T459 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T439 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> 7'h0;
  assign s2_data_uncorrected = T219;
  assign T219 = {T278, T220};
  assign T220 = s2_data_muxed[6'h3f:1'h0];
  assign s2_data_muxed = T237 | T221;
  assign T221 = T236 ? s2_data_3 : 128'h0;
  assign s2_data_3 = T222;
  assign T222 = T223;
  assign T223 = {R229, R224};
  assign T431 = T225[6'h3f:1'h0];
  assign T225 = T227 ? T226 : T432;
  assign T432 = {64'h0, R224};
  assign T226 = data_io_resp_3 >> 1'h0;
  assign T227 = s1_clk_en & T228;
  assign T228 = s1_tag_eq_way[2'h3:2'h3];
  assign T230 = T232 ? T231 : R229;
  assign T231 = data_io_resp_3 >> 7'h40;
  assign T232 = T227 & s1_writeback;
  assign s1_writeback = T234 & T233;
  assign T233 = s1_replay ^ 1'h1;
  assign T234 = s1_clk_en & T235;
  assign T235 = s1_valid ^ 1'h1;
  assign T236 = s2_tag_match_way[2'h3:2'h3];
  assign T237 = T251 | T238;
  assign T238 = T250 ? s2_data_2 : 128'h0;
  assign s2_data_2 = T239;
  assign T239 = T240;
  assign T240 = {R246, R241};
  assign T433 = T242[6'h3f:1'h0];
  assign T242 = T244 ? T243 : T434;
  assign T434 = {64'h0, R241};
  assign T243 = data_io_resp_2 >> 1'h0;
  assign T244 = s1_clk_en & T245;
  assign T245 = s1_tag_eq_way[2'h2:2'h2];
  assign T247 = T249 ? T248 : R246;
  assign T248 = data_io_resp_2 >> 7'h40;
  assign T249 = T244 & s1_writeback;
  assign T250 = s2_tag_match_way[2'h2:2'h2];
  assign T251 = T265 | T252;
  assign T252 = T264 ? s2_data_1 : 128'h0;
  assign s2_data_1 = T253;
  assign T253 = T254;
  assign T254 = {R260, R255};
  assign T435 = T256[6'h3f:1'h0];
  assign T256 = T258 ? T257 : T436;
  assign T436 = {64'h0, R255};
  assign T257 = data_io_resp_1 >> 1'h0;
  assign T258 = s1_clk_en & T259;
  assign T259 = s1_tag_eq_way[1'h1:1'h1];
  assign T261 = T263 ? T262 : R260;
  assign T262 = data_io_resp_1 >> 7'h40;
  assign T263 = T258 & s1_writeback;
  assign T264 = s2_tag_match_way[1'h1:1'h1];
  assign T265 = T277 ? s2_data_0 : 128'h0;
  assign s2_data_0 = T266;
  assign T266 = T267;
  assign T267 = {R273, R268};
  assign T437 = T269[6'h3f:1'h0];
  assign T269 = T271 ? T270 : T438;
  assign T438 = {64'h0, R268};
  assign T270 = data_io_resp_0 >> 1'h0;
  assign T271 = s1_clk_en & T272;
  assign T272 = s1_tag_eq_way[1'h0:1'h0];
  assign T274 = T276 ? T275 : R273;
  assign T275 = data_io_resp_0 >> 7'h40;
  assign T276 = T271 & s1_writeback;
  assign T277 = s2_tag_match_way[1'h0:1'h0];
  assign T278 = s2_data_muxed[7'h7f:7'h40];
  assign T439 = {64'h0, s2_store_bypass_data};
  assign T279 = T339 ? T280 : s2_store_bypass_data;
  assign T280 = T324 ? amoalu_io_out : T281;
  assign T281 = T310 ? s3_req_data : s4_req_data;
  assign T282 = T283 ? s3_req_data : s4_req_data;
  assign T283 = s3_valid & metaReadArb_io_out_valid;
  assign T440 = reset ? 1'h0 : T284;
  assign T284 = T292 & T285;
  assign T285 = T289 | T286;
  assign T286 = T288 | T287;
  assign T287 = s2_req_cmd == 5'h4;
  assign T288 = s2_req_cmd[2'h3:2'h3];
  assign T289 = T291 | T290;
  assign T290 = s2_req_cmd == 5'h7;
  assign T291 = s2_req_cmd == 5'h1;
  assign T292 = T294 & T293;
  assign T293 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T204;
  assign T204 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T205;
  assign T205 = lrsc_addr == T206;
  assign T206 = s2_req_addr >> 3'h6;
  assign T207 = T16 ? T208 : lrsc_addr;
  assign T208 = s2_req_addr >> 3'h6;
  assign T16 = T123 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T123 = T124 | s2_replay;
  assign T124 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T125;
  assign T125 = s2_valid & T126;
  assign T126 = s2_nack ^ 1'h1;
  assign s2_nack = T129 | s2_nack_miss;
  assign s2_nack_miss = T128 & T127;
  assign T127 = mshrs_io_req_ready ^ 1'h1;
  assign T128 = s2_hit ^ 1'h1;
  assign T129 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T130 = T136 ? s1_nack : s2_nack_hit;
  assign s1_nack = T135 | T131;
  assign T131 = T133 & T132;
  assign T132 = prober_io_req_ready ^ 1'h1;
  assign T133 = T134 == prober_io_meta_write_bits_idx;
  assign T134 = s1_req_addr[4'hc:3'h6];
  assign T135 = T492 & dtlb_io_resp_miss;
  assign T136 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T420 = reset ? 5'h0 : T9;
  assign T9 = io_cpu_ptw_sret ? 5'h0 : T10;
  assign T10 = T137 ? 5'h0 : T11;
  assign T11 = T14 ? 5'h1f : T12;
  assign T12 = lrsc_valid ? T13 : lrsc_count;
  assign T13 = lrsc_count - 5'h1;
  assign T14 = T16 & T15;
  assign T15 = lrsc_valid ^ 1'h1;
  assign T137 = T123 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T294 = T295 | s2_replay;
  assign T295 = s2_valid_masked & s2_hit;
  assign T441 = T296[6'h3f:1'h0];
  assign T296 = T300 ? T298 : T442;
  assign T442 = {64'h0, T297};
  assign T297 = T300 ? s2_req_data : s3_req_data;
  assign T298 = s2_data_correctable ? s2_data_corrected : T443;
  assign T443 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T299;
  assign T299 = {T278, T220};
  assign T300 = T309 & T301;
  assign T301 = T302 | s2_data_correctable;
  assign T302 = T306 | T303;
  assign T303 = T305 | T304;
  assign T304 = s2_req_cmd == 5'h4;
  assign T305 = s2_req_cmd[2'h3:2'h3];
  assign T306 = T308 | T307;
  assign T307 = s2_req_cmd == 5'h7;
  assign T308 = s2_req_cmd == 5'h1;
  assign T309 = s2_valid | s2_replay;
  assign T310 = T319 & T311;
  assign T311 = T316 | T312;
  assign T312 = T315 | T313;
  assign T313 = s3_req_cmd == 5'h4;
  assign T314 = T300 ? s2_req_cmd : s3_req_cmd;
  assign T315 = s3_req_cmd[2'h3:2'h3];
  assign T316 = T318 | T317;
  assign T317 = s3_req_cmd == 5'h7;
  assign T318 = s3_req_cmd == 5'h1;
  assign T319 = s3_valid & T320;
  assign T320 = T444 == T321;
  assign T321 = s3_req_addr >> 2'h3;
  assign T322 = T300 ? s2_req_addr : s3_req_addr;
  assign T444 = {12'h0, T323};
  assign T323 = s1_addr >> 2'h3;
  assign T324 = T332 & T325;
  assign T325 = T329 | T326;
  assign T326 = T328 | T327;
  assign T327 = s2_req_cmd == 5'h4;
  assign T328 = s2_req_cmd[2'h3:2'h3];
  assign T329 = T331 | T330;
  assign T330 = s2_req_cmd == 5'h7;
  assign T331 = s2_req_cmd == 5'h1;
  assign T332 = T336 & T333;
  assign T333 = T445 == T334;
  assign T334 = s2_req_addr >> 2'h3;
  assign T445 = {12'h0, T335};
  assign T335 = s1_addr >> 2'h3;
  assign T336 = T338 & T337;
  assign T337 = s2_sc_fail ^ 1'h1;
  assign T338 = s2_valid_masked | s2_replay;
  assign T339 = s1_clk_en & T340;
  assign T340 = T355 | T341;
  assign T341 = T350 & T342;
  assign T342 = T347 | T343;
  assign T343 = T346 | T344;
  assign T344 = s4_req_cmd == 5'h4;
  assign T345 = T283 ? s3_req_cmd : s4_req_cmd;
  assign T346 = s4_req_cmd[2'h3:2'h3];
  assign T347 = T349 | T348;
  assign T348 = s4_req_cmd == 5'h7;
  assign T349 = s4_req_cmd == 5'h1;
  assign T350 = s4_valid & T351;
  assign T351 = T446 == T352;
  assign T352 = s4_req_addr >> 2'h3;
  assign T353 = T283 ? s3_req_addr : s4_req_addr;
  assign T446 = {12'h0, T354};
  assign T354 = s1_addr >> 2'h3;
  assign T447 = reset ? 1'h0 : s3_valid;
  assign T355 = T324 | T310;
  assign T356 = T339 ? 1'h1 : T357;
  assign T357 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T173 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T170 = s2_recycle ? s2_req_typ : T171;
  assign T171 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T172;
  assign T172 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T460 = s2_req_cmd[2'h3:1'h0];
  assign T461 = s2_req_addr[3'h5:1'h0];
  assign T462 = {s3_req_data, s3_req_data};
  assign T463 = 1'h1 << T464;
  assign T464 = T465;
  assign T465 = s3_req_addr[2'h3:2'h3];
  assign T466 = s3_req_addr[4'hc:1'h0];
  assign T467 = T300 ? s2_tag_match_way : s3_way;
  assign T468 = FlowThroughSerializer_0_io_out_bits_payload_data[7'h7f:1'h0];
  assign T469 = FlowThroughSerializer_0_io_out_valid & T470;
  assign T470 = FlowThroughSerializer_0_io_out_bits_payload_uncached ? 1'h0 : T471;
  assign T471 = T473 | T472;
  assign T472 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 2'h2;
  assign T473 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 2'h1;
  assign T474 = T475 | T452;
  assign T475 = FlowThroughSerializer_0_io_out_valid ^ 1'h1;
  assign T476 = s2_req_addr[4'hc:1'h0];
  assign T477 = mshrs_io_replay_bits_addr[4'hc:1'h0];
  assign T478 = io_cpu_req_bits_addr[4'hc:1'h0];
  assign T479 = T480;
  assign T480 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T481 = T482[3'h6:1'h0];
  assign T482 = s2_req_addr >> 3'h6;
  assign T483 = T484[3'h6:1'h0];
  assign T484 = io_cpu_req_bits_addr >> 3'h6;
  assign T485 = s2_recycle ? s2_req_phys : T486;
  assign T486 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T487;
  assign T487 = prober_io_meta_read_valid ? 1'h1 : T488;
  assign T488 = wb_io_meta_read_valid ? 1'h1 : T489;
  assign T489 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T490 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T491 = s1_req_addr >> 4'hd;
  assign T492 = T494 & T493;
  assign T493 = s1_req_phys ^ 1'h1;
  assign T494 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T498 | T495;
  assign T495 = T497 | T496;
  assign T496 = s1_req_cmd == 5'h3;
  assign T497 = s1_req_cmd == 5'h2;
  assign T498 = s1_read | s1_write;
  assign s1_read = T162 | T159;
  assign T159 = T161 | T160;
  assign T160 = s1_req_cmd == 5'h4;
  assign T161 = s1_req_cmd[2'h3:2'h3];
  assign T162 = T164 | T163;
  assign T163 = s1_req_cmd == 5'h6;
  assign T164 = s1_req_cmd == 5'h0;
  assign T499 = T452 & FlowThroughSerializer_0_io_out_valid;
  assign T500 = io_mem_acquire_ready;
  assign T501 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R502;
  assign T503 = s1_clk_en ? T504 : R502;
  assign T504 = R505[1'h1:1'h0];
  assign T506 = reset ? 16'h1 : T507;
  assign T507 = T517 ? T508 : R505;
  assign T508 = {T510, T509};
  assign T509 = R505[4'hf:1'h1];
  assign T510 = T512 ^ T511;
  assign T511 = R505[3'h5:3'h5];
  assign T512 = T514 ^ T513;
  assign T513 = R505[2'h3:2'h3];
  assign T514 = T516 ^ T515;
  assign T515 = R505[2'h2:2'h2];
  assign T516 = R505[1'h0:1'h0];
  assign T517 = T518;
  assign T518 = mshrs_io_req_ready & T573;
  assign T519 = s2_tag_match ? T565 : T520;
  assign T520 = T521[1'h1:1'h0];
  assign T521 = T533 | T522;
  assign T522 = T532 ? T523 : 21'h0;
  assign T523 = T524;
  assign T524 = {R530, R525};
  assign T526 = T527 ? meta_io_resp_3_coh_state : R525;
  assign T527 = s1_clk_en & T528;
  assign T528 = s1_replaced_way_en[2'h3:2'h3];
  assign s1_replaced_way_en = 1'h1 << T529;
  assign T529 = R505[1'h1:1'h0];
  assign T531 = T527 ? meta_io_resp_3_tag : R530;
  assign T532 = s2_replaced_way_en[2'h3:2'h3];
  assign T533 = T544 | T534;
  assign T534 = T543 ? T535 : 21'h0;
  assign T535 = T536;
  assign T536 = {R541, R537};
  assign T538 = T539 ? meta_io_resp_2_coh_state : R537;
  assign T539 = s1_clk_en & T540;
  assign T540 = s1_replaced_way_en[2'h2:2'h2];
  assign T542 = T539 ? meta_io_resp_2_tag : R541;
  assign T543 = s2_replaced_way_en[2'h2:2'h2];
  assign T544 = T555 | T545;
  assign T545 = T554 ? T546 : 21'h0;
  assign T546 = T547;
  assign T547 = {R552, R548};
  assign T549 = T550 ? meta_io_resp_1_coh_state : R548;
  assign T550 = s1_clk_en & T551;
  assign T551 = s1_replaced_way_en[1'h1:1'h1];
  assign T553 = T550 ? meta_io_resp_1_tag : R552;
  assign T554 = s2_replaced_way_en[1'h1:1'h1];
  assign T555 = T564 ? T556 : 21'h0;
  assign T556 = T557;
  assign T557 = {R562, R558};
  assign T559 = T560 ? meta_io_resp_0_coh_state : R558;
  assign T560 = s1_clk_en & T561;
  assign T561 = s1_replaced_way_en[1'h0:1'h0];
  assign T563 = T560 ? meta_io_resp_0_tag : R562;
  assign T564 = s2_replaced_way_en[1'h0:1'h0];
  assign T565 = T40;
  assign T566 = s2_tag_match ? T568 : T567;
  assign T567 = T521[5'h14:2'h2];
  assign T568 = T567;
  assign T191 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T188 = s2_recycle ? s2_req_tag : T189;
  assign T189 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T190;
  assign T190 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T569 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T570 = s2_recycle ? s2_req_kill : T571;
  assign T571 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T572;
  assign T572 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T573 = s2_nack_hit ? 1'h0 : T574;
  assign T574 = T594 & T575;
  assign T575 = T583 | T576;
  assign T576 = T580 | T577;
  assign T577 = T579 | T578;
  assign T578 = s2_req_cmd == 5'h4;
  assign T579 = s2_req_cmd[2'h3:2'h3];
  assign T580 = T582 | T581;
  assign T581 = s2_req_cmd == 5'h7;
  assign T582 = s2_req_cmd == 5'h1;
  assign T583 = T591 | T584;
  assign T584 = T588 | T585;
  assign T585 = T587 | T586;
  assign T586 = s2_req_cmd == 5'h4;
  assign T587 = s2_req_cmd[2'h3:2'h3];
  assign T588 = T590 | T589;
  assign T589 = s2_req_cmd == 5'h6;
  assign T590 = s2_req_cmd == 5'h0;
  assign T591 = T593 | T592;
  assign T592 = s2_req_cmd == 5'h3;
  assign T593 = s2_req_cmd == 5'h2;
  assign T594 = s2_valid_masked & T595;
  assign T595 = s2_hit ^ 1'h1;
  assign probe_bits_p_type = io_mem_probe_bits_payload_p_type;
  assign probe_bits_addr = io_mem_probe_bits_payload_addr;
  assign T596 = probe_valid & T597;
  assign T597 = lrsc_valid ^ 1'h1;
  assign probe_valid = io_mem_probe_valid;
  assign io_mem_release_bits_payload_r_type = T0;
  assign T0 = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_payload_data = T1;
  assign T1 = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_payload_client_xact_id = T2;
  assign T2 = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_payload_addr = T3;
  assign T3 = releaseArb_io_out_bits_addr;
  assign io_mem_release_bits_header_dst = T4;
  assign T4 = 2'h0;
  assign io_mem_release_bits_header_src = T5;
  assign T5 = 2'h0;
  assign io_mem_release_valid = T6;
  assign T6 = releaseArb_io_out_valid;
  assign io_mem_probe_ready = probe_ready;
  assign probe_ready = T7;
  assign T7 = prober_io_req_ready & T8;
  assign T8 = lrsc_valid ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = mshrs_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mshrs_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = mshrs_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_0_io_in_ready;
  assign io_mem_acquire_bits_payload_subblock = T138;
  assign T138 = mshrs_io_mem_req_bits_subblock;
  assign io_mem_acquire_bits_payload_a_type = T139;
  assign T139 = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_payload_uncached = T140;
  assign T140 = mshrs_io_mem_req_bits_uncached;
  assign io_mem_acquire_bits_payload_data = T141;
  assign T141 = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_payload_client_xact_id = T142;
  assign T142 = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = T143;
  assign T143 = mshrs_io_mem_req_bits_addr;
  assign io_mem_acquire_bits_header_dst = T144;
  assign T144 = 2'h0;
  assign io_mem_acquire_bits_header_src = T145;
  assign T145 = 2'h0;
  assign io_mem_acquire_valid = T146;
  assign T146 = mshrs_io_mem_req_valid;
  assign io_cpu_ordered = T147;
  assign T147 = T149 & T148;
  assign T148 = s2_valid ^ 1'h1;
  assign T149 = mshrs_io_fence_rdy & T150;
  assign T150 = s1_valid ^ 1'h1;
  assign io_cpu_ptw_req_bits = dtlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_xcpt_pf_st = T151;
  assign T151 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T158;
  assign T158 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T165;
  assign T165 = s1_write & misaligned;
  assign misaligned = T174 | T166;
  assign T166 = T169 & T167;
  assign T167 = T168 != 3'h0;
  assign T168 = s1_req_addr[2'h2:1'h0];
  assign T169 = s1_req_typ == 3'h3;
  assign T174 = T181 | T175;
  assign T175 = T178 & T176;
  assign T176 = T177 != 2'h0;
  assign T177 = s1_req_addr[1'h1:1'h0];
  assign T178 = T180 | T179;
  assign T179 = s1_req_typ == 3'h6;
  assign T180 = s1_req_typ == 3'h2;
  assign T181 = T184 & T182;
  assign T182 = T183 != 1'h0;
  assign T183 = s1_req_addr[1'h0:1'h0];
  assign T184 = T186 | T185;
  assign T185 = s1_req_typ == 3'h5;
  assign T186 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T187;
  assign T187 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T192;
  assign T192 = s1_replay & T193;
  assign T193 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_cmd = T429;
  assign T429 = s2_req_cmd[2'h3:1'h0];
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data_subword = T203;
  assign T203 = T209 | T430;
  assign T430 = {63'h0, s2_sc_fail};
  assign T209 = {T387, T210};
  assign T210 = s2_sc ? 8'h0 : T211;
  assign T211 = T386 ? T385 : T212;
  assign T212 = T213[3'h7:1'h0];
  assign T213 = {T377, T214};
  assign T214 = T376 ? T375 : T215;
  assign T215 = T216[4'hf:1'h0];
  assign T216 = {T360, T217};
  assign T217 = T359 ? T358 : T218;
  assign T218 = s2_data_word[5'h1f:1'h0];
  assign T358 = s2_data_word[6'h3f:6'h20];
  assign T359 = s2_req_addr[2'h2:2'h2];
  assign T360 = T372 ? T362 : T361;
  assign T361 = s2_data_word[6'h3f:6'h20];
  assign T362 = 32'h0 - T448;
  assign T448 = {31'h0, T363};
  assign T363 = T365 & T364;
  assign T364 = T217[5'h1f:5'h1f];
  assign T365 = T367 | T366;
  assign T366 = s2_req_typ == 3'h3;
  assign T367 = T369 | T368;
  assign T368 = s2_req_typ == 3'h2;
  assign T369 = T371 | T370;
  assign T370 = s2_req_typ == 3'h1;
  assign T371 = s2_req_typ == 3'h0;
  assign T372 = T374 | T373;
  assign T373 = s2_req_typ == 3'h6;
  assign T374 = s2_req_typ == 3'h2;
  assign T375 = T216[5'h1f:5'h10];
  assign T376 = s2_req_addr[1'h1:1'h1];
  assign T377 = T382 ? T379 : T378;
  assign T378 = T216[6'h3f:5'h10];
  assign T379 = 48'h0 - T449;
  assign T449 = {47'h0, T380};
  assign T380 = T365 & T381;
  assign T381 = T214[4'hf:4'hf];
  assign T382 = T384 | T383;
  assign T383 = s2_req_typ == 3'h5;
  assign T384 = s2_req_typ == 3'h1;
  assign T385 = T213[4'hf:4'h8];
  assign T386 = s2_req_addr[1'h0:1'h0];
  assign T387 = T392 ? T389 : T388;
  assign T388 = T213[6'h3f:4'h8];
  assign T389 = 56'h0 - T450;
  assign T450 = {55'h0, T390};
  assign T390 = T365 & T391;
  assign T391 = T210[3'h7:3'h7];
  assign T392 = s2_sc | T393;
  assign T393 = T395 | T394;
  assign T394 = s2_req_typ == 3'h4;
  assign T395 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_has_data = T396;
  assign T396 = T397 | s2_sc;
  assign T397 = T401 | T398;
  assign T398 = T400 | T399;
  assign T399 = s2_req_cmd == 5'h4;
  assign T400 = s2_req_cmd[2'h3:2'h3];
  assign T401 = T403 | T402;
  assign T402 = s2_req_cmd == 5'h6;
  assign T403 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T404;
  assign T404 = s2_valid & s2_nack;
  assign io_cpu_resp_bits_data = T216;
  assign io_cpu_resp_valid = T405;
  assign T405 = T407 & T406;
  assign T406 = s2_data_correctable ^ 1'h1;
  assign T407 = s2_replay | T408;
  assign T408 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T409;
  assign T409 = block_miss ? 1'h0 : T410;
  assign T410 = T417 ? 1'h0 : T411;
  assign T411 = T416 ? 1'h0 : T412;
  assign T412 = T413 == 1'h0;
  assign T413 = T415 & T414;
  assign T414 = io_cpu_req_bits_phys ^ 1'h1;
  assign T415 = dtlb_io_req_ready ^ 1'h1;
  assign T416 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T417 = readArb_io_in_3_ready ^ 1'h1;
  assign T451 = reset ? 1'h0 : T418;
  assign T418 = T419 & s2_nack_miss;
  assign T419 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_tag( wbArb_io_out_bits_tag ),
       .io_req_bits_idx( wbArb_io_out_bits_idx ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr( wb_io_release_bits_addr ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T596 ),
       .io_req_bits_addr( probe_bits_addr ),
       .io_req_bits_p_type( probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr( prober_io_rep_bits_addr ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_tag( prober_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( prober_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_line_state_state( T40 )
  );
  `ifndef SYNTHESIS
    assign prober.io_req_bits_client_xact_id = {1{$random}};
  `endif
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T573 ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T566 ),
       .io_req_bits_old_meta_coh_state( T519 ),
       .io_req_bits_way_en( T501 ),
       .io_req_bits_data( s2_req_data ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( T500 ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr( mshrs_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_uncached( mshrs_io_mem_req_bits_uncached ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_subblock( mshrs_io_mem_req_bits_subblock ),
       .io_mem_resp_way_en( mshrs_io_mem_resp_way_en ),
       .io_mem_resp_addr( mshrs_io_mem_resp_addr ),
       //.io_mem_resp_wmask(  )
       //.io_mem_resp_data(  )
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_mem_grant_valid( T499 ),
       .io_mem_grant_bits_header_src( FlowThroughSerializer_0_io_out_bits_header_src ),
       .io_mem_grant_bits_header_dst( FlowThroughSerializer_0_io_out_bits_header_dst ),
       .io_mem_grant_bits_payload_data( FlowThroughSerializer_0_io_out_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( FlowThroughSerializer_0_io_out_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( FlowThroughSerializer_0_io_out_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( FlowThroughSerializer_0_io_out_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( FlowThroughSerializer_0_io_out_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( mshrs_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( mshrs_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( mshrs_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( mshrs_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T492 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T491 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_resp_miss( dtlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits( dtlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_3_tag( meta_io_resp_3_tag ),
       .io_resp_3_coh_state( meta_io_resp_3_coh_state ),
       .io_resp_2_tag( meta_io_resp_2_tag ),
       .io_resp_2_coh_state( meta_io_resp_2_coh_state ),
       .io_resp_1_tag( meta_io_resp_1_tag ),
       .io_resp_1_coh_state( meta_io_resp_1_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T483 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T481 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T479 ),
       .io_resp_3( data_io_resp_3 ),
       .io_resp_2( data_io_resp_2 ),
       .io_resp_1( data_io_resp_1 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 4'hf ),
       .io_in_3_bits_addr( T478 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 4'hf ),
       .io_in_1_bits_addr( T477 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 4'hf ),
       .io_in_0_bits_addr( T476 ),
       .io_out_ready( T474 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T469 ),
       .io_in_1_bits_way_en( mshrs_io_mem_resp_way_en ),
       .io_in_1_bits_addr( mshrs_io_mem_resp_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( T468 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T466 ),
       .io_in_0_bits_wmask( T463 ),
       .io_in_0_bits_data( T462 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T461 ),
       .io_cmd( T460 ),
       .io_typ( s2_req_typ ),
       .io_lhs( T459 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  Arbiter_4 releaseArb(
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr( prober_io_rep_bits_addr ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr( wb_io_release_bits_addr ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_out_ready( T458 ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr( releaseArb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  FlowThroughSerializer_0 FlowThroughSerializer_0(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_0_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( T452 ),
       .io_out_valid( FlowThroughSerializer_0_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( FlowThroughSerializer_0_io_out_bits_header_dst ),
       .io_out_bits_payload_data( FlowThroughSerializer_0_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( FlowThroughSerializer_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_uncached( FlowThroughSerializer_0_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_0_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_5 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_tag( prober_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( prober_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_tag( wbArb_io_out_bits_tag ),
       .io_out_bits_idx( wbArb_io_out_bits_idx ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(T201) begin
      s2_req_data <= s1_req_data;
    end else if(T197) begin
      s2_req_data <= T196;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T25;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T27) begin
      s2_recycle_next <= T23;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T26;
    end
    if(s1_clk_en) begin
      R44 <= meta_io_resp_3_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T425;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T424;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T426;
    end
    if(s1_clk_en) begin
      R88 <= meta_io_resp_2_coh_state;
    end
    if(s1_clk_en) begin
      R94 <= meta_io_resp_1_coh_state;
    end
    if(s1_clk_en) begin
      R99 <= meta_io_resp_0_coh_state;
    end
    if(reset) begin
      R121 <= 1'h0;
    end else begin
      R121 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R224 <= T431;
    if(T232) begin
      R229 <= T231;
    end
    R241 <= T433;
    if(T249) begin
      R246 <= T248;
    end
    R255 <= T435;
    if(T263) begin
      R260 <= T262;
    end
    R268 <= T437;
    if(T276) begin
      R273 <= T275;
    end
    if(T339) begin
      s2_store_bypass_data <= T280;
    end
    if(T283) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T284;
    end
    if(T16) begin
      lrsc_addr <= T208;
    end
    if(T136) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_ptw_sret) begin
      lrsc_count <= 5'h0;
    end else if(T137) begin
      lrsc_count <= 5'h0;
    end else if(T14) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T13;
    end
    s3_req_data <= T441;
    if(T300) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T300) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T283) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T283) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T339) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T300) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R502 <= T504;
    end
    if(reset) begin
      R505 <= 16'h1;
    end else if(T517) begin
      R505 <= T508;
    end
    if(T527) begin
      R525 <= meta_io_resp_3_coh_state;
    end
    if(T527) begin
      R530 <= meta_io_resp_3_tag;
    end
    if(T539) begin
      R537 <= meta_io_resp_2_coh_state;
    end
    if(T539) begin
      R541 <= meta_io_resp_2_tag;
    end
    if(T550) begin
      R548 <= meta_io_resp_1_coh_state;
    end
    if(T550) begin
      R552 <= meta_io_resp_1_tag;
    end
    if(T560) begin
      R558 <= meta_io_resp_0_coh_state;
    end
    if(T560) begin
      R562 <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T418;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [29:0] io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [29:0] io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [29:0] io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [29:0] io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [29:0] io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output[29:0] io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  reg [2:0] R11;
  wire[2:0] T111;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[29:0] T20;
  wire[29:0] T21;
  wire[29:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[29:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R11 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T18 ? 3'h1 : T2;
  assign T2 = T16 ? 3'h2 : T3;
  assign T3 = T14 ? 3'h3 : T4;
  assign T4 = T9 ? 3'h4 : T5;
  assign T5 = io_in_0_valid ? 3'h0 : T6;
  assign T6 = io_in_1_valid ? 3'h1 : T7;
  assign T7 = io_in_2_valid ? 3'h2 : T8;
  assign T8 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T9 = io_in_4_valid & T10;
  assign T10 = R11 < 3'h4;
  assign T111 = reset ? 3'h0 : T12;
  assign T12 = T13 ? T0 : R11;
  assign T13 = io_out_ready & io_out_valid;
  assign T14 = io_in_3_valid & T15;
  assign T15 = R11 < 3'h3;
  assign T16 = io_in_2_valid & T17;
  assign T17 = R11 < 3'h2;
  assign T18 = io_in_1_valid & T19;
  assign T19 = R11 < 3'h1;
  assign io_out_bits = T20;
  assign T20 = T28 ? io_in_4_bits : T21;
  assign T21 = T27 ? T25 : T22;
  assign T22 = T23 ? io_in_1_bits : io_in_0_bits;
  assign T23 = T24[1'h0:1'h0];
  assign T24 = T0;
  assign T25 = T26 ? io_in_3_bits : io_in_2_bits;
  assign T26 = T24[1'h0:1'h0];
  assign T27 = T24[1'h1:1'h1];
  assign T28 = T24[2'h2:2'h2];
  assign io_out_valid = T29;
  assign T29 = T36 ? io_in_4_valid : T30;
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_1_valid : io_in_0_valid;
  assign T32 = T24[1'h0:1'h0];
  assign T33 = T34 ? io_in_3_valid : io_in_2_valid;
  assign T34 = T24[1'h0:1'h0];
  assign T35 = T24[1'h1:1'h1];
  assign T36 = T24[2'h2:2'h2];
  assign io_in_0_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = T54 | T39;
  assign T39 = T40 ^ 1'h1;
  assign T40 = T43 | T41;
  assign T41 = io_in_4_valid & T42;
  assign T42 = R11 < 3'h4;
  assign T43 = T46 | T44;
  assign T44 = io_in_3_valid & T45;
  assign T45 = R11 < 3'h3;
  assign T46 = T49 | T47;
  assign T47 = io_in_2_valid & T48;
  assign T48 = R11 < 3'h2;
  assign T49 = T52 | T50;
  assign T50 = io_in_1_valid & T51;
  assign T51 = R11 < 3'h1;
  assign T52 = io_in_0_valid & T53;
  assign T53 = R11 < 3'h0;
  assign T54 = R11 < 3'h0;
  assign io_in_1_ready = T55;
  assign T55 = T56 & io_out_ready;
  assign T56 = T63 | T57;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T59 | io_in_0_valid;
  assign T59 = T60 | T41;
  assign T60 = T61 | T44;
  assign T61 = T62 | T47;
  assign T62 = T52 | T50;
  assign T63 = T65 & T64;
  assign T64 = R11 < 3'h1;
  assign T65 = T52 ^ 1'h1;
  assign io_in_2_ready = T66;
  assign T66 = T67 & io_out_ready;
  assign T67 = T75 | T68;
  assign T68 = T69 ^ 1'h1;
  assign T69 = T70 | io_in_1_valid;
  assign T70 = T71 | io_in_0_valid;
  assign T71 = T72 | T41;
  assign T72 = T73 | T44;
  assign T73 = T74 | T47;
  assign T74 = T52 | T50;
  assign T75 = T77 & T76;
  assign T76 = R11 < 3'h2;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T52 | T50;
  assign io_in_3_ready = T79;
  assign T79 = T80 & io_out_ready;
  assign T80 = T89 | T81;
  assign T81 = T82 ^ 1'h1;
  assign T82 = T83 | io_in_2_valid;
  assign T83 = T84 | io_in_1_valid;
  assign T84 = T85 | io_in_0_valid;
  assign T85 = T86 | T41;
  assign T86 = T87 | T44;
  assign T87 = T88 | T47;
  assign T88 = T52 | T50;
  assign T89 = T91 & T90;
  assign T90 = R11 < 3'h3;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T93 | T47;
  assign T93 = T52 | T50;
  assign io_in_4_ready = T94;
  assign T94 = T95 & io_out_ready;
  assign T95 = T105 | T96;
  assign T96 = T97 ^ 1'h1;
  assign T97 = T98 | io_in_3_valid;
  assign T98 = T99 | io_in_2_valid;
  assign T99 = T100 | io_in_1_valid;
  assign T100 = T101 | io_in_0_valid;
  assign T101 = T102 | T41;
  assign T102 = T103 | T44;
  assign T103 = T104 | T47;
  assign T104 = T52 | T50;
  assign T105 = T107 & T106;
  assign T106 = R11 < 3'h4;
  assign T107 = T108 ^ 1'h1;
  assign T108 = T109 | T44;
  assign T109 = T110 | T47;
  assign T110 = T52 | T50;

  always @(posedge clk) begin
    if(reset) begin
      R11 <= 3'h0;
    end else if(T13) begin
      R11 <= T0;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_4_req_ready,
    input  io_requestor_4_req_valid,
    input [29:0] io_requestor_4_req_bits,
    output io_requestor_4_resp_valid,
    output io_requestor_4_resp_bits_error,
    output[18:0] io_requestor_4_resp_bits_ppn,
    output[5:0] io_requestor_4_resp_bits_perm,
    output[7:0] io_requestor_4_status_ip,
    output[7:0] io_requestor_4_status_im,
    output[6:0] io_requestor_4_status_zero,
    output io_requestor_4_status_er,
    output io_requestor_4_status_vm,
    output io_requestor_4_status_s64,
    output io_requestor_4_status_u64,
    output io_requestor_4_status_ef,
    output io_requestor_4_status_pei,
    output io_requestor_4_status_ei,
    output io_requestor_4_status_ps,
    output io_requestor_4_status_s,
    output io_requestor_4_invalidate,
    output io_requestor_4_sret,
    output io_requestor_3_req_ready,
    input  io_requestor_3_req_valid,
    input [29:0] io_requestor_3_req_bits,
    output io_requestor_3_resp_valid,
    output io_requestor_3_resp_bits_error,
    output[18:0] io_requestor_3_resp_bits_ppn,
    output[5:0] io_requestor_3_resp_bits_perm,
    output[7:0] io_requestor_3_status_ip,
    output[7:0] io_requestor_3_status_im,
    output[6:0] io_requestor_3_status_zero,
    output io_requestor_3_status_er,
    output io_requestor_3_status_vm,
    output io_requestor_3_status_s64,
    output io_requestor_3_status_u64,
    output io_requestor_3_status_ef,
    output io_requestor_3_status_pei,
    output io_requestor_3_status_ei,
    output io_requestor_3_status_ps,
    output io_requestor_3_status_s,
    output io_requestor_3_invalidate,
    output io_requestor_3_sret,
    output io_requestor_2_req_ready,
    input  io_requestor_2_req_valid,
    input [29:0] io_requestor_2_req_bits,
    output io_requestor_2_resp_valid,
    output io_requestor_2_resp_bits_error,
    output[18:0] io_requestor_2_resp_bits_ppn,
    output[5:0] io_requestor_2_resp_bits_perm,
    output[7:0] io_requestor_2_status_ip,
    output[7:0] io_requestor_2_status_im,
    output[6:0] io_requestor_2_status_zero,
    output io_requestor_2_status_er,
    output io_requestor_2_status_vm,
    output io_requestor_2_status_s64,
    output io_requestor_2_status_u64,
    output io_requestor_2_status_ef,
    output io_requestor_2_status_pei,
    output io_requestor_2_status_ei,
    output io_requestor_2_status_ps,
    output io_requestor_2_status_s,
    output io_requestor_2_invalidate,
    output io_requestor_2_sret,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [29:0] io_requestor_1_req_bits,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[18:0] io_requestor_1_resp_bits_ppn,
    output[5:0] io_requestor_1_resp_bits_perm,
    output[7:0] io_requestor_1_status_ip,
    output[7:0] io_requestor_1_status_im,
    output[6:0] io_requestor_1_status_zero,
    output io_requestor_1_status_er,
    output io_requestor_1_status_vm,
    output io_requestor_1_status_s64,
    output io_requestor_1_status_u64,
    output io_requestor_1_status_ef,
    output io_requestor_1_status_pei,
    output io_requestor_1_status_ei,
    output io_requestor_1_status_ps,
    output io_requestor_1_status_s,
    output io_requestor_1_invalidate,
    output io_requestor_1_sret,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [29:0] io_requestor_0_req_bits,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[18:0] io_requestor_0_resp_bits_ppn,
    output[5:0] io_requestor_0_resp_bits_perm,
    output[7:0] io_requestor_0_status_ip,
    output[7:0] io_requestor_0_status_im,
    output[6:0] io_requestor_0_status_zero,
    output io_requestor_0_status_er,
    output io_requestor_0_status_vm,
    output io_requestor_0_status_s64,
    output io_requestor_0_status_u64,
    output io_requestor_0_status_ef,
    output io_requestor_0_status_pei,
    output io_requestor_0_status_ei,
    output io_requestor_0_status_ps,
    output io_requestor_0_status_s,
    output io_requestor_0_invalidate,
    output io_requestor_0_sret,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    //output[8:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    //output[63:0] io_mem_req_bits_data
    input  io_mem_resp_valid,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [8:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    //input  io_mem_ptw_req_valid
    //input [29:0] io_mem_ptw_req_bits
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_sret,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s
);

  wire T94;
  reg [2:0] state;
  wire[2:0] T87;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T14;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T37;
  wire T38;
  wire T39;
  reg [1:0] count;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T36;
  wire T40;
  wire T34;
  wire T35;
  wire[43:0] T86;
  wire[31:0] T0;
  wire[28:0] T1;
  wire[28:0] T2;
  wire[9:0] vpn_idx;
  wire[9:0] T3;
  wire[9:0] T4;
  wire[9:0] T5;
  reg [29:0] r_req_vpn;
  wire[29:0] T6;
  wire T7;
  wire[9:0] T8;
  wire[19:0] T9;
  wire T10;
  wire[1:0] T11;
  wire[9:0] T41;
  wire[29:0] T42;
  wire T43;
  wire[18:0] T44;
  reg [63:0] r_pte;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] T88;
  wire[31:0] T47;
  wire[12:0] T48;
  wire[18:0] T49;
  wire T50;
  wire[5:0] T51;
  wire[18:0] T89;
  wire[30:0] T52;
  wire[30:0] resp_ppn;
  wire[30:0] T53;
  wire[30:0] T54;
  wire[19:0] T55;
  wire[10:0] T56;
  wire[30:0] T57;
  wire[9:0] T58;
  wire[20:0] T59;
  wire T60;
  wire[1:0] T61;
  wire[30:0] r_resp_ppn;
  wire T62;
  wire resp_err;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  reg [2:0] r_req_dest;
  wire[2:0] T67;
  wire resp_val;
  wire T68;
  wire T69;
  wire[5:0] T70;
  wire[18:0] T90;
  wire[30:0] T71;
  wire T72;
  wire T73;
  wire[5:0] T74;
  wire[18:0] T91;
  wire[30:0] T75;
  wire T76;
  wire T77;
  wire[5:0] T78;
  wire[18:0] T92;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[5:0] T82;
  wire[18:0] T93;
  wire[30:0] T83;
  wire T84;
  wire T85;
  wire arb_io_in_4_ready;
  wire arb_io_in_3_ready;
  wire arb_io_in_2_ready;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[29:0] arb_io_out_bits;
  wire[2:0] arb_io_chosen;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    r_req_vpn = {1{$random}};
    r_pte = {2{$random}};
    r_req_dest = {1{$random}};
  end
`endif

  assign T94 = state == 3'h0;
  assign T87 = reset ? 3'h0 : T15;
  assign T15 = T35 ? 3'h0 : T16;
  assign T16 = T34 ? 3'h0 : T17;
  assign T17 = T37 ? 3'h1 : T18;
  assign T18 = T29 ? 3'h3 : T19;
  assign T19 = T28 ? 3'h4 : T20;
  assign T20 = T26 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h1 : state;
  assign T23 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T24 = T25 & io_mem_req_ready;
  assign T25 = 3'h1 == state;
  assign T26 = T27 & io_mem_resp_bits_nack;
  assign T27 = 3'h2 == state;
  assign T28 = T27 & io_mem_resp_valid;
  assign T29 = T32 & T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_mem_resp_bits_data[1'h1:1'h1];
  assign T32 = T28 & T33;
  assign T33 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T37 = T32 & T38;
  assign T38 = T40 & T39;
  assign T39 = count < 2'h2;
  assign T12 = T37 ? T36 : T13;
  assign T13 = T14 ? 2'h0 : count;
  assign T36 = count + 2'h1;
  assign T40 = T30 ^ 1'h1;
  assign T34 = 3'h3 == state;
  assign T35 = 3'h4 == state;
  assign io_mem_req_bits_cmd = 5'h0;
  assign io_mem_req_bits_addr = T86;
  assign T86 = {12'h0, T0};
  assign T0 = T1 << 2'h3;
  assign T1 = T2;
  assign T2 = {T44, vpn_idx};
  assign vpn_idx = T43 ? T41 : T3;
  assign T3 = T10 ? T8 : T4;
  assign T4 = T5[4'h9:1'h0];
  assign T5 = r_req_vpn >> 5'h14;
  assign T6 = T7 ? arb_io_out_bits : r_req_vpn;
  assign T7 = T94 & arb_io_out_valid;
  assign T8 = T9[4'h9:1'h0];
  assign T9 = r_req_vpn >> 4'ha;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = count;
  assign T41 = T42[4'h9:1'h0];
  assign T42 = r_req_vpn >> 1'h0;
  assign T43 = T11[1'h1:1'h1];
  assign T44 = r_pte[5'h1f:4'hd];
  assign T45 = io_mem_resp_valid ? io_mem_resp_bits_data : T46;
  assign T46 = T7 ? T88 : r_pte;
  assign T88 = {32'h0, T47};
  assign T47 = {T49, T48};
  assign T48 = io_mem_resp_bits_data[4'hc:1'h0];
  assign T49 = io_dpath_ptbr[5'h1f:4'hd];
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T50;
  assign T50 = state == 3'h1;
  assign io_requestor_0_sret = io_dpath_sret;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_s = io_dpath_status_s;
  assign io_requestor_0_status_ps = io_dpath_status_ps;
  assign io_requestor_0_status_ei = io_dpath_status_ei;
  assign io_requestor_0_status_pei = io_dpath_status_pei;
  assign io_requestor_0_status_ef = io_dpath_status_ef;
  assign io_requestor_0_status_u64 = io_dpath_status_u64;
  assign io_requestor_0_status_s64 = io_dpath_status_s64;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_er = io_dpath_status_er;
  assign io_requestor_0_status_zero = io_dpath_status_zero;
  assign io_requestor_0_status_im = io_dpath_status_im;
  assign io_requestor_0_status_ip = io_dpath_status_ip;
  assign io_requestor_0_resp_bits_perm = T51;
  assign T51 = r_pte[4'h8:2'h3];
  assign io_requestor_0_resp_bits_ppn = T89;
  assign T89 = T52[5'h12:1'h0];
  assign T52 = resp_ppn;
  assign resp_ppn = T62 ? r_resp_ppn : T53;
  assign T53 = T60 ? T57 : T54;
  assign T54 = {T56, T55};
  assign T55 = r_req_vpn[5'h13:1'h0];
  assign T56 = r_resp_ppn >> 5'h14;
  assign T57 = {T59, T58};
  assign T58 = r_req_vpn[4'h9:1'h0];
  assign T59 = r_resp_ppn >> 4'ha;
  assign T60 = T61[1'h0:1'h0];
  assign T61 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hd;
  assign T62 = T61[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = T64 | T63;
  assign T63 = state == 3'h2;
  assign T64 = state == 3'h4;
  assign io_requestor_0_resp_valid = T65;
  assign T65 = resp_val & T66;
  assign T66 = r_req_dest == 3'h0;
  assign T67 = T7 ? arb_io_chosen : r_req_dest;
  assign resp_val = T69 | T68;
  assign T68 = state == 3'h4;
  assign T69 = state == 3'h3;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_sret = io_dpath_sret;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_s = io_dpath_status_s;
  assign io_requestor_1_status_ps = io_dpath_status_ps;
  assign io_requestor_1_status_ei = io_dpath_status_ei;
  assign io_requestor_1_status_pei = io_dpath_status_pei;
  assign io_requestor_1_status_ef = io_dpath_status_ef;
  assign io_requestor_1_status_u64 = io_dpath_status_u64;
  assign io_requestor_1_status_s64 = io_dpath_status_s64;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_er = io_dpath_status_er;
  assign io_requestor_1_status_zero = io_dpath_status_zero;
  assign io_requestor_1_status_im = io_dpath_status_im;
  assign io_requestor_1_status_ip = io_dpath_status_ip;
  assign io_requestor_1_resp_bits_perm = T70;
  assign T70 = r_pte[4'h8:2'h3];
  assign io_requestor_1_resp_bits_ppn = T90;
  assign T90 = T71[5'h12:1'h0];
  assign T71 = resp_ppn;
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T72;
  assign T72 = resp_val & T73;
  assign T73 = r_req_dest == 3'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  assign io_requestor_2_sret = io_dpath_sret;
  assign io_requestor_2_invalidate = io_dpath_invalidate;
  assign io_requestor_2_status_s = io_dpath_status_s;
  assign io_requestor_2_status_ps = io_dpath_status_ps;
  assign io_requestor_2_status_ei = io_dpath_status_ei;
  assign io_requestor_2_status_pei = io_dpath_status_pei;
  assign io_requestor_2_status_ef = io_dpath_status_ef;
  assign io_requestor_2_status_u64 = io_dpath_status_u64;
  assign io_requestor_2_status_s64 = io_dpath_status_s64;
  assign io_requestor_2_status_vm = io_dpath_status_vm;
  assign io_requestor_2_status_er = io_dpath_status_er;
  assign io_requestor_2_status_zero = io_dpath_status_zero;
  assign io_requestor_2_status_im = io_dpath_status_im;
  assign io_requestor_2_status_ip = io_dpath_status_ip;
  assign io_requestor_2_resp_bits_perm = T74;
  assign T74 = r_pte[4'h8:2'h3];
  assign io_requestor_2_resp_bits_ppn = T91;
  assign T91 = T75[5'h12:1'h0];
  assign T75 = resp_ppn;
  assign io_requestor_2_resp_bits_error = resp_err;
  assign io_requestor_2_resp_valid = T76;
  assign T76 = resp_val & T77;
  assign T77 = r_req_dest == 3'h2;
  assign io_requestor_2_req_ready = arb_io_in_2_ready;
  assign io_requestor_3_sret = io_dpath_sret;
  assign io_requestor_3_invalidate = io_dpath_invalidate;
  assign io_requestor_3_status_s = io_dpath_status_s;
  assign io_requestor_3_status_ps = io_dpath_status_ps;
  assign io_requestor_3_status_ei = io_dpath_status_ei;
  assign io_requestor_3_status_pei = io_dpath_status_pei;
  assign io_requestor_3_status_ef = io_dpath_status_ef;
  assign io_requestor_3_status_u64 = io_dpath_status_u64;
  assign io_requestor_3_status_s64 = io_dpath_status_s64;
  assign io_requestor_3_status_vm = io_dpath_status_vm;
  assign io_requestor_3_status_er = io_dpath_status_er;
  assign io_requestor_3_status_zero = io_dpath_status_zero;
  assign io_requestor_3_status_im = io_dpath_status_im;
  assign io_requestor_3_status_ip = io_dpath_status_ip;
  assign io_requestor_3_resp_bits_perm = T78;
  assign T78 = r_pte[4'h8:2'h3];
  assign io_requestor_3_resp_bits_ppn = T92;
  assign T92 = T79[5'h12:1'h0];
  assign T79 = resp_ppn;
  assign io_requestor_3_resp_bits_error = resp_err;
  assign io_requestor_3_resp_valid = T80;
  assign T80 = resp_val & T81;
  assign T81 = r_req_dest == 3'h3;
  assign io_requestor_3_req_ready = arb_io_in_3_ready;
  assign io_requestor_4_sret = io_dpath_sret;
  assign io_requestor_4_invalidate = io_dpath_invalidate;
  assign io_requestor_4_status_s = io_dpath_status_s;
  assign io_requestor_4_status_ps = io_dpath_status_ps;
  assign io_requestor_4_status_ei = io_dpath_status_ei;
  assign io_requestor_4_status_pei = io_dpath_status_pei;
  assign io_requestor_4_status_ef = io_dpath_status_ef;
  assign io_requestor_4_status_u64 = io_dpath_status_u64;
  assign io_requestor_4_status_s64 = io_dpath_status_s64;
  assign io_requestor_4_status_vm = io_dpath_status_vm;
  assign io_requestor_4_status_er = io_dpath_status_er;
  assign io_requestor_4_status_zero = io_dpath_status_zero;
  assign io_requestor_4_status_im = io_dpath_status_im;
  assign io_requestor_4_status_ip = io_dpath_status_ip;
  assign io_requestor_4_resp_bits_perm = T82;
  assign T82 = r_pte[4'h8:2'h3];
  assign io_requestor_4_resp_bits_ppn = T93;
  assign T93 = T83[5'h12:1'h0];
  assign T83 = resp_ppn;
  assign io_requestor_4_resp_bits_error = resp_err;
  assign io_requestor_4_resp_valid = T84;
  assign T84 = resp_val & T85;
  assign T85 = r_req_dest == 3'h4;
  assign io_requestor_4_req_ready = arb_io_in_4_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_4_ready( arb_io_in_4_ready ),
       .io_in_4_valid( io_requestor_4_req_valid ),
       .io_in_4_bits( io_requestor_4_req_bits ),
       .io_in_3_ready( arb_io_in_3_ready ),
       .io_in_3_valid( io_requestor_3_req_valid ),
       .io_in_3_bits( io_requestor_3_req_bits ),
       .io_in_2_ready( arb_io_in_2_ready ),
       .io_in_2_valid( io_requestor_2_req_valid ),
       .io_in_2_bits( io_requestor_2_req_bits ),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits( io_requestor_1_req_bits ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits( io_requestor_0_req_bits ),
       .io_out_ready( T94 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits( arb_io_out_bits ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h0;
    end else if(T37) begin
      state <= 3'h1;
    end else if(T29) begin
      state <= 3'h3;
    end else if(T28) begin
      state <= 3'h4;
    end else if(T26) begin
      state <= 3'h1;
    end else if(T24) begin
      state <= 3'h2;
    end else if(T23) begin
      state <= 3'h1;
    end
    if(T37) begin
      count <= T36;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T7) begin
      r_req_vpn <= arb_io_out_bits;
    end
    if(io_mem_resp_valid) begin
      r_pte <= io_mem_resp_bits_data;
    end else if(T7) begin
      r_pte <= T88;
    end
    if(T7) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module Control(input clk, input reset,
    output[2:0] io_dpath_sel_pc,
    output io_dpath_killd,
    output io_dpath_ren_1,
    output io_dpath_ren_0,
    output[2:0] io_dpath_sel_alu2,
    output[1:0] io_dpath_sel_alu1,
    output[2:0] io_dpath_sel_imm,
    output io_dpath_fn_dw,
    output[3:0] io_dpath_fn_alu,
    output io_dpath_div_mul_val,
    output io_dpath_div_mul_kill,
    //output io_dpath_div_val
    //output io_dpath_div_kill
    output[2:0] io_dpath_csr,
    output io_dpath_sret,
    output io_dpath_mem_load,
    output io_dpath_wb_load,
    output io_dpath_ex_fp_val,
    output io_dpath_mem_fp_val,
    output io_dpath_ex_wen,
    output io_dpath_ex_valid,
    output io_dpath_mem_jalr,
    output io_dpath_mem_branch,
    output io_dpath_mem_wen,
    output io_dpath_wb_wen,
    output[2:0] io_dpath_ex_mem_type,
    output io_dpath_ex_rs2_val,
    output io_dpath_ex_rocc_val,
    output io_dpath_mem_rocc_val,
    output io_dpath_bypass_1,
    output io_dpath_bypass_0,
    output[1:0] io_dpath_bypass_src_1,
    output[1:0] io_dpath_bypass_src_0,
    output io_dpath_ll_ready,
    output io_dpath_retire,
    output io_dpath_exception,
    output[63:0] io_dpath_cause,
    output io_dpath_badvaddr_wen,
    input [31:0] io_dpath_inst,
    //input  io_dpath_jalr_eq
    input  io_dpath_mem_br_taken,
    input  io_dpath_mem_misprediction,
    input  io_dpath_div_mul_rdy,
    input  io_dpath_ll_wen,
    input [4:0] io_dpath_ll_waddr,
    input [4:0] io_dpath_ex_waddr,
    input  io_dpath_mem_rs1_ra,
    input [4:0] io_dpath_mem_waddr,
    input [4:0] io_dpath_wb_waddr,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s,
    input  io_dpath_fp_sboard_clr,
    input [4:0] io_dpath_fp_sboard_clra,
    input  io_dpath_csr_replay,
    output io_imem_req_valid,
    //output[43:0] io_imem_req_bits_pc
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_btb_update_bits_pc
    //output[42:0] io_imem_btb_update_bits_target
    //output[42:0] io_imem_btb_update_bits_returnAddr
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_mispredict,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    //output[43:0] io_dmem_req_bits_addr
    //output[8:0] io_dmem_req_bits_tag
    output[4:0] io_dmem_req_bits_cmd,
    //output[63:0] io_dmem_req_bits_data
    input  io_dmem_resp_valid,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [8:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [8:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output io_fpu_valid,
    input  io_fpu_fcsr_rdy,
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    input [4:0] io_fpu_dec_cmd,
    input  io_fpu_dec_ldst,
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    input  io_fpu_dec_swap23,
    input  io_fpu_dec_single,
    input  io_fpu_dec_fromint,
    input  io_fpu_dec_toint,
    input  io_fpu_dec_fastpipe,
    input  io_fpu_dec_fma,
    input  io_fpu_dec_round,
    input  io_fpu_sboard_set,
    input  io_fpu_sboard_clr,
    input [4:0] io_fpu_sboard_clra,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [2:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [511:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[2:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire T0;
  reg  wb_reg_xcpt;
  wire T1;
  wire T2;
  wire take_pc_wb;
  wire T3;
  reg  wb_reg_sret;
  wire T4;
  wire T5;
  wire T6;
  reg  mem_reg_replay;
  wire T7;
  wire replay_ex;
  wire replay_ex_other;
  reg  mem_reg_replay_next;
  wire T8;
  reg  ex_reg_replay_next;
  wire T9;
  wire T10;
  wire id_csr_flush;
  wire T11;
  wire T12;
  wire T13;
  wire[11:0] T14;
  wire[11:0] id_csr_addr;
  wire T15;
  wire[11:0] T16;
  wire T17;
  wire id_csr_wen;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] id_csr;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[4:0] id_raddr1;
  wire id_csr_en;
  wire id_replay_next;
  wire[31:0] T27;
  wire ctrl_killd;
  wire T28;
  wire ctrl_draind;
  wire id_interrupt;
  wire id_interrupt_unmasked;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire ctrl_stalld;
  wire id_do_fence;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire id_rocc_val;
  wire T65;
  wire[31:0] T66;
  wire T67;
  wire[31:0] T68;
  wire id_mem_val;
  wire T69;
  wire[31:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T76;
  wire T77;
  wire T78;
  wire[31:0] T79;
  wire T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire[31:0] T87;
  reg  id_reg_fence;
  wire T838;
  wire T88;
  wire T89;
  wire id_fence_next;
  wire T90;
  wire id_amo_rl;
  wire id_amo;
  wire[31:0] T91;
  wire id_fence;
  wire[31:0] T92;
  wire T93;
  wire id_fence_i;
  wire[31:0] T94;
  wire T95;
  wire id_amo_aq;
  wire id_mem_busy;
  reg  ex_reg_mem_val;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire id_rocc_busy;
  reg  wb_reg_rocc_val;
  wire T100;
  reg  mem_reg_rocc_val;
  wire T101;
  reg  ex_reg_rocc_val;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire id_stall_fpu;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[4:0] T115;
  wire[4:0] T116;
  wire[4:0] id_waddr;
  wire T117;
  reg [31:0] R118;
  wire[31:0] T839;
  wire[31:0] T119;
  wire[31:0] T120;
  wire[31:0] T121;
  wire[31:0] T122;
  wire[31:0] T123;
  wire[31:0] T124;
  wire T125;
  wire T126;
  wire replay_wb;
  wire T127;
  wire T128;
  wire replay_wb_common;
  wire T129;
  reg  wb_reg_replay;
  wire T130;
  wire T131;
  wire replay_mem;
  wire fpu_kill_mem;
  reg  mem_reg_fp_val;
  wire T132;
  reg  ex_reg_fp_val;
  wire T133;
  wire T134;
  wire dcache_kill_mem;
  reg  mem_reg_wen;
  wire T135;
  reg  ex_reg_wen;
  wire T136;
  wire id_wen;
  wire T137;
  wire[31:0] T138;
  wire T139;
  wire T140;
  wire[31:0] T141;
  wire T142;
  wire T143;
  wire[31:0] T144;
  wire T145;
  wire T146;
  wire[31:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[31:0] T151;
  wire T152;
  wire id_jal;
  wire[31:0] T153;
  wire T154;
  wire T155;
  wire[31:0] T156;
  wire T157;
  wire T158;
  wire[31:0] T159;
  wire T160;
  wire[31:0] T161;
  wire T162;
  wire T163;
  reg  wb_reg_fp_wen;
  wire T164;
  reg  mem_reg_fp_wen;
  wire T165;
  reg  ex_reg_fp_wen;
  wire T166;
  wire T167;
  wire wb_dcache_miss;
  wire T168;
  reg  wb_reg_mem_val;
  wire T169;
  reg  mem_reg_mem_val;
  wire T170;
  wire[31:0] T171;
  wire[31:0] T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire T175;
  wire[31:0] T176;
  wire[31:0] T177;
  wire[31:0] T178;
  wire[31:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[4:0] T186;
  wire[4:0] T187;
  wire[4:0] id_raddr3;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[4:0] T194;
  wire[4:0] T195;
  wire[4:0] id_raddr2;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[4:0] T202;
  wire[4:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire id_fp_val;
  wire T207;
  wire[31:0] T208;
  wire T209;
  wire T210;
  wire[31:0] T211;
  wire T212;
  wire[31:0] T213;
  wire T214;
  wire id_sboard_hazard;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire[4:0] T219;
  wire[4:0] T220;
  wire T221;
  wire[31:0] T222;
  wire[31:0] T223;
  wire[31:0] T224;
  wire[31:0] T225;
  reg [31:0] R226;
  wire[31:0] T840;
  wire[31:0] T227;
  wire[31:0] T228;
  wire[31:0] T229;
  wire[31:0] T230;
  wire[31:0] T231;
  wire T232;
  wire wb_set_sboard;
  wire T233;
  reg  wb_reg_div_mul_val;
  wire T234;
  reg  mem_reg_div_mul_val;
  wire T235;
  reg  ex_reg_div_mul_val;
  wire T236;
  wire T237;
  wire id_div_val;
  wire[31:0] T238;
  wire id_mul_val;
  wire[31:0] T239;
  wire T240;
  wire id_wen_not0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[4:0] T247;
  wire[4:0] T248;
  wire T249;
  wire id_renx2_not0;
  wire T250;
  wire id_renx2;
  wire T251;
  wire[31:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire[31:0] T256;
  wire T257;
  wire T258;
  wire[31:0] T259;
  wire T260;
  wire[31:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire[4:0] T266;
  wire[4:0] T267;
  wire T268;
  wire id_renx1_not0;
  wire T269;
  wire id_renx1;
  wire T270;
  wire[31:0] T271;
  wire T272;
  wire T273;
  wire[31:0] T274;
  wire T275;
  wire T276;
  wire[31:0] T277;
  wire T278;
  wire T279;
  wire[31:0] T280;
  wire T281;
  wire T282;
  wire[31:0] T283;
  wire T284;
  wire T285;
  wire[31:0] T286;
  wire T287;
  wire T288;
  wire[31:0] T289;
  wire T290;
  wire[31:0] T291;
  wire T292;
  wire id_wb_hazard;
  wire T293;
  wire T294;
  reg  wb_reg_fp_val;
  wire T295;
  wire fp_data_hazard_wb;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire data_hazard_wb;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  reg  wb_reg_wen;
  wire T316;
  wire T317;
  wire id_mem_hazard;
  wire T318;
  wire fp_data_hazard_mem;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  reg  mem_mem_cmd_bh;
  wire T336;
  wire ex_slow_bypass;
  wire T337;
  wire T338;
  reg [2:0] ex_reg_mem_type;
  wire[2:0] T339;
  wire[2:0] T340;
  wire[2:0] id_mem_type;
  wire[1:0] T341;
  wire T342;
  wire[31:0] T343;
  wire T344;
  wire[31:0] T345;
  wire T346;
  wire[31:0] T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  reg [4:0] ex_reg_mem_cmd;
  wire[4:0] T355;
  wire[4:0] id_mem_cmd;
  wire[3:0] T356;
  wire[2:0] T357;
  wire[1:0] T358;
  wire T359;
  wire T360;
  wire[31:0] T361;
  wire T362;
  wire T363;
  wire[31:0] T364;
  wire T365;
  wire[31:0] T366;
  wire T367;
  wire T368;
  wire[31:0] T369;
  wire T370;
  wire[31:0] T371;
  wire T372;
  wire T373;
  wire[31:0] T374;
  wire T375;
  wire T376;
  wire[31:0] T377;
  wire T378;
  wire[31:0] T379;
  wire T380;
  wire T381;
  reg [1:0] mem_reg_csr;
  wire[1:0] T382;
  reg [1:0] ex_reg_csr;
  wire[1:0] T383;
  wire data_hazard_mem;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire id_ex_hazard;
  wire T392;
  wire T393;
  wire fp_data_hazard_ex;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  reg  ex_reg_jalr;
  wire T411;
  wire id_jalr;
  wire[31:0] T412;
  wire T413;
  wire data_hazard_ex;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire take_pc;
  wire take_pc_mem;
  wire T423;
  reg  mem_reg_jal;
  wire T424;
  reg  ex_reg_jal;
  wire T425;
  wire T426;
  reg  mem_reg_jalr;
  wire T427;
  reg  mem_reg_branch;
  wire T428;
  reg  ex_reg_branch;
  wire T429;
  wire id_branch;
  wire[31:0] T430;
  wire T431;
  wire ctrl_killx;
  wire T432;
  wire T433;
  reg  ex_reg_load_use;
  wire T434;
  wire id_load_use;
  wire T435;
  wire T436;
  wire replay_ex_structural;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  reg  mem_reg_sret;
  wire T442;
  reg  ex_reg_sret;
  wire T443;
  wire id_sret;
  wire[31:0] T444;
  wire ctrl_killm;
  wire T445;
  wire T446;
  wire killm_common;
  wire T447;
  reg  mem_reg_valid;
  wire T448;
  reg  ex_reg_valid;
  wire T449;
  wire T450;
  reg  mem_reg_xcpt;
  wire T451;
  wire ex_xcpt;
  wire T452;
  wire T453;
  reg  ex_reg_xcpt;
  wire T454;
  wire id_xcpt;
  wire T455;
  wire T456;
  wire T457;
  wire id_syscall;
  wire[31:0] T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire id_csr_fp;
  wire T463;
  wire[11:0] T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire id_csr_privileged;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire[1:0] T474;
  wire T475;
  wire T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire[1:0] T482;
  wire T483;
  wire T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire[1:0] T488;
  wire T489;
  wire T490;
  wire id_csr_invalid;
  wire T491;
  reg  T492;
  wire T494;
  wire id_int_val;
  wire T495;
  wire[31:0] T496;
  wire T497;
  wire T498;
  wire[31:0] T499;
  wire T500;
  wire T501;
  wire[31:0] T502;
  wire T503;
  wire T504;
  wire[31:0] T505;
  wire T506;
  wire T507;
  wire[31:0] T508;
  wire T509;
  wire T510;
  wire[31:0] T511;
  wire T512;
  wire T513;
  wire[31:0] T514;
  wire T515;
  wire T516;
  wire[31:0] T517;
  wire T518;
  wire T519;
  wire[31:0] T520;
  wire T521;
  wire T522;
  wire[31:0] T523;
  wire T524;
  wire T525;
  wire[31:0] T526;
  wire T527;
  wire T528;
  wire[31:0] T529;
  wire T530;
  wire T531;
  wire[31:0] T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire[31:0] T537;
  wire T538;
  wire T539;
  wire[31:0] T540;
  wire T541;
  wire T542;
  wire[31:0] T543;
  wire T544;
  wire T545;
  wire[31:0] T546;
  wire T547;
  wire T548;
  wire[31:0] T549;
  wire T550;
  wire T551;
  wire[31:0] T552;
  wire T553;
  wire T554;
  wire T555;
  wire[31:0] T556;
  wire T557;
  wire T558;
  wire[31:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[31:0] T563;
  wire T564;
  wire T565;
  wire[31:0] T566;
  wire T567;
  wire T568;
  wire[31:0] T569;
  wire T570;
  wire T571;
  wire[31:0] T572;
  wire T573;
  wire T574;
  wire[31:0] T575;
  wire T576;
  wire T577;
  wire[31:0] T578;
  wire T579;
  wire T580;
  wire[31:0] T581;
  wire T582;
  wire T583;
  wire[31:0] T584;
  wire T585;
  wire T586;
  wire[31:0] T587;
  wire T588;
  wire T589;
  wire[31:0] T590;
  wire T591;
  wire T592;
  wire[31:0] T593;
  wire T594;
  wire T595;
  wire[31:0] T596;
  wire T597;
  wire T598;
  wire[31:0] T599;
  wire T600;
  wire T601;
  wire[31:0] T602;
  wire T603;
  wire T604;
  wire[31:0] T605;
  wire T606;
  wire T607;
  reg  ex_reg_xcpt_interrupt;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire mem_xcpt;
  wire T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  reg  mem_reg_xcpt_interrupt;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire wb_rocc_val;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  reg  wb_reg_flush_inst;
  wire T629;
  reg  mem_reg_flush_inst;
  wire T630;
  reg  ex_reg_flush_inst;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T638;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T639;
  wire T640;
  wire T641;
  reg  ex_reg_btb_hit;
  wire T642;
  reg [6:0] mem_reg_btb_resp_bht_history;
  wire[6:0] T643;
  reg [6:0] ex_reg_btb_resp_bht_history;
  wire[6:0] T644;
  reg [5:0] mem_reg_btb_resp_entry;
  wire[5:0] T645;
  reg [5:0] ex_reg_btb_resp_entry;
  wire[5:0] T646;
  reg [42:0] mem_reg_btb_resp_target;
  wire[42:0] T647;
  reg [42:0] ex_reg_btb_resp_target;
  wire[42:0] T648;
  reg  mem_reg_btb_resp_taken;
  wire T649;
  reg  ex_reg_btb_resp_taken;
  wire T650;
  reg  mem_reg_btb_hit;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  reg [63:0] wb_reg_cause;
  wire[63:0] T657;
  wire[63:0] mem_cause;
  wire[63:0] T841;
  wire[3:0] T658;
  wire[3:0] T659;
  wire[3:0] T660;
  reg [63:0] mem_reg_cause;
  wire[63:0] T661;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T662;
  wire[63:0] id_cause;
  wire[63:0] T842;
  wire[3:0] T663;
  wire[3:0] T664;
  wire[3:0] T665;
  wire[3:0] T666;
  wire[3:0] T667;
  wire[3:0] T668;
  wire[3:0] T669;
  wire[63:0] id_interrupt_cause;
  wire[63:0] T670;
  wire[63:0] T671;
  wire[63:0] T672;
  wire[63:0] T673;
  wire[63:0] T674;
  wire[63:0] T675;
  wire T676;
  wire T677;
  reg  wb_reg_valid;
  wire T678;
  wire T679;
  wire[1:0] T680;
  wire[1:0] T681;
  wire[1:0] T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire[1:0] T690;
  wire[1:0] T691;
  wire[1:0] T692;
  wire T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire T720;
  wire[2:0] T843;
  reg [1:0] wb_reg_csr;
  wire[1:0] T721;
  wire T722;
  wire[3:0] T723;
  wire[3:0] id_fn_alu;
  wire[2:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire[31:0] T728;
  wire T729;
  wire T730;
  wire[31:0] T731;
  wire T732;
  wire[31:0] T733;
  wire T734;
  wire T735;
  wire[31:0] T736;
  wire T737;
  wire T738;
  wire[31:0] T739;
  wire T740;
  wire T741;
  wire[31:0] T742;
  wire T743;
  wire T744;
  wire[31:0] T745;
  wire T746;
  wire[31:0] T747;
  wire T748;
  wire T749;
  wire[31:0] T750;
  wire T751;
  wire T752;
  wire[31:0] T753;
  wire T754;
  wire T755;
  wire[31:0] T756;
  wire T757;
  wire[31:0] T758;
  wire T759;
  wire T760;
  wire[31:0] T761;
  wire T762;
  wire T763;
  wire T764;
  wire[31:0] T765;
  wire T766;
  wire[31:0] T767;
  wire T768;
  wire id_fn_dw;
  wire T769;
  wire[31:0] T770;
  wire T771;
  wire T772;
  wire[31:0] T773;
  wire T774;
  wire[31:0] T775;
  wire[2:0] T776;
  wire[2:0] id_sel_imm;
  wire[1:0] T777;
  wire T778;
  wire T779;
  wire[31:0] T780;
  wire T781;
  wire[31:0] T782;
  wire T783;
  wire T784;
  wire[31:0] T785;
  wire T786;
  wire T787;
  wire[31:0] T788;
  wire T789;
  wire T790;
  wire[31:0] T791;
  wire T792;
  wire[31:0] T793;
  wire[1:0] T794;
  wire[1:0] id_sel_alu1;
  wire T795;
  wire T796;
  wire[31:0] T797;
  wire T798;
  wire T799;
  wire[31:0] T800;
  wire T801;
  wire T802;
  wire[31:0] T803;
  wire T804;
  wire T805;
  wire[31:0] T806;
  wire T807;
  wire T808;
  wire[31:0] T809;
  wire T810;
  wire[31:0] T811;
  wire T812;
  wire T813;
  wire[31:0] T814;
  wire T815;
  wire[31:0] T816;
  wire[2:0] T844;
  wire[1:0] T817;
  wire[1:0] id_sel_alu2;
  wire T818;
  wire T819;
  wire[31:0] T820;
  wire T821;
  wire T822;
  wire T823;
  wire[31:0] T824;
  wire T825;
  wire T826;
  wire[31:0] T827;
  wire T828;
  wire T829;
  wire[31:0] T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire[2:0] T845;
  wire[1:0] T835;
  wire[1:0] T836;
  wire[1:0] T837;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_xcpt = {1{$random}};
    wb_reg_sret = {1{$random}};
    mem_reg_replay = {1{$random}};
    mem_reg_replay_next = {1{$random}};
    ex_reg_replay_next = {1{$random}};
    id_reg_fence = {1{$random}};
    ex_reg_mem_val = {1{$random}};
    wb_reg_rocc_val = {1{$random}};
    mem_reg_rocc_val = {1{$random}};
    ex_reg_rocc_val = {1{$random}};
    R118 = {1{$random}};
    wb_reg_replay = {1{$random}};
    mem_reg_fp_val = {1{$random}};
    ex_reg_fp_val = {1{$random}};
    mem_reg_wen = {1{$random}};
    ex_reg_wen = {1{$random}};
    wb_reg_fp_wen = {1{$random}};
    mem_reg_fp_wen = {1{$random}};
    ex_reg_fp_wen = {1{$random}};
    wb_reg_mem_val = {1{$random}};
    mem_reg_mem_val = {1{$random}};
    R226 = {1{$random}};
    wb_reg_div_mul_val = {1{$random}};
    mem_reg_div_mul_val = {1{$random}};
    ex_reg_div_mul_val = {1{$random}};
    wb_reg_fp_val = {1{$random}};
    wb_reg_wen = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_reg_mem_type = {1{$random}};
    ex_reg_mem_cmd = {1{$random}};
    mem_reg_csr = {1{$random}};
    ex_reg_csr = {1{$random}};
    ex_reg_jalr = {1{$random}};
    mem_reg_jal = {1{$random}};
    ex_reg_jal = {1{$random}};
    mem_reg_jalr = {1{$random}};
    mem_reg_branch = {1{$random}};
    ex_reg_branch = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_reg_sret = {1{$random}};
    ex_reg_sret = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    wb_reg_flush_inst = {1{$random}};
    mem_reg_flush_inst = {1{$random}};
    ex_reg_flush_inst = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_valid = {1{$random}};
    wb_reg_csr = {1{$random}};
  end
`endif

  assign io_rocc_exception = T0;
  assign T0 = wb_reg_xcpt & io_dpath_status_er;
  assign T1 = mem_xcpt & T2;
  assign T2 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T3;
  assign T3 = T612 | wb_reg_sret;
  assign T4 = ctrl_killm ? 1'h0 : T5;
  assign T5 = mem_reg_sret & T6;
  assign T6 = mem_reg_replay ^ 1'h1;
  assign T7 = T441 & replay_ex;
  assign replay_ex = replay_ex_structural | replay_ex_other;
  assign replay_ex_other = T433 | mem_reg_replay_next;
  assign T8 = ctrl_killx ? 1'h0 : ex_reg_replay_next;
  assign T9 = ctrl_killd ? 1'h0 : T10;
  assign T10 = id_replay_next | id_csr_flush;
  assign id_csr_flush = T17 & T11;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T15 | T13;
  assign T13 = T14 == 12'h400;
  assign T14 = id_csr_addr & 12'hc2d;
  assign id_csr_addr = io_dpath_inst[5'h1f:5'h14];
  assign T15 = T16 == 12'h400;
  assign T16 = id_csr_addr & 12'hc2e;
  assign T17 = id_csr_en & id_csr_wen;
  assign id_csr_wen = T26 | T18;
  assign T18 = T19 ^ 1'h1;
  assign T19 = T25 | T20;
  assign T20 = 2'h3 == id_csr;
  assign id_csr = {T23, T21};
  assign T21 = T22 == 32'h1070;
  assign T22 = io_dpath_inst & 32'h1078;
  assign T23 = T24 == 32'h2070;
  assign T24 = io_dpath_inst & 32'h2078;
  assign T25 = 2'h2 == id_csr;
  assign T26 = id_raddr1 != 5'h0;
  assign id_raddr1 = io_dpath_inst[5'h13:4'hf];
  assign id_csr_en = id_csr != 2'h0;
  assign id_replay_next = T27 == 32'h1008;
  assign T27 = io_dpath_inst & 32'h3058;
  assign ctrl_killd = T28;
  assign T28 = T59 | ctrl_draind;
  assign ctrl_draind = id_interrupt | ex_reg_replay_next;
  assign id_interrupt = io_dpath_status_ei & id_interrupt_unmasked;
  assign id_interrupt_unmasked = T32 | T29;
  assign T29 = T31 & T30;
  assign T30 = io_dpath_status_ip[3'h7:3'h7];
  assign T31 = io_dpath_status_im[3'h7:3'h7];
  assign T32 = T36 | T33;
  assign T33 = T35 & T34;
  assign T34 = io_dpath_status_ip[3'h6:3'h6];
  assign T35 = io_dpath_status_im[3'h6:3'h6];
  assign T36 = T40 | T37;
  assign T37 = T39 & T38;
  assign T38 = io_dpath_status_ip[3'h5:3'h5];
  assign T39 = io_dpath_status_im[3'h5:3'h5];
  assign T40 = T44 | T41;
  assign T41 = T43 & T42;
  assign T42 = io_dpath_status_ip[3'h4:3'h4];
  assign T43 = io_dpath_status_im[3'h4:3'h4];
  assign T44 = T48 | T45;
  assign T45 = T47 & T46;
  assign T46 = io_dpath_status_ip[2'h3:2'h3];
  assign T47 = io_dpath_status_im[2'h3:2'h3];
  assign T48 = T52 | T49;
  assign T49 = T51 & T50;
  assign T50 = io_dpath_status_ip[2'h2:2'h2];
  assign T51 = io_dpath_status_im[2'h2:2'h2];
  assign T52 = T56 | T53;
  assign T53 = T55 & T54;
  assign T54 = io_dpath_status_ip[1'h1:1'h1];
  assign T55 = io_dpath_status_im[1'h1:1'h1];
  assign T56 = T58 & T57;
  assign T57 = io_dpath_status_ip[1'h0:1'h0];
  assign T58 = io_dpath_status_im[1'h0:1'h0];
  assign T59 = T422 | ctrl_stalld;
  assign ctrl_stalld = T106 | id_do_fence;
  assign id_do_fence = T99 | T60;
  assign T60 = id_mem_busy & T61;
  assign T61 = T62 | id_csr_flush;
  assign T62 = T93 | T63;
  assign T63 = id_reg_fence & T64;
  assign T64 = id_mem_val | id_rocc_val;
  assign id_rocc_val = T67 | T65;
  assign T65 = T66 == 32'h58;
  assign T66 = io_dpath_inst & 32'h58;
  assign T67 = T68 == 32'h8;
  assign T68 = io_dpath_inst & 32'h5c;
  assign id_mem_val = T71 | T69;
  assign T69 = T70 == 32'h1000202f;
  assign T70 = io_dpath_inst & 32'hf9f0607f;
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h800202f;
  assign T73 = io_dpath_inst & 32'he800607f;
  assign T74 = T77 | T75;
  assign T75 = T76 == 32'h202f;
  assign T76 = io_dpath_inst & 32'h1800607f;
  assign T77 = T80 | T78;
  assign T78 = T79 == 32'h2003;
  assign T79 = io_dpath_inst & 32'h605b;
  assign T80 = T83 | T81;
  assign T81 = T82 == 32'h3;
  assign T82 = io_dpath_inst & 32'h107f;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h3;
  assign T85 = io_dpath_inst & 32'h207f;
  assign T86 = T87 == 32'h3;
  assign T87 = io_dpath_inst & 32'h405f;
  assign T838 = reset ? 1'h0 : T88;
  assign T88 = id_fence_next | T89;
  assign T89 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_fence | T90;
  assign T90 = id_amo & id_amo_rl;
  assign id_amo_rl = io_dpath_inst[5'h19:5'h19];
  assign id_amo = T91 == 32'h200c;
  assign T91 = io_dpath_inst & 32'h204c;
  assign id_fence = T92 == 32'h4;
  assign T92 = io_dpath_inst & 32'h3054;
  assign T93 = T95 | id_fence_i;
  assign id_fence_i = T94 == 32'h100f;
  assign T94 = io_dpath_inst & 32'h707f;
  assign T95 = id_amo & id_amo_aq;
  assign id_amo_aq = io_dpath_inst[5'h1a:5'h1a];
  assign id_mem_busy = T98 | ex_reg_mem_val;
  assign T96 = ctrl_killd ? 1'h0 : T97;
  assign T97 = id_mem_val;
  assign T98 = io_dmem_ordered ^ 1'h1;
  assign T99 = id_rocc_busy & id_fence;
  assign id_rocc_busy = T104 | wb_reg_rocc_val;
  assign T100 = ctrl_killm ? 1'h0 : mem_reg_rocc_val;
  assign T101 = ctrl_killx ? 1'h0 : ex_reg_rocc_val;
  assign T102 = ctrl_killd ? 1'h0 : T103;
  assign T103 = id_rocc_val;
  assign T104 = T105 | mem_reg_rocc_val;
  assign T105 = io_rocc_busy | ex_reg_rocc_val;
  assign T106 = T109 | T107;
  assign T107 = id_mem_val & T108;
  assign T108 = io_dmem_req_ready ^ 1'h1;
  assign T109 = T214 | T110;
  assign T110 = id_fp_val & id_stall_fpu;
  assign id_stall_fpu = T181 | T111;
  assign T111 = io_fpu_dec_wen & T112;
  assign T112 = T117 & T113;
  assign T113 = T114 - 1'h1;
  assign T114 = 1'h1 << T115;
  assign T115 = T116 + 5'h1;
  assign T116 = id_waddr - id_waddr;
  assign id_waddr = io_dpath_inst[4'hb:3'h7];
  assign T117 = R118 >> id_waddr;
  assign T839 = reset ? 32'h0 : T119;
  assign T119 = T180 ? T176 : T120;
  assign T120 = T175 ? T171 : T121;
  assign T121 = T125 ? T122 : R118;
  assign T122 = R118 | T123;
  assign T123 = T125 ? T124 : 32'h0;
  assign T124 = 1'h1 << io_dpath_wb_waddr;
  assign T125 = T162 & T126;
  assign T126 = replay_wb ^ 1'h1;
  assign replay_wb = replay_wb_common | T127;
  assign T127 = wb_reg_rocc_val & T128;
  assign T128 = io_rocc_cmd_ready ^ 1'h1;
  assign replay_wb_common = T129 | io_dpath_csr_replay;
  assign T129 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T130 = replay_mem & T131;
  assign T131 = take_pc_wb ^ 1'h1;
  assign replay_mem = T134 | fpu_kill_mem;
  assign fpu_kill_mem = mem_reg_fp_val & io_fpu_nack_mem;
  assign T132 = ctrl_killx ? 1'h0 : ex_reg_fp_val;
  assign T133 = ctrl_killd ? 1'h0 : id_fp_val;
  assign T134 = dcache_kill_mem | mem_reg_replay;
  assign dcache_kill_mem = mem_reg_wen & io_dmem_replay_next_valid;
  assign T135 = ctrl_killx ? 1'h0 : ex_reg_wen;
  assign T136 = ctrl_killd ? 1'h0 : id_wen;
  assign id_wen = T139 | T137;
  assign T137 = T138 == 32'h80000010;
  assign T138 = io_dpath_inst & 32'h90000038;
  assign T139 = T142 | T140;
  assign T140 = T141 == 32'h4018;
  assign T141 = io_dpath_inst & 32'h4018;
  assign T142 = T145 | T143;
  assign T143 = T144 == 32'h4000;
  assign T144 = io_dpath_inst & 32'h4040;
  assign T145 = T148 | T146;
  assign T146 = T147 == 32'h2030;
  assign T147 = io_dpath_inst & 32'h2038;
  assign T148 = T149 | id_amo;
  assign T149 = T152 | T150;
  assign T150 = T151 == 32'h1030;
  assign T151 = io_dpath_inst & 32'h1038;
  assign T152 = T154 | id_jal;
  assign id_jal = T153 == 32'h68;
  assign T153 = io_dpath_inst & 32'h78;
  assign T154 = T157 | T155;
  assign T155 = T156 == 32'h24;
  assign T156 = io_dpath_inst & 32'h2024;
  assign T157 = T160 | T158;
  assign T158 = T159 == 32'h10;
  assign T159 = io_dpath_inst & 32'h50;
  assign T160 = T161 == 32'h0;
  assign T161 = io_dpath_inst & 32'h6c;
  assign T162 = T163 | io_fpu_sboard_set;
  assign T163 = wb_dcache_miss & wb_reg_fp_wen;
  assign T164 = ctrl_killm ? 1'h0 : mem_reg_fp_wen;
  assign T165 = ctrl_killx ? 1'h0 : ex_reg_fp_wen;
  assign T166 = ctrl_killd ? 1'h0 : T167;
  assign T167 = id_fp_val & io_fpu_dec_wen;
  assign wb_dcache_miss = wb_reg_mem_val & T168;
  assign T168 = io_dmem_resp_valid ^ 1'h1;
  assign T169 = ctrl_killm ? 1'h0 : mem_reg_mem_val;
  assign T170 = ctrl_killx ? 1'h0 : ex_reg_mem_val;
  assign T171 = T122 & T172;
  assign T172 = ~ T173;
  assign T173 = io_dpath_fp_sboard_clr ? T174 : 32'h0;
  assign T174 = 1'h1 << io_dpath_fp_sboard_clra;
  assign T175 = T125 | io_dpath_fp_sboard_clr;
  assign T176 = T171 & T177;
  assign T177 = ~ T178;
  assign T178 = io_fpu_sboard_clr ? T179 : 32'h0;
  assign T179 = 1'h1 << io_fpu_sboard_clra;
  assign T180 = T175 | io_fpu_sboard_clr;
  assign T181 = T189 | T182;
  assign T182 = io_fpu_dec_ren3 & T183;
  assign T183 = T188 & T184;
  assign T184 = T185 - 1'h1;
  assign T185 = 1'h1 << T186;
  assign T186 = T187 + 5'h1;
  assign T187 = id_raddr3 - id_raddr3;
  assign id_raddr3 = io_dpath_inst[5'h1f:5'h1b];
  assign T188 = R118 >> id_raddr3;
  assign T189 = T197 | T190;
  assign T190 = io_fpu_dec_ren2 & T191;
  assign T191 = T196 & T192;
  assign T192 = T193 - 1'h1;
  assign T193 = 1'h1 << T194;
  assign T194 = T195 + 5'h1;
  assign T195 = id_raddr2 - id_raddr2;
  assign id_raddr2 = io_dpath_inst[5'h18:5'h14];
  assign T196 = R118 >> id_raddr2;
  assign T197 = T205 | T198;
  assign T198 = io_fpu_dec_ren1 & T199;
  assign T199 = T204 & T200;
  assign T200 = T201 - 1'h1;
  assign T201 = 1'h1 << T202;
  assign T202 = T203 + 5'h1;
  assign T203 = id_raddr1 - id_raddr1;
  assign T204 = R118 >> id_raddr1;
  assign T205 = id_csr_en & T206;
  assign T206 = io_fpu_fcsr_rdy ^ 1'h1;
  assign id_fp_val = T209 | T207;
  assign T207 = T208 == 32'h40;
  assign T208 = io_dpath_inst & 32'h68;
  assign T209 = T212 | T210;
  assign T210 = T211 == 32'h40;
  assign T211 = io_dpath_inst & 32'h70;
  assign T212 = T213 == 32'h4;
  assign T213 = io_dpath_inst & 32'h5c;
  assign T214 = T292 | id_sboard_hazard;
  assign id_sboard_hazard = T242 | T215;
  assign T215 = id_wen_not0 & T216;
  assign T216 = T221 & T217;
  assign T217 = T218 - 1'h1;
  assign T218 = 1'h1 << T219;
  assign T219 = T220 + 5'h1;
  assign T220 = id_waddr - id_waddr;
  assign T221 = T222 >> id_waddr;
  assign T222 = R226 & T223;
  assign T223 = ~ T224;
  assign T224 = io_dpath_ll_wen ? T225 : 32'h0;
  assign T225 = 1'h1 << io_dpath_ll_waddr;
  assign T840 = reset ? 32'h0 : T227;
  assign T227 = T240 ? T229 : T228;
  assign T228 = io_dpath_ll_wen ? T222 : R226;
  assign T229 = T222 | T230;
  assign T230 = T232 ? T231 : 32'h0;
  assign T231 = 1'h1 << io_dpath_wb_waddr;
  assign T232 = wb_set_sboard & io_dpath_wb_wen;
  assign wb_set_sboard = T233 | wb_reg_rocc_val;
  assign T233 = wb_reg_div_mul_val | wb_dcache_miss;
  assign T234 = ctrl_killm ? 1'h0 : mem_reg_div_mul_val;
  assign T235 = ex_reg_div_mul_val & io_dpath_div_mul_rdy;
  assign T236 = ctrl_killd ? 1'h0 : T237;
  assign T237 = id_mul_val | id_div_val;
  assign id_div_val = T238 == 32'h2004030;
  assign T238 = io_dpath_inst & 32'h2004074;
  assign id_mul_val = T239 == 32'h2000030;
  assign T239 = io_dpath_inst & 32'h2004074;
  assign T240 = io_dpath_ll_wen | T232;
  assign id_wen_not0 = id_wen & T241;
  assign T241 = id_waddr != 5'h0;
  assign T242 = T262 | T243;
  assign T243 = id_renx2_not0 & T244;
  assign T244 = T249 & T245;
  assign T245 = T246 - 1'h1;
  assign T246 = 1'h1 << T247;
  assign T247 = T248 + 5'h1;
  assign T248 = id_raddr2 - id_raddr2;
  assign T249 = T222 >> id_raddr2;
  assign id_renx2_not0 = id_renx2 & T250;
  assign T250 = id_raddr2 != 5'h0;
  assign id_renx2 = T253 | T251;
  assign T251 = T252 == 32'h3018;
  assign T252 = io_dpath_inst & 32'h3018;
  assign T253 = T254 | id_amo;
  assign T254 = T257 | T255;
  assign T255 = T256 == 32'h1008;
  assign T256 = io_dpath_inst & 32'h105c;
  assign T257 = T260 | T258;
  assign T258 = T259 == 32'h30;
  assign T259 = io_dpath_inst & 32'h74;
  assign T260 = T261 == 32'h20;
  assign T261 = io_dpath_inst & 32'h3c;
  assign T262 = id_renx1_not0 & T263;
  assign T263 = T268 & T264;
  assign T264 = T265 - 1'h1;
  assign T265 = 1'h1 << T266;
  assign T266 = T267 + 5'h1;
  assign T267 = id_raddr1 - id_raddr1;
  assign T268 = T222 >> id_raddr1;
  assign id_renx1_not0 = id_renx1 & T269;
  assign T269 = id_raddr1 != 5'h0;
  assign id_renx1 = T272 | T270;
  assign T270 = T271 == 32'h0;
  assign T271 = io_dpath_inst & 32'h58;
  assign T272 = T275 | T273;
  assign T273 = T274 == 32'h90000010;
  assign T274 = io_dpath_inst & 32'h9000003c;
  assign T275 = T278 | T276;
  assign T276 = T277 == 32'h2020;
  assign T277 = io_dpath_inst & 32'h6024;
  assign T278 = T281 | T279;
  assign T279 = T280 == 32'h2018;
  assign T280 = io_dpath_inst & 32'h2018;
  assign T281 = T284 | T282;
  assign T282 = T283 == 32'h2000;
  assign T283 = io_dpath_inst & 32'h2050;
  assign T284 = T287 | T285;
  assign T285 = T286 == 32'h1020;
  assign T286 = io_dpath_inst & 32'h5024;
  assign T287 = T290 | T288;
  assign T288 = T289 == 32'h20;
  assign T289 = io_dpath_inst & 32'h38;
  assign T290 = T291 == 32'h10;
  assign T291 = io_dpath_inst & 32'h54;
  assign T292 = T317 | id_wb_hazard;
  assign id_wb_hazard = T307 | T293;
  assign T293 = fp_data_hazard_wb & T294;
  assign T294 = wb_dcache_miss | wb_reg_fp_val;
  assign T295 = ctrl_killm ? 1'h0 : mem_reg_fp_val;
  assign fp_data_hazard_wb = wb_reg_fp_wen & T296;
  assign T296 = T299 | T297;
  assign T297 = io_fpu_dec_wen & T298;
  assign T298 = id_waddr == io_dpath_wb_waddr;
  assign T299 = T302 | T300;
  assign T300 = io_fpu_dec_ren3 & T301;
  assign T301 = id_raddr3 == io_dpath_wb_waddr;
  assign T302 = T305 | T303;
  assign T303 = io_fpu_dec_ren2 & T304;
  assign T304 = id_raddr2 == io_dpath_wb_waddr;
  assign T305 = io_fpu_dec_ren1 & T306;
  assign T306 = id_raddr1 == io_dpath_wb_waddr;
  assign T307 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_reg_wen & T308;
  assign T308 = T311 | T309;
  assign T309 = id_wen_not0 & T310;
  assign T310 = id_waddr == io_dpath_wb_waddr;
  assign T311 = T314 | T312;
  assign T312 = id_renx2_not0 & T313;
  assign T313 = id_raddr2 == io_dpath_wb_waddr;
  assign T314 = id_renx1_not0 & T315;
  assign T315 = id_raddr1 == io_dpath_wb_waddr;
  assign T316 = ctrl_killm ? 1'h0 : mem_reg_wen;
  assign T317 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = T330 | T318;
  assign T318 = fp_data_hazard_mem & mem_reg_fp_val;
  assign fp_data_hazard_mem = mem_reg_fp_wen & T319;
  assign T319 = T322 | T320;
  assign T320 = io_fpu_dec_wen & T321;
  assign T321 = id_waddr == io_dpath_mem_waddr;
  assign T322 = T325 | T323;
  assign T323 = io_fpu_dec_ren3 & T324;
  assign T324 = id_raddr3 == io_dpath_mem_waddr;
  assign T325 = T328 | T326;
  assign T326 = io_fpu_dec_ren2 & T327;
  assign T327 = id_raddr2 == io_dpath_mem_waddr;
  assign T328 = io_fpu_dec_ren1 & T329;
  assign T329 = id_raddr1 == io_dpath_mem_waddr;
  assign T330 = data_hazard_mem & T331;
  assign T331 = T332 | mem_reg_rocc_val;
  assign T332 = T333 | mem_reg_fp_val;
  assign T333 = T334 | mem_reg_div_mul_val;
  assign T334 = T381 | T335;
  assign T335 = mem_reg_mem_val & mem_mem_cmd_bh;
  assign T336 = T380 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T354 | T337;
  assign T337 = T349 | T338;
  assign T338 = 3'h5 == ex_reg_mem_type;
  assign T339 = T348 ? T340 : ex_reg_mem_type;
  assign T340 = id_mem_type;
  assign id_mem_type = {T346, T341};
  assign T341 = {T344, T342};
  assign T342 = T343 == 32'h1000;
  assign T343 = io_dpath_inst & 32'h1000;
  assign T344 = T345 == 32'h2000;
  assign T345 = io_dpath_inst & 32'h2000;
  assign T346 = T347 == 32'h4000;
  assign T347 = io_dpath_inst & 32'h4000;
  assign T348 = ctrl_killd ^ 1'h1;
  assign T349 = T351 | T350;
  assign T350 = 3'h1 == ex_reg_mem_type;
  assign T351 = T353 | T352;
  assign T352 = 3'h4 == ex_reg_mem_type;
  assign T353 = 3'h0 == ex_reg_mem_type;
  assign T354 = ex_reg_mem_cmd == 5'h7;
  assign T355 = T348 ? id_mem_cmd : ex_reg_mem_cmd;
  assign id_mem_cmd = {1'h0, T356};
  assign T356 = {T378, T357};
  assign T357 = {T372, T358};
  assign T358 = {T367, T359};
  assign T359 = T362 | T360;
  assign T360 = T361 == 32'h20000020;
  assign T361 = io_dpath_inst & 32'h20000020;
  assign T362 = T365 | T363;
  assign T363 = T364 == 32'h18000020;
  assign T364 = io_dpath_inst & 32'h18000020;
  assign T365 = T366 == 32'h20;
  assign T366 = io_dpath_inst & 32'h28;
  assign T367 = T370 | T368;
  assign T368 = T369 == 32'h40000008;
  assign T369 = io_dpath_inst & 32'h40000008;
  assign T370 = T371 == 32'h10000008;
  assign T371 = io_dpath_inst & 32'h10000008;
  assign T372 = T375 | T373;
  assign T373 = T374 == 32'h80000008;
  assign T374 = io_dpath_inst & 32'h80000008;
  assign T375 = T376 | T370;
  assign T376 = T377 == 32'h8000008;
  assign T377 = io_dpath_inst & 32'h8000008;
  assign T378 = T379 == 32'h8;
  assign T379 = io_dpath_inst & 32'h18000008;
  assign T380 = ctrl_killx ^ 1'h1;
  assign T381 = mem_reg_csr != 2'h0;
  assign T382 = ctrl_killx ? 2'h0 : ex_reg_csr;
  assign T383 = ctrl_killd ? 2'h0 : id_csr;
  assign data_hazard_mem = mem_reg_wen & T384;
  assign T384 = T387 | T385;
  assign T385 = id_wen_not0 & T386;
  assign T386 = id_waddr == io_dpath_mem_waddr;
  assign T387 = T390 | T388;
  assign T388 = id_renx2_not0 & T389;
  assign T389 = id_raddr2 == io_dpath_mem_waddr;
  assign T390 = id_renx1_not0 & T391;
  assign T391 = id_raddr1 == io_dpath_mem_waddr;
  assign id_ex_hazard = T405 | T392;
  assign T392 = fp_data_hazard_ex & T393;
  assign T393 = ex_reg_mem_val | ex_reg_fp_val;
  assign fp_data_hazard_ex = ex_reg_fp_wen & T394;
  assign T394 = T397 | T395;
  assign T395 = io_fpu_dec_wen & T396;
  assign T396 = id_waddr == io_dpath_ex_waddr;
  assign T397 = T400 | T398;
  assign T398 = io_fpu_dec_ren3 & T399;
  assign T399 = id_raddr3 == io_dpath_ex_waddr;
  assign T400 = T403 | T401;
  assign T401 = io_fpu_dec_ren2 & T402;
  assign T402 = id_raddr2 == io_dpath_ex_waddr;
  assign T403 = io_fpu_dec_ren1 & T404;
  assign T404 = id_raddr1 == io_dpath_ex_waddr;
  assign T405 = data_hazard_ex & T406;
  assign T406 = T407 | ex_reg_rocc_val;
  assign T407 = T408 | ex_reg_fp_val;
  assign T408 = T409 | ex_reg_div_mul_val;
  assign T409 = T410 | ex_reg_mem_val;
  assign T410 = T413 | ex_reg_jalr;
  assign T411 = ctrl_killd ? 1'h0 : id_jalr;
  assign id_jalr = T412 == 32'h24;
  assign T412 = io_dpath_inst & 32'h203c;
  assign T413 = ex_reg_csr != 2'h0;
  assign data_hazard_ex = ex_reg_wen & T414;
  assign T414 = T417 | T415;
  assign T415 = id_wen_not0 & T416;
  assign T416 = id_waddr == io_dpath_ex_waddr;
  assign T417 = T420 | T418;
  assign T418 = id_renx2_not0 & T419;
  assign T419 = id_raddr2 == io_dpath_ex_waddr;
  assign T420 = id_renx1_not0 & T421;
  assign T421 = id_raddr1 == io_dpath_ex_waddr;
  assign T422 = T431 | take_pc;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = io_dpath_mem_misprediction & T423;
  assign T423 = T426 | mem_reg_jal;
  assign T424 = ctrl_killx ? 1'h0 : ex_reg_jal;
  assign T425 = ctrl_killd ? 1'h0 : id_jal;
  assign T426 = mem_reg_branch | mem_reg_jalr;
  assign T427 = ctrl_killx ? 1'h0 : ex_reg_jalr;
  assign T428 = ctrl_killx ? 1'h0 : ex_reg_branch;
  assign T429 = ctrl_killd ? 1'h0 : id_branch;
  assign id_branch = T430 == 32'h60;
  assign T430 = io_dpath_inst & 32'h74;
  assign T431 = io_imem_resp_valid ^ 1'h1;
  assign ctrl_killx = T432;
  assign T432 = take_pc | replay_ex;
  assign T433 = wb_dcache_miss & ex_reg_load_use;
  assign T434 = ctrl_killd ? 1'h0 : id_load_use;
  assign id_load_use = T435;
  assign T435 = mem_reg_mem_val & T436;
  assign T436 = data_hazard_mem | fp_data_hazard_mem;
  assign replay_ex_structural = T439 | T437;
  assign T437 = ex_reg_div_mul_val & T438;
  assign T438 = io_dpath_div_mul_rdy ^ 1'h1;
  assign T439 = ex_reg_mem_val & T440;
  assign T440 = io_dmem_req_ready ^ 1'h1;
  assign T441 = take_pc ^ 1'h1;
  assign T442 = ctrl_killx ? 1'h0 : ex_reg_sret;
  assign T443 = ctrl_killd ? 1'h0 : id_sret;
  assign id_sret = T444 == 32'h80000050;
  assign T444 = io_dpath_inst & 32'he0003058;
  assign ctrl_killm = T445;
  assign T445 = T446 | fpu_kill_mem;
  assign T446 = killm_common | mem_xcpt;
  assign killm_common = T450 | T447;
  assign T447 = mem_reg_valid ^ 1'h1;
  assign T448 = ctrl_killx ? 1'h0 : ex_reg_valid;
  assign T449 = ctrl_killd ? 1'h0 : 1'h1;
  assign T450 = T611 | mem_reg_xcpt;
  assign T451 = ctrl_killx ? 1'h0 : ex_xcpt;
  assign ex_xcpt = T453 | T452;
  assign T452 = ex_reg_fp_val & io_fpu_illegal_rm;
  assign T453 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T454 = ctrl_killd ? 1'h0 : id_xcpt;
  assign id_xcpt = T457 | T455;
  assign T455 = id_rocc_val & T456;
  assign T456 = io_dpath_status_er ^ 1'h1;
  assign T457 = T459 | id_syscall;
  assign id_syscall = T458 == 32'h70;
  assign T458 = io_dpath_inst & 32'h80003078;
  assign T459 = T465 | T460;
  assign T460 = T462 & T461;
  assign T461 = io_dpath_status_ef ^ 1'h1;
  assign T462 = id_fp_val | id_csr_fp;
  assign id_csr_fp = id_csr_en & T463;
  assign T463 = T464 == 12'h0;
  assign T464 = id_csr_addr & 12'h480;
  assign T465 = T468 | T466;
  assign T466 = id_sret & T467;
  assign T467 = io_dpath_status_s ^ 1'h1;
  assign T468 = T489 | id_csr_privileged;
  assign id_csr_privileged = id_csr_en & T469;
  assign T469 = T475 | T470;
  assign T470 = T471 & id_csr_wen;
  assign T471 = T473 & T472;
  assign T472 = io_dpath_status_s ^ 1'h1;
  assign T473 = T474 == 2'h1;
  assign T474 = id_csr_addr[4'h9:4'h8];
  assign T475 = T478 | T476;
  assign T476 = 2'h2 <= T477;
  assign T477 = id_csr_addr[4'h9:4'h8];
  assign T478 = T483 | T479;
  assign T479 = T481 & T480;
  assign T480 = io_dpath_status_s ^ 1'h1;
  assign T481 = T482 == 2'h1;
  assign T482 = id_csr_addr[4'hb:4'ha];
  assign T483 = T486 | T484;
  assign T484 = T485 == 2'h2;
  assign T485 = id_csr_addr[4'hb:4'ha];
  assign T486 = T487 & id_csr_wen;
  assign T487 = T488 == 2'h3;
  assign T488 = id_csr_addr[4'hb:4'ha];
  assign T489 = T606 | T490;
  assign T490 = T494 | id_csr_invalid;
  assign id_csr_invalid = id_csr_en & T491;
  assign T491 = T492 ^ 1'h1;
  always @(*) case (id_csr_addr)
    0: T492 = 1'h0;
    1: T492 = 1'h1;
    2: T492 = 1'h1;
    3: T492 = 1'h1;
    4: T492 = 1'h0;
    5: T492 = 1'h0;
    6: T492 = 1'h0;
    7: T492 = 1'h0;
    8: T492 = 1'h0;
    9: T492 = 1'h0;
    10: T492 = 1'h0;
    11: T492 = 1'h0;
    12: T492 = 1'h0;
    13: T492 = 1'h0;
    14: T492 = 1'h0;
    15: T492 = 1'h0;
    16: T492 = 1'h0;
    17: T492 = 1'h0;
    18: T492 = 1'h0;
    19: T492 = 1'h0;
    20: T492 = 1'h0;
    21: T492 = 1'h0;
    22: T492 = 1'h0;
    23: T492 = 1'h0;
    24: T492 = 1'h0;
    25: T492 = 1'h0;
    26: T492 = 1'h0;
    27: T492 = 1'h0;
    28: T492 = 1'h0;
    29: T492 = 1'h0;
    30: T492 = 1'h0;
    31: T492 = 1'h0;
    32: T492 = 1'h0;
    33: T492 = 1'h0;
    34: T492 = 1'h0;
    35: T492 = 1'h0;
    36: T492 = 1'h0;
    37: T492 = 1'h0;
    38: T492 = 1'h0;
    39: T492 = 1'h0;
    40: T492 = 1'h0;
    41: T492 = 1'h0;
    42: T492 = 1'h0;
    43: T492 = 1'h0;
    44: T492 = 1'h0;
    45: T492 = 1'h0;
    46: T492 = 1'h0;
    47: T492 = 1'h0;
    48: T492 = 1'h0;
    49: T492 = 1'h0;
    50: T492 = 1'h0;
    51: T492 = 1'h0;
    52: T492 = 1'h0;
    53: T492 = 1'h0;
    54: T492 = 1'h0;
    55: T492 = 1'h0;
    56: T492 = 1'h0;
    57: T492 = 1'h0;
    58: T492 = 1'h0;
    59: T492 = 1'h0;
    60: T492 = 1'h0;
    61: T492 = 1'h0;
    62: T492 = 1'h0;
    63: T492 = 1'h0;
    64: T492 = 1'h0;
    65: T492 = 1'h0;
    66: T492 = 1'h0;
    67: T492 = 1'h0;
    68: T492 = 1'h0;
    69: T492 = 1'h0;
    70: T492 = 1'h0;
    71: T492 = 1'h0;
    72: T492 = 1'h0;
    73: T492 = 1'h0;
    74: T492 = 1'h0;
    75: T492 = 1'h0;
    76: T492 = 1'h0;
    77: T492 = 1'h0;
    78: T492 = 1'h0;
    79: T492 = 1'h0;
    80: T492 = 1'h0;
    81: T492 = 1'h0;
    82: T492 = 1'h0;
    83: T492 = 1'h0;
    84: T492 = 1'h0;
    85: T492 = 1'h0;
    86: T492 = 1'h0;
    87: T492 = 1'h0;
    88: T492 = 1'h0;
    89: T492 = 1'h0;
    90: T492 = 1'h0;
    91: T492 = 1'h0;
    92: T492 = 1'h0;
    93: T492 = 1'h0;
    94: T492 = 1'h0;
    95: T492 = 1'h0;
    96: T492 = 1'h0;
    97: T492 = 1'h0;
    98: T492 = 1'h0;
    99: T492 = 1'h0;
    100: T492 = 1'h0;
    101: T492 = 1'h0;
    102: T492 = 1'h0;
    103: T492 = 1'h0;
    104: T492 = 1'h0;
    105: T492 = 1'h0;
    106: T492 = 1'h0;
    107: T492 = 1'h0;
    108: T492 = 1'h0;
    109: T492 = 1'h0;
    110: T492 = 1'h0;
    111: T492 = 1'h0;
    112: T492 = 1'h0;
    113: T492 = 1'h0;
    114: T492 = 1'h0;
    115: T492 = 1'h0;
    116: T492 = 1'h0;
    117: T492 = 1'h0;
    118: T492 = 1'h0;
    119: T492 = 1'h0;
    120: T492 = 1'h0;
    121: T492 = 1'h0;
    122: T492 = 1'h0;
    123: T492 = 1'h0;
    124: T492 = 1'h0;
    125: T492 = 1'h0;
    126: T492 = 1'h0;
    127: T492 = 1'h0;
    128: T492 = 1'h0;
    129: T492 = 1'h0;
    130: T492 = 1'h0;
    131: T492 = 1'h0;
    132: T492 = 1'h0;
    133: T492 = 1'h0;
    134: T492 = 1'h0;
    135: T492 = 1'h0;
    136: T492 = 1'h0;
    137: T492 = 1'h0;
    138: T492 = 1'h0;
    139: T492 = 1'h0;
    140: T492 = 1'h0;
    141: T492 = 1'h0;
    142: T492 = 1'h0;
    143: T492 = 1'h0;
    144: T492 = 1'h0;
    145: T492 = 1'h0;
    146: T492 = 1'h0;
    147: T492 = 1'h0;
    148: T492 = 1'h0;
    149: T492 = 1'h0;
    150: T492 = 1'h0;
    151: T492 = 1'h0;
    152: T492 = 1'h0;
    153: T492 = 1'h0;
    154: T492 = 1'h0;
    155: T492 = 1'h0;
    156: T492 = 1'h0;
    157: T492 = 1'h0;
    158: T492 = 1'h0;
    159: T492 = 1'h0;
    160: T492 = 1'h0;
    161: T492 = 1'h0;
    162: T492 = 1'h0;
    163: T492 = 1'h0;
    164: T492 = 1'h0;
    165: T492 = 1'h0;
    166: T492 = 1'h0;
    167: T492 = 1'h0;
    168: T492 = 1'h0;
    169: T492 = 1'h0;
    170: T492 = 1'h0;
    171: T492 = 1'h0;
    172: T492 = 1'h0;
    173: T492 = 1'h0;
    174: T492 = 1'h0;
    175: T492 = 1'h0;
    176: T492 = 1'h0;
    177: T492 = 1'h0;
    178: T492 = 1'h0;
    179: T492 = 1'h0;
    180: T492 = 1'h0;
    181: T492 = 1'h0;
    182: T492 = 1'h0;
    183: T492 = 1'h0;
    184: T492 = 1'h0;
    185: T492 = 1'h0;
    186: T492 = 1'h0;
    187: T492 = 1'h0;
    188: T492 = 1'h0;
    189: T492 = 1'h0;
    190: T492 = 1'h0;
    191: T492 = 1'h0;
    192: T492 = 1'h1;
    193: T492 = 1'h0;
    194: T492 = 1'h0;
    195: T492 = 1'h0;
    196: T492 = 1'h0;
    197: T492 = 1'h0;
    198: T492 = 1'h0;
    199: T492 = 1'h0;
    200: T492 = 1'h0;
    201: T492 = 1'h0;
    202: T492 = 1'h0;
    203: T492 = 1'h0;
    204: T492 = 1'h0;
    205: T492 = 1'h0;
    206: T492 = 1'h0;
    207: T492 = 1'h0;
    208: T492 = 1'h0;
    209: T492 = 1'h0;
    210: T492 = 1'h0;
    211: T492 = 1'h0;
    212: T492 = 1'h0;
    213: T492 = 1'h0;
    214: T492 = 1'h0;
    215: T492 = 1'h0;
    216: T492 = 1'h0;
    217: T492 = 1'h0;
    218: T492 = 1'h0;
    219: T492 = 1'h0;
    220: T492 = 1'h0;
    221: T492 = 1'h0;
    222: T492 = 1'h0;
    223: T492 = 1'h0;
    224: T492 = 1'h0;
    225: T492 = 1'h0;
    226: T492 = 1'h0;
    227: T492 = 1'h0;
    228: T492 = 1'h0;
    229: T492 = 1'h0;
    230: T492 = 1'h0;
    231: T492 = 1'h0;
    232: T492 = 1'h0;
    233: T492 = 1'h0;
    234: T492 = 1'h0;
    235: T492 = 1'h0;
    236: T492 = 1'h0;
    237: T492 = 1'h0;
    238: T492 = 1'h0;
    239: T492 = 1'h0;
    240: T492 = 1'h0;
    241: T492 = 1'h0;
    242: T492 = 1'h0;
    243: T492 = 1'h0;
    244: T492 = 1'h0;
    245: T492 = 1'h0;
    246: T492 = 1'h0;
    247: T492 = 1'h0;
    248: T492 = 1'h0;
    249: T492 = 1'h0;
    250: T492 = 1'h0;
    251: T492 = 1'h0;
    252: T492 = 1'h0;
    253: T492 = 1'h0;
    254: T492 = 1'h0;
    255: T492 = 1'h0;
    256: T492 = 1'h0;
    257: T492 = 1'h0;
    258: T492 = 1'h0;
    259: T492 = 1'h0;
    260: T492 = 1'h0;
    261: T492 = 1'h0;
    262: T492 = 1'h0;
    263: T492 = 1'h0;
    264: T492 = 1'h0;
    265: T492 = 1'h0;
    266: T492 = 1'h0;
    267: T492 = 1'h0;
    268: T492 = 1'h0;
    269: T492 = 1'h0;
    270: T492 = 1'h0;
    271: T492 = 1'h0;
    272: T492 = 1'h0;
    273: T492 = 1'h0;
    274: T492 = 1'h0;
    275: T492 = 1'h0;
    276: T492 = 1'h0;
    277: T492 = 1'h0;
    278: T492 = 1'h0;
    279: T492 = 1'h0;
    280: T492 = 1'h0;
    281: T492 = 1'h0;
    282: T492 = 1'h0;
    283: T492 = 1'h0;
    284: T492 = 1'h0;
    285: T492 = 1'h0;
    286: T492 = 1'h0;
    287: T492 = 1'h0;
    288: T492 = 1'h0;
    289: T492 = 1'h0;
    290: T492 = 1'h0;
    291: T492 = 1'h0;
    292: T492 = 1'h0;
    293: T492 = 1'h0;
    294: T492 = 1'h0;
    295: T492 = 1'h0;
    296: T492 = 1'h0;
    297: T492 = 1'h0;
    298: T492 = 1'h0;
    299: T492 = 1'h0;
    300: T492 = 1'h0;
    301: T492 = 1'h0;
    302: T492 = 1'h0;
    303: T492 = 1'h0;
    304: T492 = 1'h0;
    305: T492 = 1'h0;
    306: T492 = 1'h0;
    307: T492 = 1'h0;
    308: T492 = 1'h0;
    309: T492 = 1'h0;
    310: T492 = 1'h0;
    311: T492 = 1'h0;
    312: T492 = 1'h0;
    313: T492 = 1'h0;
    314: T492 = 1'h0;
    315: T492 = 1'h0;
    316: T492 = 1'h0;
    317: T492 = 1'h0;
    318: T492 = 1'h0;
    319: T492 = 1'h0;
    320: T492 = 1'h0;
    321: T492 = 1'h0;
    322: T492 = 1'h0;
    323: T492 = 1'h0;
    324: T492 = 1'h0;
    325: T492 = 1'h0;
    326: T492 = 1'h0;
    327: T492 = 1'h0;
    328: T492 = 1'h0;
    329: T492 = 1'h0;
    330: T492 = 1'h0;
    331: T492 = 1'h0;
    332: T492 = 1'h0;
    333: T492 = 1'h0;
    334: T492 = 1'h0;
    335: T492 = 1'h0;
    336: T492 = 1'h0;
    337: T492 = 1'h0;
    338: T492 = 1'h0;
    339: T492 = 1'h0;
    340: T492 = 1'h0;
    341: T492 = 1'h0;
    342: T492 = 1'h0;
    343: T492 = 1'h0;
    344: T492 = 1'h0;
    345: T492 = 1'h0;
    346: T492 = 1'h0;
    347: T492 = 1'h0;
    348: T492 = 1'h0;
    349: T492 = 1'h0;
    350: T492 = 1'h0;
    351: T492 = 1'h0;
    352: T492 = 1'h0;
    353: T492 = 1'h0;
    354: T492 = 1'h0;
    355: T492 = 1'h0;
    356: T492 = 1'h0;
    357: T492 = 1'h0;
    358: T492 = 1'h0;
    359: T492 = 1'h0;
    360: T492 = 1'h0;
    361: T492 = 1'h0;
    362: T492 = 1'h0;
    363: T492 = 1'h0;
    364: T492 = 1'h0;
    365: T492 = 1'h0;
    366: T492 = 1'h0;
    367: T492 = 1'h0;
    368: T492 = 1'h0;
    369: T492 = 1'h0;
    370: T492 = 1'h0;
    371: T492 = 1'h0;
    372: T492 = 1'h0;
    373: T492 = 1'h0;
    374: T492 = 1'h0;
    375: T492 = 1'h0;
    376: T492 = 1'h0;
    377: T492 = 1'h0;
    378: T492 = 1'h0;
    379: T492 = 1'h0;
    380: T492 = 1'h0;
    381: T492 = 1'h0;
    382: T492 = 1'h0;
    383: T492 = 1'h0;
    384: T492 = 1'h0;
    385: T492 = 1'h0;
    386: T492 = 1'h0;
    387: T492 = 1'h0;
    388: T492 = 1'h0;
    389: T492 = 1'h0;
    390: T492 = 1'h0;
    391: T492 = 1'h0;
    392: T492 = 1'h0;
    393: T492 = 1'h0;
    394: T492 = 1'h0;
    395: T492 = 1'h0;
    396: T492 = 1'h0;
    397: T492 = 1'h0;
    398: T492 = 1'h0;
    399: T492 = 1'h0;
    400: T492 = 1'h0;
    401: T492 = 1'h0;
    402: T492 = 1'h0;
    403: T492 = 1'h0;
    404: T492 = 1'h0;
    405: T492 = 1'h0;
    406: T492 = 1'h0;
    407: T492 = 1'h0;
    408: T492 = 1'h0;
    409: T492 = 1'h0;
    410: T492 = 1'h0;
    411: T492 = 1'h0;
    412: T492 = 1'h0;
    413: T492 = 1'h0;
    414: T492 = 1'h0;
    415: T492 = 1'h0;
    416: T492 = 1'h0;
    417: T492 = 1'h0;
    418: T492 = 1'h0;
    419: T492 = 1'h0;
    420: T492 = 1'h0;
    421: T492 = 1'h0;
    422: T492 = 1'h0;
    423: T492 = 1'h0;
    424: T492 = 1'h0;
    425: T492 = 1'h0;
    426: T492 = 1'h0;
    427: T492 = 1'h0;
    428: T492 = 1'h0;
    429: T492 = 1'h0;
    430: T492 = 1'h0;
    431: T492 = 1'h0;
    432: T492 = 1'h0;
    433: T492 = 1'h0;
    434: T492 = 1'h0;
    435: T492 = 1'h0;
    436: T492 = 1'h0;
    437: T492 = 1'h0;
    438: T492 = 1'h0;
    439: T492 = 1'h0;
    440: T492 = 1'h0;
    441: T492 = 1'h0;
    442: T492 = 1'h0;
    443: T492 = 1'h0;
    444: T492 = 1'h0;
    445: T492 = 1'h0;
    446: T492 = 1'h0;
    447: T492 = 1'h0;
    448: T492 = 1'h0;
    449: T492 = 1'h0;
    450: T492 = 1'h0;
    451: T492 = 1'h0;
    452: T492 = 1'h0;
    453: T492 = 1'h0;
    454: T492 = 1'h0;
    455: T492 = 1'h0;
    456: T492 = 1'h0;
    457: T492 = 1'h0;
    458: T492 = 1'h0;
    459: T492 = 1'h0;
    460: T492 = 1'h0;
    461: T492 = 1'h0;
    462: T492 = 1'h0;
    463: T492 = 1'h0;
    464: T492 = 1'h0;
    465: T492 = 1'h0;
    466: T492 = 1'h0;
    467: T492 = 1'h0;
    468: T492 = 1'h0;
    469: T492 = 1'h0;
    470: T492 = 1'h0;
    471: T492 = 1'h0;
    472: T492 = 1'h0;
    473: T492 = 1'h0;
    474: T492 = 1'h0;
    475: T492 = 1'h0;
    476: T492 = 1'h0;
    477: T492 = 1'h0;
    478: T492 = 1'h0;
    479: T492 = 1'h0;
    480: T492 = 1'h0;
    481: T492 = 1'h0;
    482: T492 = 1'h0;
    483: T492 = 1'h0;
    484: T492 = 1'h0;
    485: T492 = 1'h0;
    486: T492 = 1'h0;
    487: T492 = 1'h0;
    488: T492 = 1'h0;
    489: T492 = 1'h0;
    490: T492 = 1'h0;
    491: T492 = 1'h0;
    492: T492 = 1'h0;
    493: T492 = 1'h0;
    494: T492 = 1'h0;
    495: T492 = 1'h0;
    496: T492 = 1'h0;
    497: T492 = 1'h0;
    498: T492 = 1'h0;
    499: T492 = 1'h0;
    500: T492 = 1'h0;
    501: T492 = 1'h0;
    502: T492 = 1'h0;
    503: T492 = 1'h0;
    504: T492 = 1'h0;
    505: T492 = 1'h0;
    506: T492 = 1'h0;
    507: T492 = 1'h0;
    508: T492 = 1'h0;
    509: T492 = 1'h0;
    510: T492 = 1'h0;
    511: T492 = 1'h0;
    512: T492 = 1'h0;
    513: T492 = 1'h0;
    514: T492 = 1'h0;
    515: T492 = 1'h0;
    516: T492 = 1'h0;
    517: T492 = 1'h0;
    518: T492 = 1'h0;
    519: T492 = 1'h0;
    520: T492 = 1'h0;
    521: T492 = 1'h0;
    522: T492 = 1'h0;
    523: T492 = 1'h0;
    524: T492 = 1'h0;
    525: T492 = 1'h0;
    526: T492 = 1'h0;
    527: T492 = 1'h0;
    528: T492 = 1'h0;
    529: T492 = 1'h0;
    530: T492 = 1'h0;
    531: T492 = 1'h0;
    532: T492 = 1'h0;
    533: T492 = 1'h0;
    534: T492 = 1'h0;
    535: T492 = 1'h0;
    536: T492 = 1'h0;
    537: T492 = 1'h0;
    538: T492 = 1'h0;
    539: T492 = 1'h0;
    540: T492 = 1'h0;
    541: T492 = 1'h0;
    542: T492 = 1'h0;
    543: T492 = 1'h0;
    544: T492 = 1'h0;
    545: T492 = 1'h0;
    546: T492 = 1'h0;
    547: T492 = 1'h0;
    548: T492 = 1'h0;
    549: T492 = 1'h0;
    550: T492 = 1'h0;
    551: T492 = 1'h0;
    552: T492 = 1'h0;
    553: T492 = 1'h0;
    554: T492 = 1'h0;
    555: T492 = 1'h0;
    556: T492 = 1'h0;
    557: T492 = 1'h0;
    558: T492 = 1'h0;
    559: T492 = 1'h0;
    560: T492 = 1'h0;
    561: T492 = 1'h0;
    562: T492 = 1'h0;
    563: T492 = 1'h0;
    564: T492 = 1'h0;
    565: T492 = 1'h0;
    566: T492 = 1'h0;
    567: T492 = 1'h0;
    568: T492 = 1'h0;
    569: T492 = 1'h0;
    570: T492 = 1'h0;
    571: T492 = 1'h0;
    572: T492 = 1'h0;
    573: T492 = 1'h0;
    574: T492 = 1'h0;
    575: T492 = 1'h0;
    576: T492 = 1'h0;
    577: T492 = 1'h0;
    578: T492 = 1'h0;
    579: T492 = 1'h0;
    580: T492 = 1'h0;
    581: T492 = 1'h0;
    582: T492 = 1'h0;
    583: T492 = 1'h0;
    584: T492 = 1'h0;
    585: T492 = 1'h0;
    586: T492 = 1'h0;
    587: T492 = 1'h0;
    588: T492 = 1'h0;
    589: T492 = 1'h0;
    590: T492 = 1'h0;
    591: T492 = 1'h0;
    592: T492 = 1'h0;
    593: T492 = 1'h0;
    594: T492 = 1'h0;
    595: T492 = 1'h0;
    596: T492 = 1'h0;
    597: T492 = 1'h0;
    598: T492 = 1'h0;
    599: T492 = 1'h0;
    600: T492 = 1'h0;
    601: T492 = 1'h0;
    602: T492 = 1'h0;
    603: T492 = 1'h0;
    604: T492 = 1'h0;
    605: T492 = 1'h0;
    606: T492 = 1'h0;
    607: T492 = 1'h0;
    608: T492 = 1'h0;
    609: T492 = 1'h0;
    610: T492 = 1'h0;
    611: T492 = 1'h0;
    612: T492 = 1'h0;
    613: T492 = 1'h0;
    614: T492 = 1'h0;
    615: T492 = 1'h0;
    616: T492 = 1'h0;
    617: T492 = 1'h0;
    618: T492 = 1'h0;
    619: T492 = 1'h0;
    620: T492 = 1'h0;
    621: T492 = 1'h0;
    622: T492 = 1'h0;
    623: T492 = 1'h0;
    624: T492 = 1'h0;
    625: T492 = 1'h0;
    626: T492 = 1'h0;
    627: T492 = 1'h0;
    628: T492 = 1'h0;
    629: T492 = 1'h0;
    630: T492 = 1'h0;
    631: T492 = 1'h0;
    632: T492 = 1'h0;
    633: T492 = 1'h0;
    634: T492 = 1'h0;
    635: T492 = 1'h0;
    636: T492 = 1'h0;
    637: T492 = 1'h0;
    638: T492 = 1'h0;
    639: T492 = 1'h0;
    640: T492 = 1'h0;
    641: T492 = 1'h0;
    642: T492 = 1'h0;
    643: T492 = 1'h0;
    644: T492 = 1'h0;
    645: T492 = 1'h0;
    646: T492 = 1'h0;
    647: T492 = 1'h0;
    648: T492 = 1'h0;
    649: T492 = 1'h0;
    650: T492 = 1'h0;
    651: T492 = 1'h0;
    652: T492 = 1'h0;
    653: T492 = 1'h0;
    654: T492 = 1'h0;
    655: T492 = 1'h0;
    656: T492 = 1'h0;
    657: T492 = 1'h0;
    658: T492 = 1'h0;
    659: T492 = 1'h0;
    660: T492 = 1'h0;
    661: T492 = 1'h0;
    662: T492 = 1'h0;
    663: T492 = 1'h0;
    664: T492 = 1'h0;
    665: T492 = 1'h0;
    666: T492 = 1'h0;
    667: T492 = 1'h0;
    668: T492 = 1'h0;
    669: T492 = 1'h0;
    670: T492 = 1'h0;
    671: T492 = 1'h0;
    672: T492 = 1'h0;
    673: T492 = 1'h0;
    674: T492 = 1'h0;
    675: T492 = 1'h0;
    676: T492 = 1'h0;
    677: T492 = 1'h0;
    678: T492 = 1'h0;
    679: T492 = 1'h0;
    680: T492 = 1'h0;
    681: T492 = 1'h0;
    682: T492 = 1'h0;
    683: T492 = 1'h0;
    684: T492 = 1'h0;
    685: T492 = 1'h0;
    686: T492 = 1'h0;
    687: T492 = 1'h0;
    688: T492 = 1'h0;
    689: T492 = 1'h0;
    690: T492 = 1'h0;
    691: T492 = 1'h0;
    692: T492 = 1'h0;
    693: T492 = 1'h0;
    694: T492 = 1'h0;
    695: T492 = 1'h0;
    696: T492 = 1'h0;
    697: T492 = 1'h0;
    698: T492 = 1'h0;
    699: T492 = 1'h0;
    700: T492 = 1'h0;
    701: T492 = 1'h0;
    702: T492 = 1'h0;
    703: T492 = 1'h0;
    704: T492 = 1'h0;
    705: T492 = 1'h0;
    706: T492 = 1'h0;
    707: T492 = 1'h0;
    708: T492 = 1'h0;
    709: T492 = 1'h0;
    710: T492 = 1'h0;
    711: T492 = 1'h0;
    712: T492 = 1'h0;
    713: T492 = 1'h0;
    714: T492 = 1'h0;
    715: T492 = 1'h0;
    716: T492 = 1'h0;
    717: T492 = 1'h0;
    718: T492 = 1'h0;
    719: T492 = 1'h0;
    720: T492 = 1'h0;
    721: T492 = 1'h0;
    722: T492 = 1'h0;
    723: T492 = 1'h0;
    724: T492 = 1'h0;
    725: T492 = 1'h0;
    726: T492 = 1'h0;
    727: T492 = 1'h0;
    728: T492 = 1'h0;
    729: T492 = 1'h0;
    730: T492 = 1'h0;
    731: T492 = 1'h0;
    732: T492 = 1'h0;
    733: T492 = 1'h0;
    734: T492 = 1'h0;
    735: T492 = 1'h0;
    736: T492 = 1'h0;
    737: T492 = 1'h0;
    738: T492 = 1'h0;
    739: T492 = 1'h0;
    740: T492 = 1'h0;
    741: T492 = 1'h0;
    742: T492 = 1'h0;
    743: T492 = 1'h0;
    744: T492 = 1'h0;
    745: T492 = 1'h0;
    746: T492 = 1'h0;
    747: T492 = 1'h0;
    748: T492 = 1'h0;
    749: T492 = 1'h0;
    750: T492 = 1'h0;
    751: T492 = 1'h0;
    752: T492 = 1'h0;
    753: T492 = 1'h0;
    754: T492 = 1'h0;
    755: T492 = 1'h0;
    756: T492 = 1'h0;
    757: T492 = 1'h0;
    758: T492 = 1'h0;
    759: T492 = 1'h0;
    760: T492 = 1'h0;
    761: T492 = 1'h0;
    762: T492 = 1'h0;
    763: T492 = 1'h0;
    764: T492 = 1'h0;
    765: T492 = 1'h0;
    766: T492 = 1'h0;
    767: T492 = 1'h0;
    768: T492 = 1'h0;
    769: T492 = 1'h0;
    770: T492 = 1'h0;
    771: T492 = 1'h0;
    772: T492 = 1'h0;
    773: T492 = 1'h0;
    774: T492 = 1'h0;
    775: T492 = 1'h0;
    776: T492 = 1'h0;
    777: T492 = 1'h0;
    778: T492 = 1'h0;
    779: T492 = 1'h0;
    780: T492 = 1'h0;
    781: T492 = 1'h0;
    782: T492 = 1'h0;
    783: T492 = 1'h0;
    784: T492 = 1'h0;
    785: T492 = 1'h0;
    786: T492 = 1'h0;
    787: T492 = 1'h0;
    788: T492 = 1'h0;
    789: T492 = 1'h0;
    790: T492 = 1'h0;
    791: T492 = 1'h0;
    792: T492 = 1'h0;
    793: T492 = 1'h0;
    794: T492 = 1'h0;
    795: T492 = 1'h0;
    796: T492 = 1'h0;
    797: T492 = 1'h0;
    798: T492 = 1'h0;
    799: T492 = 1'h0;
    800: T492 = 1'h0;
    801: T492 = 1'h0;
    802: T492 = 1'h0;
    803: T492 = 1'h0;
    804: T492 = 1'h0;
    805: T492 = 1'h0;
    806: T492 = 1'h0;
    807: T492 = 1'h0;
    808: T492 = 1'h0;
    809: T492 = 1'h0;
    810: T492 = 1'h0;
    811: T492 = 1'h0;
    812: T492 = 1'h0;
    813: T492 = 1'h0;
    814: T492 = 1'h0;
    815: T492 = 1'h0;
    816: T492 = 1'h0;
    817: T492 = 1'h0;
    818: T492 = 1'h0;
    819: T492 = 1'h0;
    820: T492 = 1'h0;
    821: T492 = 1'h0;
    822: T492 = 1'h0;
    823: T492 = 1'h0;
    824: T492 = 1'h0;
    825: T492 = 1'h0;
    826: T492 = 1'h0;
    827: T492 = 1'h0;
    828: T492 = 1'h0;
    829: T492 = 1'h0;
    830: T492 = 1'h0;
    831: T492 = 1'h0;
    832: T492 = 1'h0;
    833: T492 = 1'h0;
    834: T492 = 1'h0;
    835: T492 = 1'h0;
    836: T492 = 1'h0;
    837: T492 = 1'h0;
    838: T492 = 1'h0;
    839: T492 = 1'h0;
    840: T492 = 1'h0;
    841: T492 = 1'h0;
    842: T492 = 1'h0;
    843: T492 = 1'h0;
    844: T492 = 1'h0;
    845: T492 = 1'h0;
    846: T492 = 1'h0;
    847: T492 = 1'h0;
    848: T492 = 1'h0;
    849: T492 = 1'h0;
    850: T492 = 1'h0;
    851: T492 = 1'h0;
    852: T492 = 1'h0;
    853: T492 = 1'h0;
    854: T492 = 1'h0;
    855: T492 = 1'h0;
    856: T492 = 1'h0;
    857: T492 = 1'h0;
    858: T492 = 1'h0;
    859: T492 = 1'h0;
    860: T492 = 1'h0;
    861: T492 = 1'h0;
    862: T492 = 1'h0;
    863: T492 = 1'h0;
    864: T492 = 1'h0;
    865: T492 = 1'h0;
    866: T492 = 1'h0;
    867: T492 = 1'h0;
    868: T492 = 1'h0;
    869: T492 = 1'h0;
    870: T492 = 1'h0;
    871: T492 = 1'h0;
    872: T492 = 1'h0;
    873: T492 = 1'h0;
    874: T492 = 1'h0;
    875: T492 = 1'h0;
    876: T492 = 1'h0;
    877: T492 = 1'h0;
    878: T492 = 1'h0;
    879: T492 = 1'h0;
    880: T492 = 1'h0;
    881: T492 = 1'h0;
    882: T492 = 1'h0;
    883: T492 = 1'h0;
    884: T492 = 1'h0;
    885: T492 = 1'h0;
    886: T492 = 1'h0;
    887: T492 = 1'h0;
    888: T492 = 1'h0;
    889: T492 = 1'h0;
    890: T492 = 1'h0;
    891: T492 = 1'h0;
    892: T492 = 1'h0;
    893: T492 = 1'h0;
    894: T492 = 1'h0;
    895: T492 = 1'h0;
    896: T492 = 1'h0;
    897: T492 = 1'h0;
    898: T492 = 1'h0;
    899: T492 = 1'h0;
    900: T492 = 1'h0;
    901: T492 = 1'h0;
    902: T492 = 1'h0;
    903: T492 = 1'h0;
    904: T492 = 1'h0;
    905: T492 = 1'h0;
    906: T492 = 1'h0;
    907: T492 = 1'h0;
    908: T492 = 1'h0;
    909: T492 = 1'h0;
    910: T492 = 1'h0;
    911: T492 = 1'h0;
    912: T492 = 1'h0;
    913: T492 = 1'h0;
    914: T492 = 1'h0;
    915: T492 = 1'h0;
    916: T492 = 1'h0;
    917: T492 = 1'h0;
    918: T492 = 1'h0;
    919: T492 = 1'h0;
    920: T492 = 1'h0;
    921: T492 = 1'h0;
    922: T492 = 1'h0;
    923: T492 = 1'h0;
    924: T492 = 1'h0;
    925: T492 = 1'h0;
    926: T492 = 1'h0;
    927: T492 = 1'h0;
    928: T492 = 1'h0;
    929: T492 = 1'h0;
    930: T492 = 1'h0;
    931: T492 = 1'h0;
    932: T492 = 1'h0;
    933: T492 = 1'h0;
    934: T492 = 1'h0;
    935: T492 = 1'h0;
    936: T492 = 1'h0;
    937: T492 = 1'h0;
    938: T492 = 1'h0;
    939: T492 = 1'h0;
    940: T492 = 1'h0;
    941: T492 = 1'h0;
    942: T492 = 1'h0;
    943: T492 = 1'h0;
    944: T492 = 1'h0;
    945: T492 = 1'h0;
    946: T492 = 1'h0;
    947: T492 = 1'h0;
    948: T492 = 1'h0;
    949: T492 = 1'h0;
    950: T492 = 1'h0;
    951: T492 = 1'h0;
    952: T492 = 1'h0;
    953: T492 = 1'h0;
    954: T492 = 1'h0;
    955: T492 = 1'h0;
    956: T492 = 1'h0;
    957: T492 = 1'h0;
    958: T492 = 1'h0;
    959: T492 = 1'h0;
    960: T492 = 1'h0;
    961: T492 = 1'h0;
    962: T492 = 1'h0;
    963: T492 = 1'h0;
    964: T492 = 1'h0;
    965: T492 = 1'h0;
    966: T492 = 1'h0;
    967: T492 = 1'h0;
    968: T492 = 1'h0;
    969: T492 = 1'h0;
    970: T492 = 1'h0;
    971: T492 = 1'h0;
    972: T492 = 1'h0;
    973: T492 = 1'h0;
    974: T492 = 1'h0;
    975: T492 = 1'h0;
    976: T492 = 1'h0;
    977: T492 = 1'h0;
    978: T492 = 1'h0;
    979: T492 = 1'h0;
    980: T492 = 1'h0;
    981: T492 = 1'h0;
    982: T492 = 1'h0;
    983: T492 = 1'h0;
    984: T492 = 1'h0;
    985: T492 = 1'h0;
    986: T492 = 1'h0;
    987: T492 = 1'h0;
    988: T492 = 1'h0;
    989: T492 = 1'h0;
    990: T492 = 1'h0;
    991: T492 = 1'h0;
    992: T492 = 1'h0;
    993: T492 = 1'h0;
    994: T492 = 1'h0;
    995: T492 = 1'h0;
    996: T492 = 1'h0;
    997: T492 = 1'h0;
    998: T492 = 1'h0;
    999: T492 = 1'h0;
    1000: T492 = 1'h0;
    1001: T492 = 1'h0;
    1002: T492 = 1'h0;
    1003: T492 = 1'h0;
    1004: T492 = 1'h0;
    1005: T492 = 1'h0;
    1006: T492 = 1'h0;
    1007: T492 = 1'h0;
    1008: T492 = 1'h0;
    1009: T492 = 1'h0;
    1010: T492 = 1'h0;
    1011: T492 = 1'h0;
    1012: T492 = 1'h0;
    1013: T492 = 1'h0;
    1014: T492 = 1'h0;
    1015: T492 = 1'h0;
    1016: T492 = 1'h0;
    1017: T492 = 1'h0;
    1018: T492 = 1'h0;
    1019: T492 = 1'h0;
    1020: T492 = 1'h0;
    1021: T492 = 1'h0;
    1022: T492 = 1'h0;
    1023: T492 = 1'h0;
    1024: T492 = 1'h0;
    1025: T492 = 1'h0;
    1026: T492 = 1'h0;
    1027: T492 = 1'h0;
    1028: T492 = 1'h0;
    1029: T492 = 1'h0;
    1030: T492 = 1'h0;
    1031: T492 = 1'h0;
    1032: T492 = 1'h0;
    1033: T492 = 1'h0;
    1034: T492 = 1'h0;
    1035: T492 = 1'h0;
    1036: T492 = 1'h0;
    1037: T492 = 1'h0;
    1038: T492 = 1'h0;
    1039: T492 = 1'h0;
    1040: T492 = 1'h0;
    1041: T492 = 1'h0;
    1042: T492 = 1'h0;
    1043: T492 = 1'h0;
    1044: T492 = 1'h0;
    1045: T492 = 1'h0;
    1046: T492 = 1'h0;
    1047: T492 = 1'h0;
    1048: T492 = 1'h0;
    1049: T492 = 1'h0;
    1050: T492 = 1'h0;
    1051: T492 = 1'h0;
    1052: T492 = 1'h0;
    1053: T492 = 1'h0;
    1054: T492 = 1'h0;
    1055: T492 = 1'h0;
    1056: T492 = 1'h0;
    1057: T492 = 1'h0;
    1058: T492 = 1'h0;
    1059: T492 = 1'h0;
    1060: T492 = 1'h0;
    1061: T492 = 1'h0;
    1062: T492 = 1'h0;
    1063: T492 = 1'h0;
    1064: T492 = 1'h0;
    1065: T492 = 1'h0;
    1066: T492 = 1'h0;
    1067: T492 = 1'h0;
    1068: T492 = 1'h0;
    1069: T492 = 1'h0;
    1070: T492 = 1'h0;
    1071: T492 = 1'h0;
    1072: T492 = 1'h0;
    1073: T492 = 1'h0;
    1074: T492 = 1'h0;
    1075: T492 = 1'h0;
    1076: T492 = 1'h0;
    1077: T492 = 1'h0;
    1078: T492 = 1'h0;
    1079: T492 = 1'h0;
    1080: T492 = 1'h0;
    1081: T492 = 1'h0;
    1082: T492 = 1'h0;
    1083: T492 = 1'h0;
    1084: T492 = 1'h0;
    1085: T492 = 1'h0;
    1086: T492 = 1'h0;
    1087: T492 = 1'h0;
    1088: T492 = 1'h0;
    1089: T492 = 1'h0;
    1090: T492 = 1'h0;
    1091: T492 = 1'h0;
    1092: T492 = 1'h0;
    1093: T492 = 1'h0;
    1094: T492 = 1'h0;
    1095: T492 = 1'h0;
    1096: T492 = 1'h0;
    1097: T492 = 1'h0;
    1098: T492 = 1'h0;
    1099: T492 = 1'h0;
    1100: T492 = 1'h0;
    1101: T492 = 1'h0;
    1102: T492 = 1'h0;
    1103: T492 = 1'h0;
    1104: T492 = 1'h0;
    1105: T492 = 1'h0;
    1106: T492 = 1'h0;
    1107: T492 = 1'h0;
    1108: T492 = 1'h0;
    1109: T492 = 1'h0;
    1110: T492 = 1'h0;
    1111: T492 = 1'h0;
    1112: T492 = 1'h0;
    1113: T492 = 1'h0;
    1114: T492 = 1'h0;
    1115: T492 = 1'h0;
    1116: T492 = 1'h0;
    1117: T492 = 1'h0;
    1118: T492 = 1'h0;
    1119: T492 = 1'h0;
    1120: T492 = 1'h0;
    1121: T492 = 1'h0;
    1122: T492 = 1'h0;
    1123: T492 = 1'h0;
    1124: T492 = 1'h0;
    1125: T492 = 1'h0;
    1126: T492 = 1'h0;
    1127: T492 = 1'h0;
    1128: T492 = 1'h0;
    1129: T492 = 1'h0;
    1130: T492 = 1'h0;
    1131: T492 = 1'h0;
    1132: T492 = 1'h0;
    1133: T492 = 1'h0;
    1134: T492 = 1'h0;
    1135: T492 = 1'h0;
    1136: T492 = 1'h0;
    1137: T492 = 1'h0;
    1138: T492 = 1'h0;
    1139: T492 = 1'h0;
    1140: T492 = 1'h0;
    1141: T492 = 1'h0;
    1142: T492 = 1'h0;
    1143: T492 = 1'h0;
    1144: T492 = 1'h0;
    1145: T492 = 1'h0;
    1146: T492 = 1'h0;
    1147: T492 = 1'h0;
    1148: T492 = 1'h0;
    1149: T492 = 1'h0;
    1150: T492 = 1'h0;
    1151: T492 = 1'h0;
    1152: T492 = 1'h0;
    1153: T492 = 1'h0;
    1154: T492 = 1'h0;
    1155: T492 = 1'h0;
    1156: T492 = 1'h0;
    1157: T492 = 1'h0;
    1158: T492 = 1'h0;
    1159: T492 = 1'h0;
    1160: T492 = 1'h0;
    1161: T492 = 1'h0;
    1162: T492 = 1'h0;
    1163: T492 = 1'h0;
    1164: T492 = 1'h0;
    1165: T492 = 1'h0;
    1166: T492 = 1'h0;
    1167: T492 = 1'h0;
    1168: T492 = 1'h0;
    1169: T492 = 1'h0;
    1170: T492 = 1'h0;
    1171: T492 = 1'h0;
    1172: T492 = 1'h0;
    1173: T492 = 1'h0;
    1174: T492 = 1'h0;
    1175: T492 = 1'h0;
    1176: T492 = 1'h0;
    1177: T492 = 1'h0;
    1178: T492 = 1'h0;
    1179: T492 = 1'h0;
    1180: T492 = 1'h0;
    1181: T492 = 1'h0;
    1182: T492 = 1'h0;
    1183: T492 = 1'h0;
    1184: T492 = 1'h0;
    1185: T492 = 1'h0;
    1186: T492 = 1'h0;
    1187: T492 = 1'h0;
    1188: T492 = 1'h0;
    1189: T492 = 1'h0;
    1190: T492 = 1'h0;
    1191: T492 = 1'h0;
    1192: T492 = 1'h0;
    1193: T492 = 1'h0;
    1194: T492 = 1'h0;
    1195: T492 = 1'h0;
    1196: T492 = 1'h0;
    1197: T492 = 1'h0;
    1198: T492 = 1'h0;
    1199: T492 = 1'h0;
    1200: T492 = 1'h0;
    1201: T492 = 1'h0;
    1202: T492 = 1'h0;
    1203: T492 = 1'h0;
    1204: T492 = 1'h0;
    1205: T492 = 1'h0;
    1206: T492 = 1'h0;
    1207: T492 = 1'h0;
    1208: T492 = 1'h0;
    1209: T492 = 1'h0;
    1210: T492 = 1'h0;
    1211: T492 = 1'h0;
    1212: T492 = 1'h0;
    1213: T492 = 1'h0;
    1214: T492 = 1'h0;
    1215: T492 = 1'h0;
    1216: T492 = 1'h0;
    1217: T492 = 1'h0;
    1218: T492 = 1'h0;
    1219: T492 = 1'h0;
    1220: T492 = 1'h0;
    1221: T492 = 1'h0;
    1222: T492 = 1'h0;
    1223: T492 = 1'h0;
    1224: T492 = 1'h0;
    1225: T492 = 1'h0;
    1226: T492 = 1'h0;
    1227: T492 = 1'h0;
    1228: T492 = 1'h0;
    1229: T492 = 1'h0;
    1230: T492 = 1'h0;
    1231: T492 = 1'h0;
    1232: T492 = 1'h0;
    1233: T492 = 1'h0;
    1234: T492 = 1'h0;
    1235: T492 = 1'h0;
    1236: T492 = 1'h0;
    1237: T492 = 1'h0;
    1238: T492 = 1'h0;
    1239: T492 = 1'h0;
    1240: T492 = 1'h0;
    1241: T492 = 1'h0;
    1242: T492 = 1'h0;
    1243: T492 = 1'h0;
    1244: T492 = 1'h0;
    1245: T492 = 1'h0;
    1246: T492 = 1'h0;
    1247: T492 = 1'h0;
    1248: T492 = 1'h0;
    1249: T492 = 1'h0;
    1250: T492 = 1'h0;
    1251: T492 = 1'h0;
    1252: T492 = 1'h0;
    1253: T492 = 1'h0;
    1254: T492 = 1'h0;
    1255: T492 = 1'h0;
    1256: T492 = 1'h0;
    1257: T492 = 1'h0;
    1258: T492 = 1'h0;
    1259: T492 = 1'h0;
    1260: T492 = 1'h0;
    1261: T492 = 1'h0;
    1262: T492 = 1'h0;
    1263: T492 = 1'h0;
    1264: T492 = 1'h0;
    1265: T492 = 1'h0;
    1266: T492 = 1'h0;
    1267: T492 = 1'h0;
    1268: T492 = 1'h0;
    1269: T492 = 1'h0;
    1270: T492 = 1'h0;
    1271: T492 = 1'h0;
    1272: T492 = 1'h0;
    1273: T492 = 1'h0;
    1274: T492 = 1'h0;
    1275: T492 = 1'h0;
    1276: T492 = 1'h0;
    1277: T492 = 1'h0;
    1278: T492 = 1'h0;
    1279: T492 = 1'h0;
    1280: T492 = 1'h1;
    1281: T492 = 1'h1;
    1282: T492 = 1'h1;
    1283: T492 = 1'h1;
    1284: T492 = 1'h1;
    1285: T492 = 1'h1;
    1286: T492 = 1'h1;
    1287: T492 = 1'h1;
    1288: T492 = 1'h1;
    1289: T492 = 1'h1;
    1290: T492 = 1'h1;
    1291: T492 = 1'h1;
    1292: T492 = 1'h1;
    1293: T492 = 1'h1;
    1294: T492 = 1'h1;
    1295: T492 = 1'h1;
    1296: T492 = 1'h0;
    1297: T492 = 1'h0;
    1298: T492 = 1'h0;
    1299: T492 = 1'h0;
    1300: T492 = 1'h0;
    1301: T492 = 1'h0;
    1302: T492 = 1'h0;
    1303: T492 = 1'h0;
    1304: T492 = 1'h0;
    1305: T492 = 1'h0;
    1306: T492 = 1'h0;
    1307: T492 = 1'h0;
    1308: T492 = 1'h0;
    1309: T492 = 1'h1;
    1310: T492 = 1'h1;
    1311: T492 = 1'h1;
    1312: T492 = 1'h1;
    1313: T492 = 1'h1;
    1314: T492 = 1'h1;
    1315: T492 = 1'h1;
    1316: T492 = 1'h0;
    1317: T492 = 1'h0;
    1318: T492 = 1'h0;
    1319: T492 = 1'h0;
    1320: T492 = 1'h0;
    1321: T492 = 1'h0;
    1322: T492 = 1'h0;
    1323: T492 = 1'h0;
    1324: T492 = 1'h0;
    1325: T492 = 1'h0;
    1326: T492 = 1'h0;
    1327: T492 = 1'h0;
    1328: T492 = 1'h0;
    1329: T492 = 1'h0;
    1330: T492 = 1'h0;
    1331: T492 = 1'h0;
    1332: T492 = 1'h0;
    1333: T492 = 1'h0;
    1334: T492 = 1'h0;
    1335: T492 = 1'h0;
    1336: T492 = 1'h0;
    1337: T492 = 1'h0;
    1338: T492 = 1'h0;
    1339: T492 = 1'h0;
    1340: T492 = 1'h0;
    1341: T492 = 1'h0;
    1342: T492 = 1'h0;
    1343: T492 = 1'h0;
    1344: T492 = 1'h0;
    1345: T492 = 1'h0;
    1346: T492 = 1'h0;
    1347: T492 = 1'h0;
    1348: T492 = 1'h0;
    1349: T492 = 1'h0;
    1350: T492 = 1'h0;
    1351: T492 = 1'h0;
    1352: T492 = 1'h0;
    1353: T492 = 1'h0;
    1354: T492 = 1'h0;
    1355: T492 = 1'h0;
    1356: T492 = 1'h0;
    1357: T492 = 1'h0;
    1358: T492 = 1'h0;
    1359: T492 = 1'h0;
    1360: T492 = 1'h0;
    1361: T492 = 1'h0;
    1362: T492 = 1'h0;
    1363: T492 = 1'h0;
    1364: T492 = 1'h0;
    1365: T492 = 1'h0;
    1366: T492 = 1'h0;
    1367: T492 = 1'h0;
    1368: T492 = 1'h0;
    1369: T492 = 1'h0;
    1370: T492 = 1'h0;
    1371: T492 = 1'h0;
    1372: T492 = 1'h0;
    1373: T492 = 1'h0;
    1374: T492 = 1'h0;
    1375: T492 = 1'h0;
    1376: T492 = 1'h0;
    1377: T492 = 1'h0;
    1378: T492 = 1'h0;
    1379: T492 = 1'h0;
    1380: T492 = 1'h0;
    1381: T492 = 1'h0;
    1382: T492 = 1'h0;
    1383: T492 = 1'h0;
    1384: T492 = 1'h0;
    1385: T492 = 1'h0;
    1386: T492 = 1'h0;
    1387: T492 = 1'h0;
    1388: T492 = 1'h0;
    1389: T492 = 1'h0;
    1390: T492 = 1'h0;
    1391: T492 = 1'h0;
    1392: T492 = 1'h0;
    1393: T492 = 1'h0;
    1394: T492 = 1'h0;
    1395: T492 = 1'h0;
    1396: T492 = 1'h0;
    1397: T492 = 1'h0;
    1398: T492 = 1'h0;
    1399: T492 = 1'h0;
    1400: T492 = 1'h0;
    1401: T492 = 1'h0;
    1402: T492 = 1'h0;
    1403: T492 = 1'h0;
    1404: T492 = 1'h0;
    1405: T492 = 1'h0;
    1406: T492 = 1'h0;
    1407: T492 = 1'h0;
    1408: T492 = 1'h0;
    1409: T492 = 1'h0;
    1410: T492 = 1'h0;
    1411: T492 = 1'h0;
    1412: T492 = 1'h0;
    1413: T492 = 1'h0;
    1414: T492 = 1'h0;
    1415: T492 = 1'h0;
    1416: T492 = 1'h0;
    1417: T492 = 1'h0;
    1418: T492 = 1'h0;
    1419: T492 = 1'h0;
    1420: T492 = 1'h0;
    1421: T492 = 1'h0;
    1422: T492 = 1'h0;
    1423: T492 = 1'h0;
    1424: T492 = 1'h0;
    1425: T492 = 1'h0;
    1426: T492 = 1'h0;
    1427: T492 = 1'h0;
    1428: T492 = 1'h0;
    1429: T492 = 1'h0;
    1430: T492 = 1'h0;
    1431: T492 = 1'h0;
    1432: T492 = 1'h0;
    1433: T492 = 1'h0;
    1434: T492 = 1'h0;
    1435: T492 = 1'h0;
    1436: T492 = 1'h0;
    1437: T492 = 1'h0;
    1438: T492 = 1'h0;
    1439: T492 = 1'h0;
    1440: T492 = 1'h0;
    1441: T492 = 1'h0;
    1442: T492 = 1'h0;
    1443: T492 = 1'h0;
    1444: T492 = 1'h0;
    1445: T492 = 1'h0;
    1446: T492 = 1'h0;
    1447: T492 = 1'h0;
    1448: T492 = 1'h0;
    1449: T492 = 1'h0;
    1450: T492 = 1'h0;
    1451: T492 = 1'h0;
    1452: T492 = 1'h0;
    1453: T492 = 1'h0;
    1454: T492 = 1'h0;
    1455: T492 = 1'h0;
    1456: T492 = 1'h0;
    1457: T492 = 1'h0;
    1458: T492 = 1'h0;
    1459: T492 = 1'h0;
    1460: T492 = 1'h0;
    1461: T492 = 1'h0;
    1462: T492 = 1'h0;
    1463: T492 = 1'h0;
    1464: T492 = 1'h0;
    1465: T492 = 1'h0;
    1466: T492 = 1'h0;
    1467: T492 = 1'h0;
    1468: T492 = 1'h0;
    1469: T492 = 1'h0;
    1470: T492 = 1'h0;
    1471: T492 = 1'h0;
    1472: T492 = 1'h0;
    1473: T492 = 1'h0;
    1474: T492 = 1'h0;
    1475: T492 = 1'h0;
    1476: T492 = 1'h0;
    1477: T492 = 1'h0;
    1478: T492 = 1'h0;
    1479: T492 = 1'h0;
    1480: T492 = 1'h0;
    1481: T492 = 1'h0;
    1482: T492 = 1'h0;
    1483: T492 = 1'h0;
    1484: T492 = 1'h0;
    1485: T492 = 1'h0;
    1486: T492 = 1'h0;
    1487: T492 = 1'h0;
    1488: T492 = 1'h0;
    1489: T492 = 1'h0;
    1490: T492 = 1'h0;
    1491: T492 = 1'h0;
    1492: T492 = 1'h0;
    1493: T492 = 1'h0;
    1494: T492 = 1'h0;
    1495: T492 = 1'h0;
    1496: T492 = 1'h0;
    1497: T492 = 1'h0;
    1498: T492 = 1'h0;
    1499: T492 = 1'h0;
    1500: T492 = 1'h0;
    1501: T492 = 1'h0;
    1502: T492 = 1'h0;
    1503: T492 = 1'h0;
    1504: T492 = 1'h0;
    1505: T492 = 1'h0;
    1506: T492 = 1'h0;
    1507: T492 = 1'h0;
    1508: T492 = 1'h0;
    1509: T492 = 1'h0;
    1510: T492 = 1'h0;
    1511: T492 = 1'h0;
    1512: T492 = 1'h0;
    1513: T492 = 1'h0;
    1514: T492 = 1'h0;
    1515: T492 = 1'h0;
    1516: T492 = 1'h0;
    1517: T492 = 1'h0;
    1518: T492 = 1'h0;
    1519: T492 = 1'h0;
    1520: T492 = 1'h0;
    1521: T492 = 1'h0;
    1522: T492 = 1'h0;
    1523: T492 = 1'h0;
    1524: T492 = 1'h0;
    1525: T492 = 1'h0;
    1526: T492 = 1'h0;
    1527: T492 = 1'h0;
    1528: T492 = 1'h0;
    1529: T492 = 1'h0;
    1530: T492 = 1'h0;
    1531: T492 = 1'h0;
    1532: T492 = 1'h0;
    1533: T492 = 1'h0;
    1534: T492 = 1'h0;
    1535: T492 = 1'h0;
    1536: T492 = 1'h0;
    1537: T492 = 1'h0;
    1538: T492 = 1'h0;
    1539: T492 = 1'h0;
    1540: T492 = 1'h0;
    1541: T492 = 1'h0;
    1542: T492 = 1'h0;
    1543: T492 = 1'h0;
    1544: T492 = 1'h0;
    1545: T492 = 1'h0;
    1546: T492 = 1'h0;
    1547: T492 = 1'h0;
    1548: T492 = 1'h0;
    1549: T492 = 1'h0;
    1550: T492 = 1'h0;
    1551: T492 = 1'h0;
    1552: T492 = 1'h0;
    1553: T492 = 1'h0;
    1554: T492 = 1'h0;
    1555: T492 = 1'h0;
    1556: T492 = 1'h0;
    1557: T492 = 1'h0;
    1558: T492 = 1'h0;
    1559: T492 = 1'h0;
    1560: T492 = 1'h0;
    1561: T492 = 1'h0;
    1562: T492 = 1'h0;
    1563: T492 = 1'h0;
    1564: T492 = 1'h0;
    1565: T492 = 1'h0;
    1566: T492 = 1'h0;
    1567: T492 = 1'h0;
    1568: T492 = 1'h0;
    1569: T492 = 1'h0;
    1570: T492 = 1'h0;
    1571: T492 = 1'h0;
    1572: T492 = 1'h0;
    1573: T492 = 1'h0;
    1574: T492 = 1'h0;
    1575: T492 = 1'h0;
    1576: T492 = 1'h0;
    1577: T492 = 1'h0;
    1578: T492 = 1'h0;
    1579: T492 = 1'h0;
    1580: T492 = 1'h0;
    1581: T492 = 1'h0;
    1582: T492 = 1'h0;
    1583: T492 = 1'h0;
    1584: T492 = 1'h0;
    1585: T492 = 1'h0;
    1586: T492 = 1'h0;
    1587: T492 = 1'h0;
    1588: T492 = 1'h0;
    1589: T492 = 1'h0;
    1590: T492 = 1'h0;
    1591: T492 = 1'h0;
    1592: T492 = 1'h0;
    1593: T492 = 1'h0;
    1594: T492 = 1'h0;
    1595: T492 = 1'h0;
    1596: T492 = 1'h0;
    1597: T492 = 1'h0;
    1598: T492 = 1'h0;
    1599: T492 = 1'h0;
    1600: T492 = 1'h0;
    1601: T492 = 1'h0;
    1602: T492 = 1'h0;
    1603: T492 = 1'h0;
    1604: T492 = 1'h0;
    1605: T492 = 1'h0;
    1606: T492 = 1'h0;
    1607: T492 = 1'h0;
    1608: T492 = 1'h0;
    1609: T492 = 1'h0;
    1610: T492 = 1'h0;
    1611: T492 = 1'h0;
    1612: T492 = 1'h0;
    1613: T492 = 1'h0;
    1614: T492 = 1'h0;
    1615: T492 = 1'h0;
    1616: T492 = 1'h0;
    1617: T492 = 1'h0;
    1618: T492 = 1'h0;
    1619: T492 = 1'h0;
    1620: T492 = 1'h0;
    1621: T492 = 1'h0;
    1622: T492 = 1'h0;
    1623: T492 = 1'h0;
    1624: T492 = 1'h0;
    1625: T492 = 1'h0;
    1626: T492 = 1'h0;
    1627: T492 = 1'h0;
    1628: T492 = 1'h0;
    1629: T492 = 1'h0;
    1630: T492 = 1'h0;
    1631: T492 = 1'h0;
    1632: T492 = 1'h0;
    1633: T492 = 1'h0;
    1634: T492 = 1'h0;
    1635: T492 = 1'h0;
    1636: T492 = 1'h0;
    1637: T492 = 1'h0;
    1638: T492 = 1'h0;
    1639: T492 = 1'h0;
    1640: T492 = 1'h0;
    1641: T492 = 1'h0;
    1642: T492 = 1'h0;
    1643: T492 = 1'h0;
    1644: T492 = 1'h0;
    1645: T492 = 1'h0;
    1646: T492 = 1'h0;
    1647: T492 = 1'h0;
    1648: T492 = 1'h0;
    1649: T492 = 1'h0;
    1650: T492 = 1'h0;
    1651: T492 = 1'h0;
    1652: T492 = 1'h0;
    1653: T492 = 1'h0;
    1654: T492 = 1'h0;
    1655: T492 = 1'h0;
    1656: T492 = 1'h0;
    1657: T492 = 1'h0;
    1658: T492 = 1'h0;
    1659: T492 = 1'h0;
    1660: T492 = 1'h0;
    1661: T492 = 1'h0;
    1662: T492 = 1'h0;
    1663: T492 = 1'h0;
    1664: T492 = 1'h0;
    1665: T492 = 1'h0;
    1666: T492 = 1'h0;
    1667: T492 = 1'h0;
    1668: T492 = 1'h0;
    1669: T492 = 1'h0;
    1670: T492 = 1'h0;
    1671: T492 = 1'h0;
    1672: T492 = 1'h0;
    1673: T492 = 1'h0;
    1674: T492 = 1'h0;
    1675: T492 = 1'h0;
    1676: T492 = 1'h0;
    1677: T492 = 1'h0;
    1678: T492 = 1'h0;
    1679: T492 = 1'h0;
    1680: T492 = 1'h0;
    1681: T492 = 1'h0;
    1682: T492 = 1'h0;
    1683: T492 = 1'h0;
    1684: T492 = 1'h0;
    1685: T492 = 1'h0;
    1686: T492 = 1'h0;
    1687: T492 = 1'h0;
    1688: T492 = 1'h0;
    1689: T492 = 1'h0;
    1690: T492 = 1'h0;
    1691: T492 = 1'h0;
    1692: T492 = 1'h0;
    1693: T492 = 1'h0;
    1694: T492 = 1'h0;
    1695: T492 = 1'h0;
    1696: T492 = 1'h0;
    1697: T492 = 1'h0;
    1698: T492 = 1'h0;
    1699: T492 = 1'h0;
    1700: T492 = 1'h0;
    1701: T492 = 1'h0;
    1702: T492 = 1'h0;
    1703: T492 = 1'h0;
    1704: T492 = 1'h0;
    1705: T492 = 1'h0;
    1706: T492 = 1'h0;
    1707: T492 = 1'h0;
    1708: T492 = 1'h0;
    1709: T492 = 1'h0;
    1710: T492 = 1'h0;
    1711: T492 = 1'h0;
    1712: T492 = 1'h0;
    1713: T492 = 1'h0;
    1714: T492 = 1'h0;
    1715: T492 = 1'h0;
    1716: T492 = 1'h0;
    1717: T492 = 1'h0;
    1718: T492 = 1'h0;
    1719: T492 = 1'h0;
    1720: T492 = 1'h0;
    1721: T492 = 1'h0;
    1722: T492 = 1'h0;
    1723: T492 = 1'h0;
    1724: T492 = 1'h0;
    1725: T492 = 1'h0;
    1726: T492 = 1'h0;
    1727: T492 = 1'h0;
    1728: T492 = 1'h0;
    1729: T492 = 1'h0;
    1730: T492 = 1'h0;
    1731: T492 = 1'h0;
    1732: T492 = 1'h0;
    1733: T492 = 1'h0;
    1734: T492 = 1'h0;
    1735: T492 = 1'h0;
    1736: T492 = 1'h0;
    1737: T492 = 1'h0;
    1738: T492 = 1'h0;
    1739: T492 = 1'h0;
    1740: T492 = 1'h0;
    1741: T492 = 1'h0;
    1742: T492 = 1'h0;
    1743: T492 = 1'h0;
    1744: T492 = 1'h0;
    1745: T492 = 1'h0;
    1746: T492 = 1'h0;
    1747: T492 = 1'h0;
    1748: T492 = 1'h0;
    1749: T492 = 1'h0;
    1750: T492 = 1'h0;
    1751: T492 = 1'h0;
    1752: T492 = 1'h0;
    1753: T492 = 1'h0;
    1754: T492 = 1'h0;
    1755: T492 = 1'h0;
    1756: T492 = 1'h0;
    1757: T492 = 1'h0;
    1758: T492 = 1'h0;
    1759: T492 = 1'h0;
    1760: T492 = 1'h0;
    1761: T492 = 1'h0;
    1762: T492 = 1'h0;
    1763: T492 = 1'h0;
    1764: T492 = 1'h0;
    1765: T492 = 1'h0;
    1766: T492 = 1'h0;
    1767: T492 = 1'h0;
    1768: T492 = 1'h0;
    1769: T492 = 1'h0;
    1770: T492 = 1'h0;
    1771: T492 = 1'h0;
    1772: T492 = 1'h0;
    1773: T492 = 1'h0;
    1774: T492 = 1'h0;
    1775: T492 = 1'h0;
    1776: T492 = 1'h0;
    1777: T492 = 1'h0;
    1778: T492 = 1'h0;
    1779: T492 = 1'h0;
    1780: T492 = 1'h0;
    1781: T492 = 1'h0;
    1782: T492 = 1'h0;
    1783: T492 = 1'h0;
    1784: T492 = 1'h0;
    1785: T492 = 1'h0;
    1786: T492 = 1'h0;
    1787: T492 = 1'h0;
    1788: T492 = 1'h0;
    1789: T492 = 1'h0;
    1790: T492 = 1'h0;
    1791: T492 = 1'h0;
    1792: T492 = 1'h0;
    1793: T492 = 1'h0;
    1794: T492 = 1'h0;
    1795: T492 = 1'h0;
    1796: T492 = 1'h0;
    1797: T492 = 1'h0;
    1798: T492 = 1'h0;
    1799: T492 = 1'h0;
    1800: T492 = 1'h0;
    1801: T492 = 1'h0;
    1802: T492 = 1'h0;
    1803: T492 = 1'h0;
    1804: T492 = 1'h0;
    1805: T492 = 1'h0;
    1806: T492 = 1'h0;
    1807: T492 = 1'h0;
    1808: T492 = 1'h0;
    1809: T492 = 1'h0;
    1810: T492 = 1'h0;
    1811: T492 = 1'h0;
    1812: T492 = 1'h0;
    1813: T492 = 1'h0;
    1814: T492 = 1'h0;
    1815: T492 = 1'h0;
    1816: T492 = 1'h0;
    1817: T492 = 1'h0;
    1818: T492 = 1'h0;
    1819: T492 = 1'h0;
    1820: T492 = 1'h0;
    1821: T492 = 1'h0;
    1822: T492 = 1'h0;
    1823: T492 = 1'h0;
    1824: T492 = 1'h0;
    1825: T492 = 1'h0;
    1826: T492 = 1'h0;
    1827: T492 = 1'h0;
    1828: T492 = 1'h0;
    1829: T492 = 1'h0;
    1830: T492 = 1'h0;
    1831: T492 = 1'h0;
    1832: T492 = 1'h0;
    1833: T492 = 1'h0;
    1834: T492 = 1'h0;
    1835: T492 = 1'h0;
    1836: T492 = 1'h0;
    1837: T492 = 1'h0;
    1838: T492 = 1'h0;
    1839: T492 = 1'h0;
    1840: T492 = 1'h0;
    1841: T492 = 1'h0;
    1842: T492 = 1'h0;
    1843: T492 = 1'h0;
    1844: T492 = 1'h0;
    1845: T492 = 1'h0;
    1846: T492 = 1'h0;
    1847: T492 = 1'h0;
    1848: T492 = 1'h0;
    1849: T492 = 1'h0;
    1850: T492 = 1'h0;
    1851: T492 = 1'h0;
    1852: T492 = 1'h0;
    1853: T492 = 1'h0;
    1854: T492 = 1'h0;
    1855: T492 = 1'h0;
    1856: T492 = 1'h0;
    1857: T492 = 1'h0;
    1858: T492 = 1'h0;
    1859: T492 = 1'h0;
    1860: T492 = 1'h0;
    1861: T492 = 1'h0;
    1862: T492 = 1'h0;
    1863: T492 = 1'h0;
    1864: T492 = 1'h0;
    1865: T492 = 1'h0;
    1866: T492 = 1'h0;
    1867: T492 = 1'h0;
    1868: T492 = 1'h0;
    1869: T492 = 1'h0;
    1870: T492 = 1'h0;
    1871: T492 = 1'h0;
    1872: T492 = 1'h0;
    1873: T492 = 1'h0;
    1874: T492 = 1'h0;
    1875: T492 = 1'h0;
    1876: T492 = 1'h0;
    1877: T492 = 1'h0;
    1878: T492 = 1'h0;
    1879: T492 = 1'h0;
    1880: T492 = 1'h0;
    1881: T492 = 1'h0;
    1882: T492 = 1'h0;
    1883: T492 = 1'h0;
    1884: T492 = 1'h0;
    1885: T492 = 1'h0;
    1886: T492 = 1'h0;
    1887: T492 = 1'h0;
    1888: T492 = 1'h0;
    1889: T492 = 1'h0;
    1890: T492 = 1'h0;
    1891: T492 = 1'h0;
    1892: T492 = 1'h0;
    1893: T492 = 1'h0;
    1894: T492 = 1'h0;
    1895: T492 = 1'h0;
    1896: T492 = 1'h0;
    1897: T492 = 1'h0;
    1898: T492 = 1'h0;
    1899: T492 = 1'h0;
    1900: T492 = 1'h0;
    1901: T492 = 1'h0;
    1902: T492 = 1'h0;
    1903: T492 = 1'h0;
    1904: T492 = 1'h0;
    1905: T492 = 1'h0;
    1906: T492 = 1'h0;
    1907: T492 = 1'h0;
    1908: T492 = 1'h0;
    1909: T492 = 1'h0;
    1910: T492 = 1'h0;
    1911: T492 = 1'h0;
    1912: T492 = 1'h0;
    1913: T492 = 1'h0;
    1914: T492 = 1'h0;
    1915: T492 = 1'h0;
    1916: T492 = 1'h0;
    1917: T492 = 1'h0;
    1918: T492 = 1'h0;
    1919: T492 = 1'h0;
    1920: T492 = 1'h0;
    1921: T492 = 1'h0;
    1922: T492 = 1'h0;
    1923: T492 = 1'h0;
    1924: T492 = 1'h0;
    1925: T492 = 1'h0;
    1926: T492 = 1'h0;
    1927: T492 = 1'h0;
    1928: T492 = 1'h0;
    1929: T492 = 1'h0;
    1930: T492 = 1'h0;
    1931: T492 = 1'h0;
    1932: T492 = 1'h0;
    1933: T492 = 1'h0;
    1934: T492 = 1'h0;
    1935: T492 = 1'h0;
    1936: T492 = 1'h0;
    1937: T492 = 1'h0;
    1938: T492 = 1'h0;
    1939: T492 = 1'h0;
    1940: T492 = 1'h0;
    1941: T492 = 1'h0;
    1942: T492 = 1'h0;
    1943: T492 = 1'h0;
    1944: T492 = 1'h0;
    1945: T492 = 1'h0;
    1946: T492 = 1'h0;
    1947: T492 = 1'h0;
    1948: T492 = 1'h0;
    1949: T492 = 1'h0;
    1950: T492 = 1'h0;
    1951: T492 = 1'h0;
    1952: T492 = 1'h0;
    1953: T492 = 1'h0;
    1954: T492 = 1'h0;
    1955: T492 = 1'h0;
    1956: T492 = 1'h0;
    1957: T492 = 1'h0;
    1958: T492 = 1'h0;
    1959: T492 = 1'h0;
    1960: T492 = 1'h0;
    1961: T492 = 1'h0;
    1962: T492 = 1'h0;
    1963: T492 = 1'h0;
    1964: T492 = 1'h0;
    1965: T492 = 1'h0;
    1966: T492 = 1'h0;
    1967: T492 = 1'h0;
    1968: T492 = 1'h0;
    1969: T492 = 1'h0;
    1970: T492 = 1'h0;
    1971: T492 = 1'h0;
    1972: T492 = 1'h0;
    1973: T492 = 1'h0;
    1974: T492 = 1'h0;
    1975: T492 = 1'h0;
    1976: T492 = 1'h0;
    1977: T492 = 1'h0;
    1978: T492 = 1'h0;
    1979: T492 = 1'h0;
    1980: T492 = 1'h0;
    1981: T492 = 1'h0;
    1982: T492 = 1'h0;
    1983: T492 = 1'h0;
    1984: T492 = 1'h0;
    1985: T492 = 1'h0;
    1986: T492 = 1'h0;
    1987: T492 = 1'h0;
    1988: T492 = 1'h0;
    1989: T492 = 1'h0;
    1990: T492 = 1'h0;
    1991: T492 = 1'h0;
    1992: T492 = 1'h0;
    1993: T492 = 1'h0;
    1994: T492 = 1'h0;
    1995: T492 = 1'h0;
    1996: T492 = 1'h0;
    1997: T492 = 1'h0;
    1998: T492 = 1'h0;
    1999: T492 = 1'h0;
    2000: T492 = 1'h0;
    2001: T492 = 1'h0;
    2002: T492 = 1'h0;
    2003: T492 = 1'h0;
    2004: T492 = 1'h0;
    2005: T492 = 1'h0;
    2006: T492 = 1'h0;
    2007: T492 = 1'h0;
    2008: T492 = 1'h0;
    2009: T492 = 1'h0;
    2010: T492 = 1'h0;
    2011: T492 = 1'h0;
    2012: T492 = 1'h0;
    2013: T492 = 1'h0;
    2014: T492 = 1'h0;
    2015: T492 = 1'h0;
    2016: T492 = 1'h0;
    2017: T492 = 1'h0;
    2018: T492 = 1'h0;
    2019: T492 = 1'h0;
    2020: T492 = 1'h0;
    2021: T492 = 1'h0;
    2022: T492 = 1'h0;
    2023: T492 = 1'h0;
    2024: T492 = 1'h0;
    2025: T492 = 1'h0;
    2026: T492 = 1'h0;
    2027: T492 = 1'h0;
    2028: T492 = 1'h0;
    2029: T492 = 1'h0;
    2030: T492 = 1'h0;
    2031: T492 = 1'h0;
    2032: T492 = 1'h0;
    2033: T492 = 1'h0;
    2034: T492 = 1'h0;
    2035: T492 = 1'h0;
    2036: T492 = 1'h0;
    2037: T492 = 1'h0;
    2038: T492 = 1'h0;
    2039: T492 = 1'h0;
    2040: T492 = 1'h0;
    2041: T492 = 1'h0;
    2042: T492 = 1'h0;
    2043: T492 = 1'h0;
    2044: T492 = 1'h0;
    2045: T492 = 1'h0;
    2046: T492 = 1'h0;
    2047: T492 = 1'h0;
    2048: T492 = 1'h0;
    2049: T492 = 1'h0;
    2050: T492 = 1'h0;
    2051: T492 = 1'h0;
    2052: T492 = 1'h0;
    2053: T492 = 1'h0;
    2054: T492 = 1'h0;
    2055: T492 = 1'h0;
    2056: T492 = 1'h0;
    2057: T492 = 1'h0;
    2058: T492 = 1'h0;
    2059: T492 = 1'h0;
    2060: T492 = 1'h0;
    2061: T492 = 1'h0;
    2062: T492 = 1'h0;
    2063: T492 = 1'h0;
    2064: T492 = 1'h0;
    2065: T492 = 1'h0;
    2066: T492 = 1'h0;
    2067: T492 = 1'h0;
    2068: T492 = 1'h0;
    2069: T492 = 1'h0;
    2070: T492 = 1'h0;
    2071: T492 = 1'h0;
    2072: T492 = 1'h0;
    2073: T492 = 1'h0;
    2074: T492 = 1'h0;
    2075: T492 = 1'h0;
    2076: T492 = 1'h0;
    2077: T492 = 1'h0;
    2078: T492 = 1'h0;
    2079: T492 = 1'h0;
    2080: T492 = 1'h0;
    2081: T492 = 1'h0;
    2082: T492 = 1'h0;
    2083: T492 = 1'h0;
    2084: T492 = 1'h0;
    2085: T492 = 1'h0;
    2086: T492 = 1'h0;
    2087: T492 = 1'h0;
    2088: T492 = 1'h0;
    2089: T492 = 1'h0;
    2090: T492 = 1'h0;
    2091: T492 = 1'h0;
    2092: T492 = 1'h0;
    2093: T492 = 1'h0;
    2094: T492 = 1'h0;
    2095: T492 = 1'h0;
    2096: T492 = 1'h0;
    2097: T492 = 1'h0;
    2098: T492 = 1'h0;
    2099: T492 = 1'h0;
    2100: T492 = 1'h0;
    2101: T492 = 1'h0;
    2102: T492 = 1'h0;
    2103: T492 = 1'h0;
    2104: T492 = 1'h0;
    2105: T492 = 1'h0;
    2106: T492 = 1'h0;
    2107: T492 = 1'h0;
    2108: T492 = 1'h0;
    2109: T492 = 1'h0;
    2110: T492 = 1'h0;
    2111: T492 = 1'h0;
    2112: T492 = 1'h0;
    2113: T492 = 1'h0;
    2114: T492 = 1'h0;
    2115: T492 = 1'h0;
    2116: T492 = 1'h0;
    2117: T492 = 1'h0;
    2118: T492 = 1'h0;
    2119: T492 = 1'h0;
    2120: T492 = 1'h0;
    2121: T492 = 1'h0;
    2122: T492 = 1'h0;
    2123: T492 = 1'h0;
    2124: T492 = 1'h0;
    2125: T492 = 1'h0;
    2126: T492 = 1'h0;
    2127: T492 = 1'h0;
    2128: T492 = 1'h0;
    2129: T492 = 1'h0;
    2130: T492 = 1'h0;
    2131: T492 = 1'h0;
    2132: T492 = 1'h0;
    2133: T492 = 1'h0;
    2134: T492 = 1'h0;
    2135: T492 = 1'h0;
    2136: T492 = 1'h0;
    2137: T492 = 1'h0;
    2138: T492 = 1'h0;
    2139: T492 = 1'h0;
    2140: T492 = 1'h0;
    2141: T492 = 1'h0;
    2142: T492 = 1'h0;
    2143: T492 = 1'h0;
    2144: T492 = 1'h0;
    2145: T492 = 1'h0;
    2146: T492 = 1'h0;
    2147: T492 = 1'h0;
    2148: T492 = 1'h0;
    2149: T492 = 1'h0;
    2150: T492 = 1'h0;
    2151: T492 = 1'h0;
    2152: T492 = 1'h0;
    2153: T492 = 1'h0;
    2154: T492 = 1'h0;
    2155: T492 = 1'h0;
    2156: T492 = 1'h0;
    2157: T492 = 1'h0;
    2158: T492 = 1'h0;
    2159: T492 = 1'h0;
    2160: T492 = 1'h0;
    2161: T492 = 1'h0;
    2162: T492 = 1'h0;
    2163: T492 = 1'h0;
    2164: T492 = 1'h0;
    2165: T492 = 1'h0;
    2166: T492 = 1'h0;
    2167: T492 = 1'h0;
    2168: T492 = 1'h0;
    2169: T492 = 1'h0;
    2170: T492 = 1'h0;
    2171: T492 = 1'h0;
    2172: T492 = 1'h0;
    2173: T492 = 1'h0;
    2174: T492 = 1'h0;
    2175: T492 = 1'h0;
    2176: T492 = 1'h0;
    2177: T492 = 1'h0;
    2178: T492 = 1'h0;
    2179: T492 = 1'h0;
    2180: T492 = 1'h0;
    2181: T492 = 1'h0;
    2182: T492 = 1'h0;
    2183: T492 = 1'h0;
    2184: T492 = 1'h0;
    2185: T492 = 1'h0;
    2186: T492 = 1'h0;
    2187: T492 = 1'h0;
    2188: T492 = 1'h0;
    2189: T492 = 1'h0;
    2190: T492 = 1'h0;
    2191: T492 = 1'h0;
    2192: T492 = 1'h0;
    2193: T492 = 1'h0;
    2194: T492 = 1'h0;
    2195: T492 = 1'h0;
    2196: T492 = 1'h0;
    2197: T492 = 1'h0;
    2198: T492 = 1'h0;
    2199: T492 = 1'h0;
    2200: T492 = 1'h0;
    2201: T492 = 1'h0;
    2202: T492 = 1'h0;
    2203: T492 = 1'h0;
    2204: T492 = 1'h0;
    2205: T492 = 1'h0;
    2206: T492 = 1'h0;
    2207: T492 = 1'h0;
    2208: T492 = 1'h0;
    2209: T492 = 1'h0;
    2210: T492 = 1'h0;
    2211: T492 = 1'h0;
    2212: T492 = 1'h0;
    2213: T492 = 1'h0;
    2214: T492 = 1'h0;
    2215: T492 = 1'h0;
    2216: T492 = 1'h0;
    2217: T492 = 1'h0;
    2218: T492 = 1'h0;
    2219: T492 = 1'h0;
    2220: T492 = 1'h0;
    2221: T492 = 1'h0;
    2222: T492 = 1'h0;
    2223: T492 = 1'h0;
    2224: T492 = 1'h0;
    2225: T492 = 1'h0;
    2226: T492 = 1'h0;
    2227: T492 = 1'h0;
    2228: T492 = 1'h0;
    2229: T492 = 1'h0;
    2230: T492 = 1'h0;
    2231: T492 = 1'h0;
    2232: T492 = 1'h0;
    2233: T492 = 1'h0;
    2234: T492 = 1'h0;
    2235: T492 = 1'h0;
    2236: T492 = 1'h0;
    2237: T492 = 1'h0;
    2238: T492 = 1'h0;
    2239: T492 = 1'h0;
    2240: T492 = 1'h0;
    2241: T492 = 1'h0;
    2242: T492 = 1'h0;
    2243: T492 = 1'h0;
    2244: T492 = 1'h0;
    2245: T492 = 1'h0;
    2246: T492 = 1'h0;
    2247: T492 = 1'h0;
    2248: T492 = 1'h0;
    2249: T492 = 1'h0;
    2250: T492 = 1'h0;
    2251: T492 = 1'h0;
    2252: T492 = 1'h0;
    2253: T492 = 1'h0;
    2254: T492 = 1'h0;
    2255: T492 = 1'h0;
    2256: T492 = 1'h0;
    2257: T492 = 1'h0;
    2258: T492 = 1'h0;
    2259: T492 = 1'h0;
    2260: T492 = 1'h0;
    2261: T492 = 1'h0;
    2262: T492 = 1'h0;
    2263: T492 = 1'h0;
    2264: T492 = 1'h0;
    2265: T492 = 1'h0;
    2266: T492 = 1'h0;
    2267: T492 = 1'h0;
    2268: T492 = 1'h0;
    2269: T492 = 1'h0;
    2270: T492 = 1'h0;
    2271: T492 = 1'h0;
    2272: T492 = 1'h0;
    2273: T492 = 1'h0;
    2274: T492 = 1'h0;
    2275: T492 = 1'h0;
    2276: T492 = 1'h0;
    2277: T492 = 1'h0;
    2278: T492 = 1'h0;
    2279: T492 = 1'h0;
    2280: T492 = 1'h0;
    2281: T492 = 1'h0;
    2282: T492 = 1'h0;
    2283: T492 = 1'h0;
    2284: T492 = 1'h0;
    2285: T492 = 1'h0;
    2286: T492 = 1'h0;
    2287: T492 = 1'h0;
    2288: T492 = 1'h0;
    2289: T492 = 1'h0;
    2290: T492 = 1'h0;
    2291: T492 = 1'h0;
    2292: T492 = 1'h0;
    2293: T492 = 1'h0;
    2294: T492 = 1'h0;
    2295: T492 = 1'h0;
    2296: T492 = 1'h0;
    2297: T492 = 1'h0;
    2298: T492 = 1'h0;
    2299: T492 = 1'h0;
    2300: T492 = 1'h0;
    2301: T492 = 1'h0;
    2302: T492 = 1'h0;
    2303: T492 = 1'h0;
    2304: T492 = 1'h0;
    2305: T492 = 1'h0;
    2306: T492 = 1'h0;
    2307: T492 = 1'h0;
    2308: T492 = 1'h0;
    2309: T492 = 1'h0;
    2310: T492 = 1'h0;
    2311: T492 = 1'h0;
    2312: T492 = 1'h0;
    2313: T492 = 1'h0;
    2314: T492 = 1'h0;
    2315: T492 = 1'h0;
    2316: T492 = 1'h0;
    2317: T492 = 1'h0;
    2318: T492 = 1'h0;
    2319: T492 = 1'h0;
    2320: T492 = 1'h0;
    2321: T492 = 1'h0;
    2322: T492 = 1'h0;
    2323: T492 = 1'h0;
    2324: T492 = 1'h0;
    2325: T492 = 1'h0;
    2326: T492 = 1'h0;
    2327: T492 = 1'h0;
    2328: T492 = 1'h0;
    2329: T492 = 1'h0;
    2330: T492 = 1'h0;
    2331: T492 = 1'h0;
    2332: T492 = 1'h0;
    2333: T492 = 1'h0;
    2334: T492 = 1'h0;
    2335: T492 = 1'h0;
    2336: T492 = 1'h0;
    2337: T492 = 1'h0;
    2338: T492 = 1'h0;
    2339: T492 = 1'h0;
    2340: T492 = 1'h0;
    2341: T492 = 1'h0;
    2342: T492 = 1'h0;
    2343: T492 = 1'h0;
    2344: T492 = 1'h0;
    2345: T492 = 1'h0;
    2346: T492 = 1'h0;
    2347: T492 = 1'h0;
    2348: T492 = 1'h0;
    2349: T492 = 1'h0;
    2350: T492 = 1'h0;
    2351: T492 = 1'h0;
    2352: T492 = 1'h0;
    2353: T492 = 1'h0;
    2354: T492 = 1'h0;
    2355: T492 = 1'h0;
    2356: T492 = 1'h0;
    2357: T492 = 1'h0;
    2358: T492 = 1'h0;
    2359: T492 = 1'h0;
    2360: T492 = 1'h0;
    2361: T492 = 1'h0;
    2362: T492 = 1'h0;
    2363: T492 = 1'h0;
    2364: T492 = 1'h0;
    2365: T492 = 1'h0;
    2366: T492 = 1'h0;
    2367: T492 = 1'h0;
    2368: T492 = 1'h0;
    2369: T492 = 1'h0;
    2370: T492 = 1'h0;
    2371: T492 = 1'h0;
    2372: T492 = 1'h0;
    2373: T492 = 1'h0;
    2374: T492 = 1'h0;
    2375: T492 = 1'h0;
    2376: T492 = 1'h0;
    2377: T492 = 1'h0;
    2378: T492 = 1'h0;
    2379: T492 = 1'h0;
    2380: T492 = 1'h0;
    2381: T492 = 1'h0;
    2382: T492 = 1'h0;
    2383: T492 = 1'h0;
    2384: T492 = 1'h0;
    2385: T492 = 1'h0;
    2386: T492 = 1'h0;
    2387: T492 = 1'h0;
    2388: T492 = 1'h0;
    2389: T492 = 1'h0;
    2390: T492 = 1'h0;
    2391: T492 = 1'h0;
    2392: T492 = 1'h0;
    2393: T492 = 1'h0;
    2394: T492 = 1'h0;
    2395: T492 = 1'h0;
    2396: T492 = 1'h0;
    2397: T492 = 1'h0;
    2398: T492 = 1'h0;
    2399: T492 = 1'h0;
    2400: T492 = 1'h0;
    2401: T492 = 1'h0;
    2402: T492 = 1'h0;
    2403: T492 = 1'h0;
    2404: T492 = 1'h0;
    2405: T492 = 1'h0;
    2406: T492 = 1'h0;
    2407: T492 = 1'h0;
    2408: T492 = 1'h0;
    2409: T492 = 1'h0;
    2410: T492 = 1'h0;
    2411: T492 = 1'h0;
    2412: T492 = 1'h0;
    2413: T492 = 1'h0;
    2414: T492 = 1'h0;
    2415: T492 = 1'h0;
    2416: T492 = 1'h0;
    2417: T492 = 1'h0;
    2418: T492 = 1'h0;
    2419: T492 = 1'h0;
    2420: T492 = 1'h0;
    2421: T492 = 1'h0;
    2422: T492 = 1'h0;
    2423: T492 = 1'h0;
    2424: T492 = 1'h0;
    2425: T492 = 1'h0;
    2426: T492 = 1'h0;
    2427: T492 = 1'h0;
    2428: T492 = 1'h0;
    2429: T492 = 1'h0;
    2430: T492 = 1'h0;
    2431: T492 = 1'h0;
    2432: T492 = 1'h0;
    2433: T492 = 1'h0;
    2434: T492 = 1'h0;
    2435: T492 = 1'h0;
    2436: T492 = 1'h0;
    2437: T492 = 1'h0;
    2438: T492 = 1'h0;
    2439: T492 = 1'h0;
    2440: T492 = 1'h0;
    2441: T492 = 1'h0;
    2442: T492 = 1'h0;
    2443: T492 = 1'h0;
    2444: T492 = 1'h0;
    2445: T492 = 1'h0;
    2446: T492 = 1'h0;
    2447: T492 = 1'h0;
    2448: T492 = 1'h0;
    2449: T492 = 1'h0;
    2450: T492 = 1'h0;
    2451: T492 = 1'h0;
    2452: T492 = 1'h0;
    2453: T492 = 1'h0;
    2454: T492 = 1'h0;
    2455: T492 = 1'h0;
    2456: T492 = 1'h0;
    2457: T492 = 1'h0;
    2458: T492 = 1'h0;
    2459: T492 = 1'h0;
    2460: T492 = 1'h0;
    2461: T492 = 1'h0;
    2462: T492 = 1'h0;
    2463: T492 = 1'h0;
    2464: T492 = 1'h0;
    2465: T492 = 1'h0;
    2466: T492 = 1'h0;
    2467: T492 = 1'h0;
    2468: T492 = 1'h0;
    2469: T492 = 1'h0;
    2470: T492 = 1'h0;
    2471: T492 = 1'h0;
    2472: T492 = 1'h0;
    2473: T492 = 1'h0;
    2474: T492 = 1'h0;
    2475: T492 = 1'h0;
    2476: T492 = 1'h0;
    2477: T492 = 1'h0;
    2478: T492 = 1'h0;
    2479: T492 = 1'h0;
    2480: T492 = 1'h0;
    2481: T492 = 1'h0;
    2482: T492 = 1'h0;
    2483: T492 = 1'h0;
    2484: T492 = 1'h0;
    2485: T492 = 1'h0;
    2486: T492 = 1'h0;
    2487: T492 = 1'h0;
    2488: T492 = 1'h0;
    2489: T492 = 1'h0;
    2490: T492 = 1'h0;
    2491: T492 = 1'h0;
    2492: T492 = 1'h0;
    2493: T492 = 1'h0;
    2494: T492 = 1'h0;
    2495: T492 = 1'h0;
    2496: T492 = 1'h0;
    2497: T492 = 1'h0;
    2498: T492 = 1'h0;
    2499: T492 = 1'h0;
    2500: T492 = 1'h0;
    2501: T492 = 1'h0;
    2502: T492 = 1'h0;
    2503: T492 = 1'h0;
    2504: T492 = 1'h0;
    2505: T492 = 1'h0;
    2506: T492 = 1'h0;
    2507: T492 = 1'h0;
    2508: T492 = 1'h0;
    2509: T492 = 1'h0;
    2510: T492 = 1'h0;
    2511: T492 = 1'h0;
    2512: T492 = 1'h0;
    2513: T492 = 1'h0;
    2514: T492 = 1'h0;
    2515: T492 = 1'h0;
    2516: T492 = 1'h0;
    2517: T492 = 1'h0;
    2518: T492 = 1'h0;
    2519: T492 = 1'h0;
    2520: T492 = 1'h0;
    2521: T492 = 1'h0;
    2522: T492 = 1'h0;
    2523: T492 = 1'h0;
    2524: T492 = 1'h0;
    2525: T492 = 1'h0;
    2526: T492 = 1'h0;
    2527: T492 = 1'h0;
    2528: T492 = 1'h0;
    2529: T492 = 1'h0;
    2530: T492 = 1'h0;
    2531: T492 = 1'h0;
    2532: T492 = 1'h0;
    2533: T492 = 1'h0;
    2534: T492 = 1'h0;
    2535: T492 = 1'h0;
    2536: T492 = 1'h0;
    2537: T492 = 1'h0;
    2538: T492 = 1'h0;
    2539: T492 = 1'h0;
    2540: T492 = 1'h0;
    2541: T492 = 1'h0;
    2542: T492 = 1'h0;
    2543: T492 = 1'h0;
    2544: T492 = 1'h0;
    2545: T492 = 1'h0;
    2546: T492 = 1'h0;
    2547: T492 = 1'h0;
    2548: T492 = 1'h0;
    2549: T492 = 1'h0;
    2550: T492 = 1'h0;
    2551: T492 = 1'h0;
    2552: T492 = 1'h0;
    2553: T492 = 1'h0;
    2554: T492 = 1'h0;
    2555: T492 = 1'h0;
    2556: T492 = 1'h0;
    2557: T492 = 1'h0;
    2558: T492 = 1'h0;
    2559: T492 = 1'h0;
    2560: T492 = 1'h0;
    2561: T492 = 1'h0;
    2562: T492 = 1'h0;
    2563: T492 = 1'h0;
    2564: T492 = 1'h0;
    2565: T492 = 1'h0;
    2566: T492 = 1'h0;
    2567: T492 = 1'h0;
    2568: T492 = 1'h0;
    2569: T492 = 1'h0;
    2570: T492 = 1'h0;
    2571: T492 = 1'h0;
    2572: T492 = 1'h0;
    2573: T492 = 1'h0;
    2574: T492 = 1'h0;
    2575: T492 = 1'h0;
    2576: T492 = 1'h0;
    2577: T492 = 1'h0;
    2578: T492 = 1'h0;
    2579: T492 = 1'h0;
    2580: T492 = 1'h0;
    2581: T492 = 1'h0;
    2582: T492 = 1'h0;
    2583: T492 = 1'h0;
    2584: T492 = 1'h0;
    2585: T492 = 1'h0;
    2586: T492 = 1'h0;
    2587: T492 = 1'h0;
    2588: T492 = 1'h0;
    2589: T492 = 1'h0;
    2590: T492 = 1'h0;
    2591: T492 = 1'h0;
    2592: T492 = 1'h0;
    2593: T492 = 1'h0;
    2594: T492 = 1'h0;
    2595: T492 = 1'h0;
    2596: T492 = 1'h0;
    2597: T492 = 1'h0;
    2598: T492 = 1'h0;
    2599: T492 = 1'h0;
    2600: T492 = 1'h0;
    2601: T492 = 1'h0;
    2602: T492 = 1'h0;
    2603: T492 = 1'h0;
    2604: T492 = 1'h0;
    2605: T492 = 1'h0;
    2606: T492 = 1'h0;
    2607: T492 = 1'h0;
    2608: T492 = 1'h0;
    2609: T492 = 1'h0;
    2610: T492 = 1'h0;
    2611: T492 = 1'h0;
    2612: T492 = 1'h0;
    2613: T492 = 1'h0;
    2614: T492 = 1'h0;
    2615: T492 = 1'h0;
    2616: T492 = 1'h0;
    2617: T492 = 1'h0;
    2618: T492 = 1'h0;
    2619: T492 = 1'h0;
    2620: T492 = 1'h0;
    2621: T492 = 1'h0;
    2622: T492 = 1'h0;
    2623: T492 = 1'h0;
    2624: T492 = 1'h0;
    2625: T492 = 1'h0;
    2626: T492 = 1'h0;
    2627: T492 = 1'h0;
    2628: T492 = 1'h0;
    2629: T492 = 1'h0;
    2630: T492 = 1'h0;
    2631: T492 = 1'h0;
    2632: T492 = 1'h0;
    2633: T492 = 1'h0;
    2634: T492 = 1'h0;
    2635: T492 = 1'h0;
    2636: T492 = 1'h0;
    2637: T492 = 1'h0;
    2638: T492 = 1'h0;
    2639: T492 = 1'h0;
    2640: T492 = 1'h0;
    2641: T492 = 1'h0;
    2642: T492 = 1'h0;
    2643: T492 = 1'h0;
    2644: T492 = 1'h0;
    2645: T492 = 1'h0;
    2646: T492 = 1'h0;
    2647: T492 = 1'h0;
    2648: T492 = 1'h0;
    2649: T492 = 1'h0;
    2650: T492 = 1'h0;
    2651: T492 = 1'h0;
    2652: T492 = 1'h0;
    2653: T492 = 1'h0;
    2654: T492 = 1'h0;
    2655: T492 = 1'h0;
    2656: T492 = 1'h0;
    2657: T492 = 1'h0;
    2658: T492 = 1'h0;
    2659: T492 = 1'h0;
    2660: T492 = 1'h0;
    2661: T492 = 1'h0;
    2662: T492 = 1'h0;
    2663: T492 = 1'h0;
    2664: T492 = 1'h0;
    2665: T492 = 1'h0;
    2666: T492 = 1'h0;
    2667: T492 = 1'h0;
    2668: T492 = 1'h0;
    2669: T492 = 1'h0;
    2670: T492 = 1'h0;
    2671: T492 = 1'h0;
    2672: T492 = 1'h0;
    2673: T492 = 1'h0;
    2674: T492 = 1'h0;
    2675: T492 = 1'h0;
    2676: T492 = 1'h0;
    2677: T492 = 1'h0;
    2678: T492 = 1'h0;
    2679: T492 = 1'h0;
    2680: T492 = 1'h0;
    2681: T492 = 1'h0;
    2682: T492 = 1'h0;
    2683: T492 = 1'h0;
    2684: T492 = 1'h0;
    2685: T492 = 1'h0;
    2686: T492 = 1'h0;
    2687: T492 = 1'h0;
    2688: T492 = 1'h0;
    2689: T492 = 1'h0;
    2690: T492 = 1'h0;
    2691: T492 = 1'h0;
    2692: T492 = 1'h0;
    2693: T492 = 1'h0;
    2694: T492 = 1'h0;
    2695: T492 = 1'h0;
    2696: T492 = 1'h0;
    2697: T492 = 1'h0;
    2698: T492 = 1'h0;
    2699: T492 = 1'h0;
    2700: T492 = 1'h0;
    2701: T492 = 1'h0;
    2702: T492 = 1'h0;
    2703: T492 = 1'h0;
    2704: T492 = 1'h0;
    2705: T492 = 1'h0;
    2706: T492 = 1'h0;
    2707: T492 = 1'h0;
    2708: T492 = 1'h0;
    2709: T492 = 1'h0;
    2710: T492 = 1'h0;
    2711: T492 = 1'h0;
    2712: T492 = 1'h0;
    2713: T492 = 1'h0;
    2714: T492 = 1'h0;
    2715: T492 = 1'h0;
    2716: T492 = 1'h0;
    2717: T492 = 1'h0;
    2718: T492 = 1'h0;
    2719: T492 = 1'h0;
    2720: T492 = 1'h0;
    2721: T492 = 1'h0;
    2722: T492 = 1'h0;
    2723: T492 = 1'h0;
    2724: T492 = 1'h0;
    2725: T492 = 1'h0;
    2726: T492 = 1'h0;
    2727: T492 = 1'h0;
    2728: T492 = 1'h0;
    2729: T492 = 1'h0;
    2730: T492 = 1'h0;
    2731: T492 = 1'h0;
    2732: T492 = 1'h0;
    2733: T492 = 1'h0;
    2734: T492 = 1'h0;
    2735: T492 = 1'h0;
    2736: T492 = 1'h0;
    2737: T492 = 1'h0;
    2738: T492 = 1'h0;
    2739: T492 = 1'h0;
    2740: T492 = 1'h0;
    2741: T492 = 1'h0;
    2742: T492 = 1'h0;
    2743: T492 = 1'h0;
    2744: T492 = 1'h0;
    2745: T492 = 1'h0;
    2746: T492 = 1'h0;
    2747: T492 = 1'h0;
    2748: T492 = 1'h0;
    2749: T492 = 1'h0;
    2750: T492 = 1'h0;
    2751: T492 = 1'h0;
    2752: T492 = 1'h0;
    2753: T492 = 1'h0;
    2754: T492 = 1'h0;
    2755: T492 = 1'h0;
    2756: T492 = 1'h0;
    2757: T492 = 1'h0;
    2758: T492 = 1'h0;
    2759: T492 = 1'h0;
    2760: T492 = 1'h0;
    2761: T492 = 1'h0;
    2762: T492 = 1'h0;
    2763: T492 = 1'h0;
    2764: T492 = 1'h0;
    2765: T492 = 1'h0;
    2766: T492 = 1'h0;
    2767: T492 = 1'h0;
    2768: T492 = 1'h0;
    2769: T492 = 1'h0;
    2770: T492 = 1'h0;
    2771: T492 = 1'h0;
    2772: T492 = 1'h0;
    2773: T492 = 1'h0;
    2774: T492 = 1'h0;
    2775: T492 = 1'h0;
    2776: T492 = 1'h0;
    2777: T492 = 1'h0;
    2778: T492 = 1'h0;
    2779: T492 = 1'h0;
    2780: T492 = 1'h0;
    2781: T492 = 1'h0;
    2782: T492 = 1'h0;
    2783: T492 = 1'h0;
    2784: T492 = 1'h0;
    2785: T492 = 1'h0;
    2786: T492 = 1'h0;
    2787: T492 = 1'h0;
    2788: T492 = 1'h0;
    2789: T492 = 1'h0;
    2790: T492 = 1'h0;
    2791: T492 = 1'h0;
    2792: T492 = 1'h0;
    2793: T492 = 1'h0;
    2794: T492 = 1'h0;
    2795: T492 = 1'h0;
    2796: T492 = 1'h0;
    2797: T492 = 1'h0;
    2798: T492 = 1'h0;
    2799: T492 = 1'h0;
    2800: T492 = 1'h0;
    2801: T492 = 1'h0;
    2802: T492 = 1'h0;
    2803: T492 = 1'h0;
    2804: T492 = 1'h0;
    2805: T492 = 1'h0;
    2806: T492 = 1'h0;
    2807: T492 = 1'h0;
    2808: T492 = 1'h0;
    2809: T492 = 1'h0;
    2810: T492 = 1'h0;
    2811: T492 = 1'h0;
    2812: T492 = 1'h0;
    2813: T492 = 1'h0;
    2814: T492 = 1'h0;
    2815: T492 = 1'h0;
    2816: T492 = 1'h0;
    2817: T492 = 1'h0;
    2818: T492 = 1'h0;
    2819: T492 = 1'h0;
    2820: T492 = 1'h0;
    2821: T492 = 1'h0;
    2822: T492 = 1'h0;
    2823: T492 = 1'h0;
    2824: T492 = 1'h0;
    2825: T492 = 1'h0;
    2826: T492 = 1'h0;
    2827: T492 = 1'h0;
    2828: T492 = 1'h0;
    2829: T492 = 1'h0;
    2830: T492 = 1'h0;
    2831: T492 = 1'h0;
    2832: T492 = 1'h0;
    2833: T492 = 1'h0;
    2834: T492 = 1'h0;
    2835: T492 = 1'h0;
    2836: T492 = 1'h0;
    2837: T492 = 1'h0;
    2838: T492 = 1'h0;
    2839: T492 = 1'h0;
    2840: T492 = 1'h0;
    2841: T492 = 1'h0;
    2842: T492 = 1'h0;
    2843: T492 = 1'h0;
    2844: T492 = 1'h0;
    2845: T492 = 1'h0;
    2846: T492 = 1'h0;
    2847: T492 = 1'h0;
    2848: T492 = 1'h0;
    2849: T492 = 1'h0;
    2850: T492 = 1'h0;
    2851: T492 = 1'h0;
    2852: T492 = 1'h0;
    2853: T492 = 1'h0;
    2854: T492 = 1'h0;
    2855: T492 = 1'h0;
    2856: T492 = 1'h0;
    2857: T492 = 1'h0;
    2858: T492 = 1'h0;
    2859: T492 = 1'h0;
    2860: T492 = 1'h0;
    2861: T492 = 1'h0;
    2862: T492 = 1'h0;
    2863: T492 = 1'h0;
    2864: T492 = 1'h0;
    2865: T492 = 1'h0;
    2866: T492 = 1'h0;
    2867: T492 = 1'h0;
    2868: T492 = 1'h0;
    2869: T492 = 1'h0;
    2870: T492 = 1'h0;
    2871: T492 = 1'h0;
    2872: T492 = 1'h0;
    2873: T492 = 1'h0;
    2874: T492 = 1'h0;
    2875: T492 = 1'h0;
    2876: T492 = 1'h0;
    2877: T492 = 1'h0;
    2878: T492 = 1'h0;
    2879: T492 = 1'h0;
    2880: T492 = 1'h0;
    2881: T492 = 1'h0;
    2882: T492 = 1'h0;
    2883: T492 = 1'h0;
    2884: T492 = 1'h0;
    2885: T492 = 1'h0;
    2886: T492 = 1'h0;
    2887: T492 = 1'h0;
    2888: T492 = 1'h0;
    2889: T492 = 1'h0;
    2890: T492 = 1'h0;
    2891: T492 = 1'h0;
    2892: T492 = 1'h0;
    2893: T492 = 1'h0;
    2894: T492 = 1'h0;
    2895: T492 = 1'h0;
    2896: T492 = 1'h0;
    2897: T492 = 1'h0;
    2898: T492 = 1'h0;
    2899: T492 = 1'h0;
    2900: T492 = 1'h0;
    2901: T492 = 1'h0;
    2902: T492 = 1'h0;
    2903: T492 = 1'h0;
    2904: T492 = 1'h0;
    2905: T492 = 1'h0;
    2906: T492 = 1'h0;
    2907: T492 = 1'h0;
    2908: T492 = 1'h0;
    2909: T492 = 1'h0;
    2910: T492 = 1'h0;
    2911: T492 = 1'h0;
    2912: T492 = 1'h0;
    2913: T492 = 1'h0;
    2914: T492 = 1'h0;
    2915: T492 = 1'h0;
    2916: T492 = 1'h0;
    2917: T492 = 1'h0;
    2918: T492 = 1'h0;
    2919: T492 = 1'h0;
    2920: T492 = 1'h0;
    2921: T492 = 1'h0;
    2922: T492 = 1'h0;
    2923: T492 = 1'h0;
    2924: T492 = 1'h0;
    2925: T492 = 1'h0;
    2926: T492 = 1'h0;
    2927: T492 = 1'h0;
    2928: T492 = 1'h0;
    2929: T492 = 1'h0;
    2930: T492 = 1'h0;
    2931: T492 = 1'h0;
    2932: T492 = 1'h0;
    2933: T492 = 1'h0;
    2934: T492 = 1'h0;
    2935: T492 = 1'h0;
    2936: T492 = 1'h0;
    2937: T492 = 1'h0;
    2938: T492 = 1'h0;
    2939: T492 = 1'h0;
    2940: T492 = 1'h0;
    2941: T492 = 1'h0;
    2942: T492 = 1'h0;
    2943: T492 = 1'h0;
    2944: T492 = 1'h0;
    2945: T492 = 1'h0;
    2946: T492 = 1'h0;
    2947: T492 = 1'h0;
    2948: T492 = 1'h0;
    2949: T492 = 1'h0;
    2950: T492 = 1'h0;
    2951: T492 = 1'h0;
    2952: T492 = 1'h0;
    2953: T492 = 1'h0;
    2954: T492 = 1'h0;
    2955: T492 = 1'h0;
    2956: T492 = 1'h0;
    2957: T492 = 1'h0;
    2958: T492 = 1'h0;
    2959: T492 = 1'h0;
    2960: T492 = 1'h0;
    2961: T492 = 1'h0;
    2962: T492 = 1'h0;
    2963: T492 = 1'h0;
    2964: T492 = 1'h0;
    2965: T492 = 1'h0;
    2966: T492 = 1'h0;
    2967: T492 = 1'h0;
    2968: T492 = 1'h0;
    2969: T492 = 1'h0;
    2970: T492 = 1'h0;
    2971: T492 = 1'h0;
    2972: T492 = 1'h0;
    2973: T492 = 1'h0;
    2974: T492 = 1'h0;
    2975: T492 = 1'h0;
    2976: T492 = 1'h0;
    2977: T492 = 1'h0;
    2978: T492 = 1'h0;
    2979: T492 = 1'h0;
    2980: T492 = 1'h0;
    2981: T492 = 1'h0;
    2982: T492 = 1'h0;
    2983: T492 = 1'h0;
    2984: T492 = 1'h0;
    2985: T492 = 1'h0;
    2986: T492 = 1'h0;
    2987: T492 = 1'h0;
    2988: T492 = 1'h0;
    2989: T492 = 1'h0;
    2990: T492 = 1'h0;
    2991: T492 = 1'h0;
    2992: T492 = 1'h0;
    2993: T492 = 1'h0;
    2994: T492 = 1'h0;
    2995: T492 = 1'h0;
    2996: T492 = 1'h0;
    2997: T492 = 1'h0;
    2998: T492 = 1'h0;
    2999: T492 = 1'h0;
    3000: T492 = 1'h0;
    3001: T492 = 1'h0;
    3002: T492 = 1'h0;
    3003: T492 = 1'h0;
    3004: T492 = 1'h0;
    3005: T492 = 1'h0;
    3006: T492 = 1'h0;
    3007: T492 = 1'h0;
    3008: T492 = 1'h0;
    3009: T492 = 1'h0;
    3010: T492 = 1'h0;
    3011: T492 = 1'h0;
    3012: T492 = 1'h0;
    3013: T492 = 1'h0;
    3014: T492 = 1'h0;
    3015: T492 = 1'h0;
    3016: T492 = 1'h0;
    3017: T492 = 1'h0;
    3018: T492 = 1'h0;
    3019: T492 = 1'h0;
    3020: T492 = 1'h0;
    3021: T492 = 1'h0;
    3022: T492 = 1'h0;
    3023: T492 = 1'h0;
    3024: T492 = 1'h0;
    3025: T492 = 1'h0;
    3026: T492 = 1'h0;
    3027: T492 = 1'h0;
    3028: T492 = 1'h0;
    3029: T492 = 1'h0;
    3030: T492 = 1'h0;
    3031: T492 = 1'h0;
    3032: T492 = 1'h0;
    3033: T492 = 1'h0;
    3034: T492 = 1'h0;
    3035: T492 = 1'h0;
    3036: T492 = 1'h0;
    3037: T492 = 1'h0;
    3038: T492 = 1'h0;
    3039: T492 = 1'h0;
    3040: T492 = 1'h0;
    3041: T492 = 1'h0;
    3042: T492 = 1'h0;
    3043: T492 = 1'h0;
    3044: T492 = 1'h0;
    3045: T492 = 1'h0;
    3046: T492 = 1'h0;
    3047: T492 = 1'h0;
    3048: T492 = 1'h0;
    3049: T492 = 1'h0;
    3050: T492 = 1'h0;
    3051: T492 = 1'h0;
    3052: T492 = 1'h0;
    3053: T492 = 1'h0;
    3054: T492 = 1'h0;
    3055: T492 = 1'h0;
    3056: T492 = 1'h0;
    3057: T492 = 1'h0;
    3058: T492 = 1'h0;
    3059: T492 = 1'h0;
    3060: T492 = 1'h0;
    3061: T492 = 1'h0;
    3062: T492 = 1'h0;
    3063: T492 = 1'h0;
    3064: T492 = 1'h0;
    3065: T492 = 1'h0;
    3066: T492 = 1'h0;
    3067: T492 = 1'h0;
    3068: T492 = 1'h0;
    3069: T492 = 1'h0;
    3070: T492 = 1'h0;
    3071: T492 = 1'h0;
    3072: T492 = 1'h1;
    3073: T492 = 1'h1;
    3074: T492 = 1'h1;
    3075: T492 = 1'h0;
    3076: T492 = 1'h0;
    3077: T492 = 1'h0;
    3078: T492 = 1'h0;
    3079: T492 = 1'h0;
    3080: T492 = 1'h0;
    3081: T492 = 1'h0;
    3082: T492 = 1'h0;
    3083: T492 = 1'h0;
    3084: T492 = 1'h0;
    3085: T492 = 1'h0;
    3086: T492 = 1'h0;
    3087: T492 = 1'h0;
    3088: T492 = 1'h0;
    3089: T492 = 1'h0;
    3090: T492 = 1'h0;
    3091: T492 = 1'h0;
    3092: T492 = 1'h0;
    3093: T492 = 1'h0;
    3094: T492 = 1'h0;
    3095: T492 = 1'h0;
    3096: T492 = 1'h0;
    3097: T492 = 1'h0;
    3098: T492 = 1'h0;
    3099: T492 = 1'h0;
    3100: T492 = 1'h0;
    3101: T492 = 1'h0;
    3102: T492 = 1'h0;
    3103: T492 = 1'h0;
    3104: T492 = 1'h0;
    3105: T492 = 1'h0;
    3106: T492 = 1'h0;
    3107: T492 = 1'h0;
    3108: T492 = 1'h0;
    3109: T492 = 1'h0;
    3110: T492 = 1'h0;
    3111: T492 = 1'h0;
    3112: T492 = 1'h0;
    3113: T492 = 1'h0;
    3114: T492 = 1'h0;
    3115: T492 = 1'h0;
    3116: T492 = 1'h0;
    3117: T492 = 1'h0;
    3118: T492 = 1'h0;
    3119: T492 = 1'h0;
    3120: T492 = 1'h0;
    3121: T492 = 1'h0;
    3122: T492 = 1'h0;
    3123: T492 = 1'h0;
    3124: T492 = 1'h0;
    3125: T492 = 1'h0;
    3126: T492 = 1'h0;
    3127: T492 = 1'h0;
    3128: T492 = 1'h0;
    3129: T492 = 1'h0;
    3130: T492 = 1'h0;
    3131: T492 = 1'h0;
    3132: T492 = 1'h0;
    3133: T492 = 1'h0;
    3134: T492 = 1'h0;
    3135: T492 = 1'h0;
    3136: T492 = 1'h0;
    3137: T492 = 1'h0;
    3138: T492 = 1'h0;
    3139: T492 = 1'h0;
    3140: T492 = 1'h0;
    3141: T492 = 1'h0;
    3142: T492 = 1'h0;
    3143: T492 = 1'h0;
    3144: T492 = 1'h0;
    3145: T492 = 1'h0;
    3146: T492 = 1'h0;
    3147: T492 = 1'h0;
    3148: T492 = 1'h0;
    3149: T492 = 1'h0;
    3150: T492 = 1'h0;
    3151: T492 = 1'h0;
    3152: T492 = 1'h0;
    3153: T492 = 1'h0;
    3154: T492 = 1'h0;
    3155: T492 = 1'h0;
    3156: T492 = 1'h0;
    3157: T492 = 1'h0;
    3158: T492 = 1'h0;
    3159: T492 = 1'h0;
    3160: T492 = 1'h0;
    3161: T492 = 1'h0;
    3162: T492 = 1'h0;
    3163: T492 = 1'h0;
    3164: T492 = 1'h0;
    3165: T492 = 1'h0;
    3166: T492 = 1'h0;
    3167: T492 = 1'h0;
    3168: T492 = 1'h0;
    3169: T492 = 1'h0;
    3170: T492 = 1'h0;
    3171: T492 = 1'h0;
    3172: T492 = 1'h0;
    3173: T492 = 1'h0;
    3174: T492 = 1'h0;
    3175: T492 = 1'h0;
    3176: T492 = 1'h0;
    3177: T492 = 1'h0;
    3178: T492 = 1'h0;
    3179: T492 = 1'h0;
    3180: T492 = 1'h0;
    3181: T492 = 1'h0;
    3182: T492 = 1'h0;
    3183: T492 = 1'h0;
    3184: T492 = 1'h0;
    3185: T492 = 1'h0;
    3186: T492 = 1'h0;
    3187: T492 = 1'h0;
    3188: T492 = 1'h0;
    3189: T492 = 1'h0;
    3190: T492 = 1'h0;
    3191: T492 = 1'h0;
    3192: T492 = 1'h0;
    3193: T492 = 1'h0;
    3194: T492 = 1'h0;
    3195: T492 = 1'h0;
    3196: T492 = 1'h0;
    3197: T492 = 1'h0;
    3198: T492 = 1'h0;
    3199: T492 = 1'h0;
    3200: T492 = 1'h0;
    3201: T492 = 1'h0;
    3202: T492 = 1'h0;
    3203: T492 = 1'h0;
    3204: T492 = 1'h0;
    3205: T492 = 1'h0;
    3206: T492 = 1'h0;
    3207: T492 = 1'h0;
    3208: T492 = 1'h0;
    3209: T492 = 1'h0;
    3210: T492 = 1'h0;
    3211: T492 = 1'h0;
    3212: T492 = 1'h0;
    3213: T492 = 1'h0;
    3214: T492 = 1'h0;
    3215: T492 = 1'h0;
    3216: T492 = 1'h0;
    3217: T492 = 1'h0;
    3218: T492 = 1'h0;
    3219: T492 = 1'h0;
    3220: T492 = 1'h0;
    3221: T492 = 1'h0;
    3222: T492 = 1'h0;
    3223: T492 = 1'h0;
    3224: T492 = 1'h0;
    3225: T492 = 1'h0;
    3226: T492 = 1'h0;
    3227: T492 = 1'h0;
    3228: T492 = 1'h0;
    3229: T492 = 1'h0;
    3230: T492 = 1'h0;
    3231: T492 = 1'h0;
    3232: T492 = 1'h0;
    3233: T492 = 1'h0;
    3234: T492 = 1'h0;
    3235: T492 = 1'h0;
    3236: T492 = 1'h0;
    3237: T492 = 1'h0;
    3238: T492 = 1'h0;
    3239: T492 = 1'h0;
    3240: T492 = 1'h0;
    3241: T492 = 1'h0;
    3242: T492 = 1'h0;
    3243: T492 = 1'h0;
    3244: T492 = 1'h0;
    3245: T492 = 1'h0;
    3246: T492 = 1'h0;
    3247: T492 = 1'h0;
    3248: T492 = 1'h0;
    3249: T492 = 1'h0;
    3250: T492 = 1'h0;
    3251: T492 = 1'h0;
    3252: T492 = 1'h0;
    3253: T492 = 1'h0;
    3254: T492 = 1'h0;
    3255: T492 = 1'h0;
    3256: T492 = 1'h0;
    3257: T492 = 1'h0;
    3258: T492 = 1'h0;
    3259: T492 = 1'h0;
    3260: T492 = 1'h0;
    3261: T492 = 1'h0;
    3262: T492 = 1'h0;
    3263: T492 = 1'h0;
    3264: T492 = 1'h1;
    3265: T492 = 1'h1;
    3266: T492 = 1'h1;
    3267: T492 = 1'h1;
    3268: T492 = 1'h1;
    3269: T492 = 1'h1;
    3270: T492 = 1'h1;
    3271: T492 = 1'h1;
    3272: T492 = 1'h1;
    3273: T492 = 1'h1;
    3274: T492 = 1'h1;
    3275: T492 = 1'h1;
    3276: T492 = 1'h1;
    3277: T492 = 1'h1;
    3278: T492 = 1'h1;
    3279: T492 = 1'h1;
    3280: T492 = 1'h0;
    3281: T492 = 1'h0;
    3282: T492 = 1'h0;
    3283: T492 = 1'h0;
    3284: T492 = 1'h0;
    3285: T492 = 1'h0;
    3286: T492 = 1'h0;
    3287: T492 = 1'h0;
    3288: T492 = 1'h0;
    3289: T492 = 1'h0;
    3290: T492 = 1'h0;
    3291: T492 = 1'h0;
    3292: T492 = 1'h0;
    3293: T492 = 1'h0;
    3294: T492 = 1'h0;
    3295: T492 = 1'h0;
    3296: T492 = 1'h0;
    3297: T492 = 1'h0;
    3298: T492 = 1'h0;
    3299: T492 = 1'h0;
    3300: T492 = 1'h0;
    3301: T492 = 1'h0;
    3302: T492 = 1'h0;
    3303: T492 = 1'h0;
    3304: T492 = 1'h0;
    3305: T492 = 1'h0;
    3306: T492 = 1'h0;
    3307: T492 = 1'h0;
    3308: T492 = 1'h0;
    3309: T492 = 1'h0;
    3310: T492 = 1'h0;
    3311: T492 = 1'h0;
    3312: T492 = 1'h0;
    3313: T492 = 1'h0;
    3314: T492 = 1'h0;
    3315: T492 = 1'h0;
    3316: T492 = 1'h0;
    3317: T492 = 1'h0;
    3318: T492 = 1'h0;
    3319: T492 = 1'h0;
    3320: T492 = 1'h0;
    3321: T492 = 1'h0;
    3322: T492 = 1'h0;
    3323: T492 = 1'h0;
    3324: T492 = 1'h0;
    3325: T492 = 1'h0;
    3326: T492 = 1'h0;
    3327: T492 = 1'h0;
    3328: T492 = 1'h0;
    3329: T492 = 1'h0;
    3330: T492 = 1'h0;
    3331: T492 = 1'h0;
    3332: T492 = 1'h0;
    3333: T492 = 1'h0;
    3334: T492 = 1'h0;
    3335: T492 = 1'h0;
    3336: T492 = 1'h0;
    3337: T492 = 1'h0;
    3338: T492 = 1'h0;
    3339: T492 = 1'h0;
    3340: T492 = 1'h0;
    3341: T492 = 1'h0;
    3342: T492 = 1'h0;
    3343: T492 = 1'h0;
    3344: T492 = 1'h0;
    3345: T492 = 1'h0;
    3346: T492 = 1'h0;
    3347: T492 = 1'h0;
    3348: T492 = 1'h0;
    3349: T492 = 1'h0;
    3350: T492 = 1'h0;
    3351: T492 = 1'h0;
    3352: T492 = 1'h0;
    3353: T492 = 1'h0;
    3354: T492 = 1'h0;
    3355: T492 = 1'h0;
    3356: T492 = 1'h0;
    3357: T492 = 1'h0;
    3358: T492 = 1'h0;
    3359: T492 = 1'h0;
    3360: T492 = 1'h0;
    3361: T492 = 1'h0;
    3362: T492 = 1'h0;
    3363: T492 = 1'h0;
    3364: T492 = 1'h0;
    3365: T492 = 1'h0;
    3366: T492 = 1'h0;
    3367: T492 = 1'h0;
    3368: T492 = 1'h0;
    3369: T492 = 1'h0;
    3370: T492 = 1'h0;
    3371: T492 = 1'h0;
    3372: T492 = 1'h0;
    3373: T492 = 1'h0;
    3374: T492 = 1'h0;
    3375: T492 = 1'h0;
    3376: T492 = 1'h0;
    3377: T492 = 1'h0;
    3378: T492 = 1'h0;
    3379: T492 = 1'h0;
    3380: T492 = 1'h0;
    3381: T492 = 1'h0;
    3382: T492 = 1'h0;
    3383: T492 = 1'h0;
    3384: T492 = 1'h0;
    3385: T492 = 1'h0;
    3386: T492 = 1'h0;
    3387: T492 = 1'h0;
    3388: T492 = 1'h0;
    3389: T492 = 1'h0;
    3390: T492 = 1'h0;
    3391: T492 = 1'h0;
    3392: T492 = 1'h0;
    3393: T492 = 1'h0;
    3394: T492 = 1'h0;
    3395: T492 = 1'h0;
    3396: T492 = 1'h0;
    3397: T492 = 1'h0;
    3398: T492 = 1'h0;
    3399: T492 = 1'h0;
    3400: T492 = 1'h0;
    3401: T492 = 1'h0;
    3402: T492 = 1'h0;
    3403: T492 = 1'h0;
    3404: T492 = 1'h0;
    3405: T492 = 1'h0;
    3406: T492 = 1'h0;
    3407: T492 = 1'h0;
    3408: T492 = 1'h0;
    3409: T492 = 1'h0;
    3410: T492 = 1'h0;
    3411: T492 = 1'h0;
    3412: T492 = 1'h0;
    3413: T492 = 1'h0;
    3414: T492 = 1'h0;
    3415: T492 = 1'h0;
    3416: T492 = 1'h0;
    3417: T492 = 1'h0;
    3418: T492 = 1'h0;
    3419: T492 = 1'h0;
    3420: T492 = 1'h0;
    3421: T492 = 1'h0;
    3422: T492 = 1'h0;
    3423: T492 = 1'h0;
    3424: T492 = 1'h0;
    3425: T492 = 1'h0;
    3426: T492 = 1'h0;
    3427: T492 = 1'h0;
    3428: T492 = 1'h0;
    3429: T492 = 1'h0;
    3430: T492 = 1'h0;
    3431: T492 = 1'h0;
    3432: T492 = 1'h0;
    3433: T492 = 1'h0;
    3434: T492 = 1'h0;
    3435: T492 = 1'h0;
    3436: T492 = 1'h0;
    3437: T492 = 1'h0;
    3438: T492 = 1'h0;
    3439: T492 = 1'h0;
    3440: T492 = 1'h0;
    3441: T492 = 1'h0;
    3442: T492 = 1'h0;
    3443: T492 = 1'h0;
    3444: T492 = 1'h0;
    3445: T492 = 1'h0;
    3446: T492 = 1'h0;
    3447: T492 = 1'h0;
    3448: T492 = 1'h0;
    3449: T492 = 1'h0;
    3450: T492 = 1'h0;
    3451: T492 = 1'h0;
    3452: T492 = 1'h0;
    3453: T492 = 1'h0;
    3454: T492 = 1'h0;
    3455: T492 = 1'h0;
    3456: T492 = 1'h0;
    3457: T492 = 1'h0;
    3458: T492 = 1'h0;
    3459: T492 = 1'h0;
    3460: T492 = 1'h0;
    3461: T492 = 1'h0;
    3462: T492 = 1'h0;
    3463: T492 = 1'h0;
    3464: T492 = 1'h0;
    3465: T492 = 1'h0;
    3466: T492 = 1'h0;
    3467: T492 = 1'h0;
    3468: T492 = 1'h0;
    3469: T492 = 1'h0;
    3470: T492 = 1'h0;
    3471: T492 = 1'h0;
    3472: T492 = 1'h0;
    3473: T492 = 1'h0;
    3474: T492 = 1'h0;
    3475: T492 = 1'h0;
    3476: T492 = 1'h0;
    3477: T492 = 1'h0;
    3478: T492 = 1'h0;
    3479: T492 = 1'h0;
    3480: T492 = 1'h0;
    3481: T492 = 1'h0;
    3482: T492 = 1'h0;
    3483: T492 = 1'h0;
    3484: T492 = 1'h0;
    3485: T492 = 1'h0;
    3486: T492 = 1'h0;
    3487: T492 = 1'h0;
    3488: T492 = 1'h0;
    3489: T492 = 1'h0;
    3490: T492 = 1'h0;
    3491: T492 = 1'h0;
    3492: T492 = 1'h0;
    3493: T492 = 1'h0;
    3494: T492 = 1'h0;
    3495: T492 = 1'h0;
    3496: T492 = 1'h0;
    3497: T492 = 1'h0;
    3498: T492 = 1'h0;
    3499: T492 = 1'h0;
    3500: T492 = 1'h0;
    3501: T492 = 1'h0;
    3502: T492 = 1'h0;
    3503: T492 = 1'h0;
    3504: T492 = 1'h0;
    3505: T492 = 1'h0;
    3506: T492 = 1'h0;
    3507: T492 = 1'h0;
    3508: T492 = 1'h0;
    3509: T492 = 1'h0;
    3510: T492 = 1'h0;
    3511: T492 = 1'h0;
    3512: T492 = 1'h0;
    3513: T492 = 1'h0;
    3514: T492 = 1'h0;
    3515: T492 = 1'h0;
    3516: T492 = 1'h0;
    3517: T492 = 1'h0;
    3518: T492 = 1'h0;
    3519: T492 = 1'h0;
    3520: T492 = 1'h0;
    3521: T492 = 1'h0;
    3522: T492 = 1'h0;
    3523: T492 = 1'h0;
    3524: T492 = 1'h0;
    3525: T492 = 1'h0;
    3526: T492 = 1'h0;
    3527: T492 = 1'h0;
    3528: T492 = 1'h0;
    3529: T492 = 1'h0;
    3530: T492 = 1'h0;
    3531: T492 = 1'h0;
    3532: T492 = 1'h0;
    3533: T492 = 1'h0;
    3534: T492 = 1'h0;
    3535: T492 = 1'h0;
    3536: T492 = 1'h0;
    3537: T492 = 1'h0;
    3538: T492 = 1'h0;
    3539: T492 = 1'h0;
    3540: T492 = 1'h0;
    3541: T492 = 1'h0;
    3542: T492 = 1'h0;
    3543: T492 = 1'h0;
    3544: T492 = 1'h0;
    3545: T492 = 1'h0;
    3546: T492 = 1'h0;
    3547: T492 = 1'h0;
    3548: T492 = 1'h0;
    3549: T492 = 1'h0;
    3550: T492 = 1'h0;
    3551: T492 = 1'h0;
    3552: T492 = 1'h0;
    3553: T492 = 1'h0;
    3554: T492 = 1'h0;
    3555: T492 = 1'h0;
    3556: T492 = 1'h0;
    3557: T492 = 1'h0;
    3558: T492 = 1'h0;
    3559: T492 = 1'h0;
    3560: T492 = 1'h0;
    3561: T492 = 1'h0;
    3562: T492 = 1'h0;
    3563: T492 = 1'h0;
    3564: T492 = 1'h0;
    3565: T492 = 1'h0;
    3566: T492 = 1'h0;
    3567: T492 = 1'h0;
    3568: T492 = 1'h0;
    3569: T492 = 1'h0;
    3570: T492 = 1'h0;
    3571: T492 = 1'h0;
    3572: T492 = 1'h0;
    3573: T492 = 1'h0;
    3574: T492 = 1'h0;
    3575: T492 = 1'h0;
    3576: T492 = 1'h0;
    3577: T492 = 1'h0;
    3578: T492 = 1'h0;
    3579: T492 = 1'h0;
    3580: T492 = 1'h0;
    3581: T492 = 1'h0;
    3582: T492 = 1'h0;
    3583: T492 = 1'h0;
    3584: T492 = 1'h0;
    3585: T492 = 1'h0;
    3586: T492 = 1'h0;
    3587: T492 = 1'h0;
    3588: T492 = 1'h0;
    3589: T492 = 1'h0;
    3590: T492 = 1'h0;
    3591: T492 = 1'h0;
    3592: T492 = 1'h0;
    3593: T492 = 1'h0;
    3594: T492 = 1'h0;
    3595: T492 = 1'h0;
    3596: T492 = 1'h0;
    3597: T492 = 1'h0;
    3598: T492 = 1'h0;
    3599: T492 = 1'h0;
    3600: T492 = 1'h0;
    3601: T492 = 1'h0;
    3602: T492 = 1'h0;
    3603: T492 = 1'h0;
    3604: T492 = 1'h0;
    3605: T492 = 1'h0;
    3606: T492 = 1'h0;
    3607: T492 = 1'h0;
    3608: T492 = 1'h0;
    3609: T492 = 1'h0;
    3610: T492 = 1'h0;
    3611: T492 = 1'h0;
    3612: T492 = 1'h0;
    3613: T492 = 1'h0;
    3614: T492 = 1'h0;
    3615: T492 = 1'h0;
    3616: T492 = 1'h0;
    3617: T492 = 1'h0;
    3618: T492 = 1'h0;
    3619: T492 = 1'h0;
    3620: T492 = 1'h0;
    3621: T492 = 1'h0;
    3622: T492 = 1'h0;
    3623: T492 = 1'h0;
    3624: T492 = 1'h0;
    3625: T492 = 1'h0;
    3626: T492 = 1'h0;
    3627: T492 = 1'h0;
    3628: T492 = 1'h0;
    3629: T492 = 1'h0;
    3630: T492 = 1'h0;
    3631: T492 = 1'h0;
    3632: T492 = 1'h0;
    3633: T492 = 1'h0;
    3634: T492 = 1'h0;
    3635: T492 = 1'h0;
    3636: T492 = 1'h0;
    3637: T492 = 1'h0;
    3638: T492 = 1'h0;
    3639: T492 = 1'h0;
    3640: T492 = 1'h0;
    3641: T492 = 1'h0;
    3642: T492 = 1'h0;
    3643: T492 = 1'h0;
    3644: T492 = 1'h0;
    3645: T492 = 1'h0;
    3646: T492 = 1'h0;
    3647: T492 = 1'h0;
    3648: T492 = 1'h0;
    3649: T492 = 1'h0;
    3650: T492 = 1'h0;
    3651: T492 = 1'h0;
    3652: T492 = 1'h0;
    3653: T492 = 1'h0;
    3654: T492 = 1'h0;
    3655: T492 = 1'h0;
    3656: T492 = 1'h0;
    3657: T492 = 1'h0;
    3658: T492 = 1'h0;
    3659: T492 = 1'h0;
    3660: T492 = 1'h0;
    3661: T492 = 1'h0;
    3662: T492 = 1'h0;
    3663: T492 = 1'h0;
    3664: T492 = 1'h0;
    3665: T492 = 1'h0;
    3666: T492 = 1'h0;
    3667: T492 = 1'h0;
    3668: T492 = 1'h0;
    3669: T492 = 1'h0;
    3670: T492 = 1'h0;
    3671: T492 = 1'h0;
    3672: T492 = 1'h0;
    3673: T492 = 1'h0;
    3674: T492 = 1'h0;
    3675: T492 = 1'h0;
    3676: T492 = 1'h0;
    3677: T492 = 1'h0;
    3678: T492 = 1'h0;
    3679: T492 = 1'h0;
    3680: T492 = 1'h0;
    3681: T492 = 1'h0;
    3682: T492 = 1'h0;
    3683: T492 = 1'h0;
    3684: T492 = 1'h0;
    3685: T492 = 1'h0;
    3686: T492 = 1'h0;
    3687: T492 = 1'h0;
    3688: T492 = 1'h0;
    3689: T492 = 1'h0;
    3690: T492 = 1'h0;
    3691: T492 = 1'h0;
    3692: T492 = 1'h0;
    3693: T492 = 1'h0;
    3694: T492 = 1'h0;
    3695: T492 = 1'h0;
    3696: T492 = 1'h0;
    3697: T492 = 1'h0;
    3698: T492 = 1'h0;
    3699: T492 = 1'h0;
    3700: T492 = 1'h0;
    3701: T492 = 1'h0;
    3702: T492 = 1'h0;
    3703: T492 = 1'h0;
    3704: T492 = 1'h0;
    3705: T492 = 1'h0;
    3706: T492 = 1'h0;
    3707: T492 = 1'h0;
    3708: T492 = 1'h0;
    3709: T492 = 1'h0;
    3710: T492 = 1'h0;
    3711: T492 = 1'h0;
    3712: T492 = 1'h0;
    3713: T492 = 1'h0;
    3714: T492 = 1'h0;
    3715: T492 = 1'h0;
    3716: T492 = 1'h0;
    3717: T492 = 1'h0;
    3718: T492 = 1'h0;
    3719: T492 = 1'h0;
    3720: T492 = 1'h0;
    3721: T492 = 1'h0;
    3722: T492 = 1'h0;
    3723: T492 = 1'h0;
    3724: T492 = 1'h0;
    3725: T492 = 1'h0;
    3726: T492 = 1'h0;
    3727: T492 = 1'h0;
    3728: T492 = 1'h0;
    3729: T492 = 1'h0;
    3730: T492 = 1'h0;
    3731: T492 = 1'h0;
    3732: T492 = 1'h0;
    3733: T492 = 1'h0;
    3734: T492 = 1'h0;
    3735: T492 = 1'h0;
    3736: T492 = 1'h0;
    3737: T492 = 1'h0;
    3738: T492 = 1'h0;
    3739: T492 = 1'h0;
    3740: T492 = 1'h0;
    3741: T492 = 1'h0;
    3742: T492 = 1'h0;
    3743: T492 = 1'h0;
    3744: T492 = 1'h0;
    3745: T492 = 1'h0;
    3746: T492 = 1'h0;
    3747: T492 = 1'h0;
    3748: T492 = 1'h0;
    3749: T492 = 1'h0;
    3750: T492 = 1'h0;
    3751: T492 = 1'h0;
    3752: T492 = 1'h0;
    3753: T492 = 1'h0;
    3754: T492 = 1'h0;
    3755: T492 = 1'h0;
    3756: T492 = 1'h0;
    3757: T492 = 1'h0;
    3758: T492 = 1'h0;
    3759: T492 = 1'h0;
    3760: T492 = 1'h0;
    3761: T492 = 1'h0;
    3762: T492 = 1'h0;
    3763: T492 = 1'h0;
    3764: T492 = 1'h0;
    3765: T492 = 1'h0;
    3766: T492 = 1'h0;
    3767: T492 = 1'h0;
    3768: T492 = 1'h0;
    3769: T492 = 1'h0;
    3770: T492 = 1'h0;
    3771: T492 = 1'h0;
    3772: T492 = 1'h0;
    3773: T492 = 1'h0;
    3774: T492 = 1'h0;
    3775: T492 = 1'h0;
    3776: T492 = 1'h0;
    3777: T492 = 1'h0;
    3778: T492 = 1'h0;
    3779: T492 = 1'h0;
    3780: T492 = 1'h0;
    3781: T492 = 1'h0;
    3782: T492 = 1'h0;
    3783: T492 = 1'h0;
    3784: T492 = 1'h0;
    3785: T492 = 1'h0;
    3786: T492 = 1'h0;
    3787: T492 = 1'h0;
    3788: T492 = 1'h0;
    3789: T492 = 1'h0;
    3790: T492 = 1'h0;
    3791: T492 = 1'h0;
    3792: T492 = 1'h0;
    3793: T492 = 1'h0;
    3794: T492 = 1'h0;
    3795: T492 = 1'h0;
    3796: T492 = 1'h0;
    3797: T492 = 1'h0;
    3798: T492 = 1'h0;
    3799: T492 = 1'h0;
    3800: T492 = 1'h0;
    3801: T492 = 1'h0;
    3802: T492 = 1'h0;
    3803: T492 = 1'h0;
    3804: T492 = 1'h0;
    3805: T492 = 1'h0;
    3806: T492 = 1'h0;
    3807: T492 = 1'h0;
    3808: T492 = 1'h0;
    3809: T492 = 1'h0;
    3810: T492 = 1'h0;
    3811: T492 = 1'h0;
    3812: T492 = 1'h0;
    3813: T492 = 1'h0;
    3814: T492 = 1'h0;
    3815: T492 = 1'h0;
    3816: T492 = 1'h0;
    3817: T492 = 1'h0;
    3818: T492 = 1'h0;
    3819: T492 = 1'h0;
    3820: T492 = 1'h0;
    3821: T492 = 1'h0;
    3822: T492 = 1'h0;
    3823: T492 = 1'h0;
    3824: T492 = 1'h0;
    3825: T492 = 1'h0;
    3826: T492 = 1'h0;
    3827: T492 = 1'h0;
    3828: T492 = 1'h0;
    3829: T492 = 1'h0;
    3830: T492 = 1'h0;
    3831: T492 = 1'h0;
    3832: T492 = 1'h0;
    3833: T492 = 1'h0;
    3834: T492 = 1'h0;
    3835: T492 = 1'h0;
    3836: T492 = 1'h0;
    3837: T492 = 1'h0;
    3838: T492 = 1'h0;
    3839: T492 = 1'h0;
    3840: T492 = 1'h0;
    3841: T492 = 1'h0;
    3842: T492 = 1'h0;
    3843: T492 = 1'h0;
    3844: T492 = 1'h0;
    3845: T492 = 1'h0;
    3846: T492 = 1'h0;
    3847: T492 = 1'h0;
    3848: T492 = 1'h0;
    3849: T492 = 1'h0;
    3850: T492 = 1'h0;
    3851: T492 = 1'h0;
    3852: T492 = 1'h0;
    3853: T492 = 1'h0;
    3854: T492 = 1'h0;
    3855: T492 = 1'h0;
    3856: T492 = 1'h0;
    3857: T492 = 1'h0;
    3858: T492 = 1'h0;
    3859: T492 = 1'h0;
    3860: T492 = 1'h0;
    3861: T492 = 1'h0;
    3862: T492 = 1'h0;
    3863: T492 = 1'h0;
    3864: T492 = 1'h0;
    3865: T492 = 1'h0;
    3866: T492 = 1'h0;
    3867: T492 = 1'h0;
    3868: T492 = 1'h0;
    3869: T492 = 1'h0;
    3870: T492 = 1'h0;
    3871: T492 = 1'h0;
    3872: T492 = 1'h0;
    3873: T492 = 1'h0;
    3874: T492 = 1'h0;
    3875: T492 = 1'h0;
    3876: T492 = 1'h0;
    3877: T492 = 1'h0;
    3878: T492 = 1'h0;
    3879: T492 = 1'h0;
    3880: T492 = 1'h0;
    3881: T492 = 1'h0;
    3882: T492 = 1'h0;
    3883: T492 = 1'h0;
    3884: T492 = 1'h0;
    3885: T492 = 1'h0;
    3886: T492 = 1'h0;
    3887: T492 = 1'h0;
    3888: T492 = 1'h0;
    3889: T492 = 1'h0;
    3890: T492 = 1'h0;
    3891: T492 = 1'h0;
    3892: T492 = 1'h0;
    3893: T492 = 1'h0;
    3894: T492 = 1'h0;
    3895: T492 = 1'h0;
    3896: T492 = 1'h0;
    3897: T492 = 1'h0;
    3898: T492 = 1'h0;
    3899: T492 = 1'h0;
    3900: T492 = 1'h0;
    3901: T492 = 1'h0;
    3902: T492 = 1'h0;
    3903: T492 = 1'h0;
    3904: T492 = 1'h0;
    3905: T492 = 1'h0;
    3906: T492 = 1'h0;
    3907: T492 = 1'h0;
    3908: T492 = 1'h0;
    3909: T492 = 1'h0;
    3910: T492 = 1'h0;
    3911: T492 = 1'h0;
    3912: T492 = 1'h0;
    3913: T492 = 1'h0;
    3914: T492 = 1'h0;
    3915: T492 = 1'h0;
    3916: T492 = 1'h0;
    3917: T492 = 1'h0;
    3918: T492 = 1'h0;
    3919: T492 = 1'h0;
    3920: T492 = 1'h0;
    3921: T492 = 1'h0;
    3922: T492 = 1'h0;
    3923: T492 = 1'h0;
    3924: T492 = 1'h0;
    3925: T492 = 1'h0;
    3926: T492 = 1'h0;
    3927: T492 = 1'h0;
    3928: T492 = 1'h0;
    3929: T492 = 1'h0;
    3930: T492 = 1'h0;
    3931: T492 = 1'h0;
    3932: T492 = 1'h0;
    3933: T492 = 1'h0;
    3934: T492 = 1'h0;
    3935: T492 = 1'h0;
    3936: T492 = 1'h0;
    3937: T492 = 1'h0;
    3938: T492 = 1'h0;
    3939: T492 = 1'h0;
    3940: T492 = 1'h0;
    3941: T492 = 1'h0;
    3942: T492 = 1'h0;
    3943: T492 = 1'h0;
    3944: T492 = 1'h0;
    3945: T492 = 1'h0;
    3946: T492 = 1'h0;
    3947: T492 = 1'h0;
    3948: T492 = 1'h0;
    3949: T492 = 1'h0;
    3950: T492 = 1'h0;
    3951: T492 = 1'h0;
    3952: T492 = 1'h0;
    3953: T492 = 1'h0;
    3954: T492 = 1'h0;
    3955: T492 = 1'h0;
    3956: T492 = 1'h0;
    3957: T492 = 1'h0;
    3958: T492 = 1'h0;
    3959: T492 = 1'h0;
    3960: T492 = 1'h0;
    3961: T492 = 1'h0;
    3962: T492 = 1'h0;
    3963: T492 = 1'h0;
    3964: T492 = 1'h0;
    3965: T492 = 1'h0;
    3966: T492 = 1'h0;
    3967: T492 = 1'h0;
    3968: T492 = 1'h0;
    3969: T492 = 1'h0;
    3970: T492 = 1'h0;
    3971: T492 = 1'h0;
    3972: T492 = 1'h0;
    3973: T492 = 1'h0;
    3974: T492 = 1'h0;
    3975: T492 = 1'h0;
    3976: T492 = 1'h0;
    3977: T492 = 1'h0;
    3978: T492 = 1'h0;
    3979: T492 = 1'h0;
    3980: T492 = 1'h0;
    3981: T492 = 1'h0;
    3982: T492 = 1'h0;
    3983: T492 = 1'h0;
    3984: T492 = 1'h0;
    3985: T492 = 1'h0;
    3986: T492 = 1'h0;
    3987: T492 = 1'h0;
    3988: T492 = 1'h0;
    3989: T492 = 1'h0;
    3990: T492 = 1'h0;
    3991: T492 = 1'h0;
    3992: T492 = 1'h0;
    3993: T492 = 1'h0;
    3994: T492 = 1'h0;
    3995: T492 = 1'h0;
    3996: T492 = 1'h0;
    3997: T492 = 1'h0;
    3998: T492 = 1'h0;
    3999: T492 = 1'h0;
    4000: T492 = 1'h0;
    4001: T492 = 1'h0;
    4002: T492 = 1'h0;
    4003: T492 = 1'h0;
    4004: T492 = 1'h0;
    4005: T492 = 1'h0;
    4006: T492 = 1'h0;
    4007: T492 = 1'h0;
    4008: T492 = 1'h0;
    4009: T492 = 1'h0;
    4010: T492 = 1'h0;
    4011: T492 = 1'h0;
    4012: T492 = 1'h0;
    4013: T492 = 1'h0;
    4014: T492 = 1'h0;
    4015: T492 = 1'h0;
    4016: T492 = 1'h0;
    4017: T492 = 1'h0;
    4018: T492 = 1'h0;
    4019: T492 = 1'h0;
    4020: T492 = 1'h0;
    4021: T492 = 1'h0;
    4022: T492 = 1'h0;
    4023: T492 = 1'h0;
    4024: T492 = 1'h0;
    4025: T492 = 1'h0;
    4026: T492 = 1'h0;
    4027: T492 = 1'h0;
    4028: T492 = 1'h0;
    4029: T492 = 1'h0;
    4030: T492 = 1'h0;
    4031: T492 = 1'h0;
    4032: T492 = 1'h0;
    4033: T492 = 1'h0;
    4034: T492 = 1'h0;
    4035: T492 = 1'h0;
    4036: T492 = 1'h0;
    4037: T492 = 1'h0;
    4038: T492 = 1'h0;
    4039: T492 = 1'h0;
    4040: T492 = 1'h0;
    4041: T492 = 1'h0;
    4042: T492 = 1'h0;
    4043: T492 = 1'h0;
    4044: T492 = 1'h0;
    4045: T492 = 1'h0;
    4046: T492 = 1'h0;
    4047: T492 = 1'h0;
    4048: T492 = 1'h0;
    4049: T492 = 1'h0;
    4050: T492 = 1'h0;
    4051: T492 = 1'h0;
    4052: T492 = 1'h0;
    4053: T492 = 1'h0;
    4054: T492 = 1'h0;
    4055: T492 = 1'h0;
    4056: T492 = 1'h0;
    4057: T492 = 1'h0;
    4058: T492 = 1'h0;
    4059: T492 = 1'h0;
    4060: T492 = 1'h0;
    4061: T492 = 1'h0;
    4062: T492 = 1'h0;
    4063: T492 = 1'h0;
    4064: T492 = 1'h0;
    4065: T492 = 1'h0;
    4066: T492 = 1'h0;
    4067: T492 = 1'h0;
    4068: T492 = 1'h0;
    4069: T492 = 1'h0;
    4070: T492 = 1'h0;
    4071: T492 = 1'h0;
    4072: T492 = 1'h0;
    4073: T492 = 1'h0;
    4074: T492 = 1'h0;
    4075: T492 = 1'h0;
    4076: T492 = 1'h0;
    4077: T492 = 1'h0;
    4078: T492 = 1'h0;
    4079: T492 = 1'h0;
    4080: T492 = 1'h0;
    4081: T492 = 1'h0;
    4082: T492 = 1'h0;
    4083: T492 = 1'h0;
    4084: T492 = 1'h0;
    4085: T492 = 1'h0;
    4086: T492 = 1'h0;
    4087: T492 = 1'h0;
    4088: T492 = 1'h0;
    4089: T492 = 1'h0;
    4090: T492 = 1'h0;
    4091: T492 = 1'h0;
    4092: T492 = 1'h0;
    4093: T492 = 1'h0;
    4094: T492 = 1'h0;
    4095: T492 = 1'h0;
`ifndef SYNTHESIS
    default: T492 = {1{$random}};
`else
    default: T492 = 1'bx;
`endif
  endcase
  assign T494 = id_int_val ^ 1'h1;
  assign id_int_val = T497 | T495;
  assign T495 = T496 == 32'h3;
  assign T496 = io_dpath_inst & 32'h7067;
  assign T497 = T500 | T498;
  assign T498 = T499 == 32'h33;
  assign T499 = io_dpath_inst & 32'hfc007077;
  assign T500 = T503 | T501;
  assign T501 = T502 == 32'h4063;
  assign T502 = io_dpath_inst & 32'h407f;
  assign T503 = T506 | T504;
  assign T504 = T505 == 32'h1063;
  assign T505 = io_dpath_inst & 32'h306f;
  assign T506 = T509 | T507;
  assign T507 = T508 == 32'h23;
  assign T508 = io_dpath_inst & 32'h603f;
  assign T509 = T512 | T510;
  assign T510 = T511 == 32'he0000053;
  assign T511 = io_dpath_inst & 32'hedf0707f;
  assign T512 = T515 | T513;
  assign T513 = T514 == 32'he0000053;
  assign T514 = io_dpath_inst & 32'hfdf0607f;
  assign T515 = T518 | T516;
  assign T516 = T517 == 32'hc0000053;
  assign T517 = io_dpath_inst & 32'hedc0007f;
  assign T518 = T521 | T519;
  assign T519 = T520 == 32'h42000053;
  assign T520 = io_dpath_inst & 32'h7ff0007f;
  assign T521 = T524 | T522;
  assign T522 = T523 == 32'h40100053;
  assign T523 = io_dpath_inst & 32'h7ff0007f;
  assign T524 = T527 | T525;
  assign T525 = T526 == 32'h20000053;
  assign T526 = io_dpath_inst & 32'h7c00507f;
  assign T527 = T530 | T528;
  assign T528 = T529 == 32'h20000053;
  assign T529 = io_dpath_inst & 32'h7c00607f;
  assign T530 = T533 | T531;
  assign T531 = T532 == 32'h20000053;
  assign T532 = io_dpath_inst & 32'hf400607f;
  assign T533 = T534 | T69;
  assign T534 = T535 | T72;
  assign T535 = T538 | T536;
  assign T536 = T537 == 32'h2004033;
  assign T537 = io_dpath_inst & 32'hfe004077;
  assign T538 = T541 | T539;
  assign T539 = T540 == 32'h5033;
  assign T540 = io_dpath_inst & 32'hbe007077;
  assign T541 = T544 | T542;
  assign T542 = T543 == 32'h501b;
  assign T543 = io_dpath_inst & 32'hbe00705f;
  assign T544 = T547 | T545;
  assign T545 = T546 == 32'h5013;
  assign T546 = io_dpath_inst & 32'hbc00707f;
  assign T547 = T550 | T548;
  assign T548 = T549 == 32'h2073;
  assign T549 = io_dpath_inst & 32'h2077;
  assign T550 = T553 | T551;
  assign T551 = T552 == 32'h205b;
  assign T552 = io_dpath_inst & 32'h205f;
  assign T553 = T554 | T75;
  assign T554 = T557 | T555;
  assign T555 = T556 == 32'h2013;
  assign T556 = io_dpath_inst & 32'h207f;
  assign T557 = T560 | T558;
  assign T558 = T559 == 32'h200b;
  assign T559 = io_dpath_inst & 32'h205f;
  assign T560 = T561 | T78;
  assign T561 = T564 | T562;
  assign T562 = T563 == 32'h101b;
  assign T563 = io_dpath_inst & 32'hfe00305f;
  assign T564 = T567 | T565;
  assign T565 = T566 == 32'h1013;
  assign T566 = io_dpath_inst & 32'hfc00305f;
  assign T567 = T570 | T568;
  assign T568 = T569 == 32'h73;
  assign T569 = io_dpath_inst & 32'h7fffffff;
  assign T570 = T573 | T571;
  assign T571 = T572 == 32'h6f;
  assign T572 = io_dpath_inst & 32'h7f;
  assign T573 = T576 | T574;
  assign T574 = T575 == 32'h63;
  assign T575 = io_dpath_inst & 32'h707b;
  assign T576 = T579 | T577;
  assign T577 = T578 == 32'h5b;
  assign T578 = io_dpath_inst & 32'h105f;
  assign T579 = T582 | T580;
  assign T580 = T581 == 32'h53;
  assign T581 = io_dpath_inst & 32'hec00007f;
  assign T582 = T585 | T583;
  assign T583 = T584 == 32'h53;
  assign T584 = io_dpath_inst & 32'hf400007f;
  assign T585 = T588 | T586;
  assign T586 = T587 == 32'h43;
  assign T587 = io_dpath_inst & 32'h4000073;
  assign T588 = T591 | T589;
  assign T589 = T590 == 32'h33;
  assign T590 = io_dpath_inst & 32'hbe007077;
  assign T591 = T594 | T592;
  assign T592 = T593 == 32'h33;
  assign T593 = io_dpath_inst & 32'hfc00007f;
  assign T594 = T597 | T595;
  assign T595 = T596 == 32'h17;
  assign T596 = io_dpath_inst & 32'h5f;
  assign T597 = T600 | T598;
  assign T598 = T599 == 32'hf;
  assign T599 = io_dpath_inst & 32'h607f;
  assign T600 = T603 | T601;
  assign T601 = T602 == 32'hb;
  assign T602 = io_dpath_inst & 32'h105f;
  assign T603 = T84 | T604;
  assign T604 = T605 == 32'h3;
  assign T605 = io_dpath_inst & 32'h106f;
  assign T606 = T607 | io_imem_resp_bits_xcpt_if;
  assign T607 = id_interrupt | io_imem_resp_bits_xcpt_ma;
  assign T608 = T609 & io_imem_resp_valid;
  assign T609 = id_interrupt & T610;
  assign T610 = take_pc ^ 1'h1;
  assign T611 = dcache_kill_mem | take_pc_wb;
  assign T612 = replay_wb | wb_reg_xcpt;
  assign mem_xcpt = T614 | T613;
  assign T613 = mem_reg_mem_val & io_dmem_xcpt_pf_st;
  assign T614 = T616 | T615;
  assign T615 = mem_reg_mem_val & io_dmem_xcpt_pf_ld;
  assign T616 = T618 | T617;
  assign T617 = mem_reg_mem_val & io_dmem_xcpt_ma_st;
  assign T618 = T620 | T619;
  assign T619 = mem_reg_mem_val & io_dmem_xcpt_ma_ld;
  assign T620 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T621 = T623 & T622;
  assign T622 = mem_reg_replay_next ^ 1'h1;
  assign T623 = T624 & ex_reg_xcpt_interrupt;
  assign T624 = take_pc ^ 1'h1;
  assign io_rocc_s = io_dpath_status_s;
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = wb_reg_rocc_val & T625;
  assign T625 = replay_wb_common ^ 1'h1;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T626;
  assign T626 = T627 & id_fp_val;
  assign T627 = ctrl_killd ^ 1'h1;
  assign io_dmem_req_bits_cmd = ex_reg_mem_cmd;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_typ = ex_reg_mem_type;
  assign io_dmem_req_bits_kill = T628;
  assign T628 = killm_common | mem_xcpt;
  assign io_dmem_req_valid = ex_reg_mem_val;
  assign io_imem_invalidate = wb_reg_flush_inst;
  assign T629 = ctrl_killm ? 1'h0 : mem_reg_flush_inst;
  assign T630 = ctrl_killx ? 1'h0 : ex_reg_flush_inst;
  assign T631 = ctrl_killd ? 1'h0 : id_fence_i;
  assign io_imem_btb_update_bits_mispredict = take_pc_mem;
  assign io_imem_btb_update_bits_isReturn = T632;
  assign T632 = mem_reg_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_btb_update_bits_isCall = T633;
  assign T633 = mem_reg_wen & T634;
  assign T634 = io_dpath_mem_waddr[1'h0:1'h0];
  assign io_imem_btb_update_bits_isJump = T635;
  assign T635 = mem_reg_jal | mem_reg_jalr;
  assign io_imem_btb_update_bits_taken = T636;
  assign T636 = T637 | io_imem_btb_update_bits_isJump;
  assign T637 = mem_reg_branch & io_dpath_mem_br_taken;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T638 = T641 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T639 = T640 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T640 = T348 & io_imem_btb_resp_valid;
  assign T641 = T380 & ex_reg_btb_hit;
  assign T642 = ctrl_killd ? 1'h0 : io_imem_btb_resp_valid;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T643 = T641 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T644 = T640 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T645 = T641 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T646 = T640 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T647 = T641 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T648 = T640 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T649 = T641 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T650 = T640 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T651 = T380 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T652;
  assign T652 = T654 & T653;
  assign T653 = take_pc_wb ^ 1'h1;
  assign T654 = mem_reg_branch | io_imem_btb_update_bits_isJump;
  assign io_imem_resp_ready = T655;
  assign T655 = T656 | ctrl_draind;
  assign T656 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_valid = take_pc;
  assign io_dpath_badvaddr_wen = wb_reg_xcpt;
  assign io_dpath_cause = wb_reg_cause;
  assign T657 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T620 ? mem_reg_cause : T841;
  assign T841 = {60'h0, T658};
  assign T658 = T619 ? 4'h8 : T659;
  assign T659 = T617 ? 4'h9 : T660;
  assign T660 = T615 ? 4'ha : 4'hb;
  assign T661 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T453 ? ex_reg_cause : 64'h2;
  assign T662 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = id_interrupt ? id_interrupt_cause : T842;
  assign T842 = {60'h0, T663};
  assign T663 = io_imem_resp_bits_xcpt_ma ? 4'h0 : T664;
  assign T664 = io_imem_resp_bits_xcpt_if ? 4'h1 : T665;
  assign T665 = T490 ? 4'h2 : T666;
  assign T666 = id_csr_privileged ? 4'h3 : T667;
  assign T667 = T466 ? 4'h3 : T668;
  assign T668 = T460 ? 4'h4 : T669;
  assign T669 = id_syscall ? 4'h6 : 4'hc;
  assign id_interrupt_cause = T56 ? 64'h8000000000000000 : T670;
  assign T670 = T53 ? 64'h8000000000000001 : T671;
  assign T671 = T49 ? 64'h8000000000000002 : T672;
  assign T672 = T45 ? 64'h8000000000000003 : T673;
  assign T673 = T41 ? 64'h8000000000000004 : T674;
  assign T674 = T37 ? 64'h8000000000000005 : T675;
  assign T675 = T33 ? 64'h8000000000000006 : 64'h8000000000000007;
  assign io_dpath_exception = wb_reg_xcpt;
  assign io_dpath_retire = T676;
  assign T676 = wb_reg_valid & T677;
  assign T677 = replay_wb ^ 1'h1;
  assign T678 = ctrl_killm ? 1'h0 : mem_reg_valid;
  assign io_dpath_ll_ready = T679;
  assign T679 = wb_reg_wen ^ 1'h1;
  assign io_dpath_bypass_src_0 = T680;
  assign T680 = T689 ? 2'h0 : T681;
  assign T681 = T687 ? 2'h1 : T682;
  assign T682 = T683 ? 2'h2 : 2'h3;
  assign T683 = T685 & T684;
  assign T684 = io_dpath_mem_waddr == id_raddr1;
  assign T685 = mem_reg_wen & T686;
  assign T686 = mem_reg_mem_val ^ 1'h1;
  assign T687 = ex_reg_wen & T688;
  assign T688 = io_dpath_ex_waddr == id_raddr1;
  assign T689 = 5'h0 == id_raddr1;
  assign io_dpath_bypass_src_1 = T690;
  assign T690 = T697 ? 2'h0 : T691;
  assign T691 = T695 ? 2'h1 : T692;
  assign T692 = T693 ? 2'h2 : 2'h3;
  assign T693 = T685 & T694;
  assign T694 = io_dpath_mem_waddr == id_raddr2;
  assign T695 = ex_reg_wen & T696;
  assign T696 = io_dpath_ex_waddr == id_raddr2;
  assign T697 = 5'h0 == id_raddr2;
  assign io_dpath_bypass_0 = T698;
  assign T698 = T701 | T699;
  assign T699 = mem_reg_wen & T700;
  assign T700 = io_dpath_mem_waddr == id_raddr1;
  assign T701 = T702 | T683;
  assign T702 = T689 | T687;
  assign io_dpath_bypass_1 = T703;
  assign T703 = T706 | T704;
  assign T704 = mem_reg_wen & T705;
  assign T705 = io_dpath_mem_waddr == id_raddr2;
  assign T706 = T707 | T693;
  assign T707 = T697 | T695;
  assign io_dpath_mem_rocc_val = mem_reg_rocc_val;
  assign io_dpath_ex_rocc_val = ex_reg_rocc_val;
  assign io_dpath_ex_rs2_val = T708;
  assign T708 = T709 | ex_reg_rocc_val;
  assign T709 = ex_reg_mem_val & T710;
  assign T710 = T714 | T711;
  assign T711 = T713 | T712;
  assign T712 = ex_reg_mem_cmd == 5'h4;
  assign T713 = ex_reg_mem_cmd[2'h3:2'h3];
  assign T714 = T716 | T715;
  assign T715 = ex_reg_mem_cmd == 5'h7;
  assign T716 = ex_reg_mem_cmd == 5'h1;
  assign io_dpath_ex_mem_type = ex_reg_mem_type;
  assign io_dpath_wb_wen = T717;
  assign T717 = wb_reg_wen & T718;
  assign T718 = replay_wb ^ 1'h1;
  assign io_dpath_mem_wen = mem_reg_wen;
  assign io_dpath_mem_branch = mem_reg_branch;
  assign io_dpath_mem_jalr = mem_reg_jalr;
  assign io_dpath_ex_valid = ex_reg_valid;
  assign io_dpath_ex_wen = ex_reg_wen;
  assign io_dpath_mem_fp_val = mem_reg_fp_val;
  assign io_dpath_ex_fp_val = ex_reg_fp_val;
  assign io_dpath_wb_load = T719;
  assign T719 = wb_reg_mem_val & wb_reg_wen;
  assign io_dpath_mem_load = T720;
  assign T720 = mem_reg_mem_val & mem_reg_wen;
  assign io_dpath_sret = wb_reg_sret;
  assign io_dpath_csr = T843;
  assign T843 = {1'h0, wb_reg_csr};
  assign T721 = ctrl_killm ? 2'h0 : mem_reg_csr;
  assign io_dpath_div_mul_kill = T722;
  assign T722 = mem_reg_div_mul_val & killm_common;
  assign io_dpath_div_mul_val = ex_reg_div_mul_val;
  assign io_dpath_fn_alu = T723;
  assign T723 = id_fn_alu;
  assign id_fn_alu = {T759, T724};
  assign T724 = {T748, T725};
  assign T725 = {T734, T726};
  assign T726 = T729 | T727;
  assign T727 = T728 == 32'h5010;
  assign T728 = io_dpath_inst & 32'h5054;
  assign T729 = T732 | T730;
  assign T730 = T731 == 32'h1040;
  assign T731 = io_dpath_inst & 32'h1058;
  assign T732 = T733 == 32'h1010;
  assign T733 = io_dpath_inst & 32'h3054;
  assign T734 = T737 | T735;
  assign T735 = T736 == 32'h40001010;
  assign T736 = io_dpath_inst & 32'h40001054;
  assign T737 = T740 | T738;
  assign T738 = T739 == 32'h40000030;
  assign T739 = io_dpath_inst & 32'h40000074;
  assign T740 = T743 | T741;
  assign T741 = T742 == 32'h6010;
  assign T742 = io_dpath_inst & 32'h6054;
  assign T743 = T746 | T744;
  assign T744 = T745 == 32'h3010;
  assign T745 = io_dpath_inst & 32'h3054;
  assign T746 = T747 == 32'h2040;
  assign T747 = io_dpath_inst & 32'h2058;
  assign T748 = T751 | T749;
  assign T749 = T750 == 32'h4040;
  assign T750 = io_dpath_inst & 32'h4058;
  assign T751 = T754 | T752;
  assign T752 = T753 == 32'h4010;
  assign T753 = io_dpath_inst & 32'h5054;
  assign T754 = T757 | T755;
  assign T755 = T756 == 32'h4010;
  assign T756 = io_dpath_inst & 32'h40004054;
  assign T757 = T758 == 32'h2010;
  assign T758 = io_dpath_inst & 32'h2054;
  assign T759 = T762 | T760;
  assign T760 = T761 == 32'h40001010;
  assign T761 = io_dpath_inst & 32'h40003054;
  assign T762 = T763 | T738;
  assign T763 = T766 | T764;
  assign T764 = T765 == 32'h2010;
  assign T765 = io_dpath_inst & 32'h6054;
  assign T766 = T767 == 32'h40;
  assign T767 = io_dpath_inst & 32'h54;
  assign io_dpath_fn_dw = T768;
  assign T768 = id_fn_dw;
  assign id_fn_dw = T771 | T769;
  assign T769 = T770 == 32'h40;
  assign T770 = io_dpath_inst & 32'h40;
  assign T771 = T774 | T772;
  assign T772 = T773 == 32'h0;
  assign T773 = io_dpath_inst & 32'h8;
  assign T774 = T775 == 32'h0;
  assign T775 = io_dpath_inst & 32'h10;
  assign io_dpath_sel_imm = T776;
  assign T776 = id_sel_imm;
  assign id_sel_imm = {T786, T777};
  assign T777 = {T783, T778};
  assign T778 = T781 | T779;
  assign T779 = T780 == 32'h40;
  assign T780 = io_dpath_inst & 32'h44;
  assign T781 = T782 == 32'h8;
  assign T782 = io_dpath_inst & 32'h18;
  assign T783 = T781 | T784;
  assign T784 = T785 == 32'h14;
  assign T785 = io_dpath_inst & 32'h14;
  assign T786 = T789 | T787;
  assign T787 = T788 == 32'h10;
  assign T788 = io_dpath_inst & 32'h14;
  assign T789 = T792 | T790;
  assign T790 = T791 == 32'h4;
  assign T791 = io_dpath_inst & 32'h201c;
  assign T792 = T793 == 32'h0;
  assign T793 = io_dpath_inst & 32'h30;
  assign io_dpath_sel_alu1 = T794;
  assign T794 = id_sel_alu1;
  assign id_sel_alu1 = {T812, T795};
  assign T795 = T798 | T796;
  assign T796 = T797 == 32'h8;
  assign T797 = io_dpath_inst & 32'hc;
  assign T798 = T801 | T799;
  assign T799 = T800 == 32'h0;
  assign T800 = io_dpath_inst & 32'h18;
  assign T801 = T804 | T802;
  assign T802 = T803 == 32'h0;
  assign T803 = io_dpath_inst & 32'h24;
  assign T804 = T807 | T805;
  assign T805 = T806 == 32'h0;
  assign T806 = io_dpath_inst & 32'h44;
  assign T807 = T810 | T808;
  assign T808 = T809 == 32'h0;
  assign T809 = io_dpath_inst & 32'h50;
  assign T810 = T811 == 32'h0;
  assign T811 = io_dpath_inst & 32'h4004;
  assign T812 = T815 | T813;
  assign T813 = T814 == 32'h48;
  assign T814 = io_dpath_inst & 32'h58;
  assign T815 = T816 == 32'h14;
  assign T816 = io_dpath_inst & 32'h34;
  assign io_dpath_sel_alu2 = T844;
  assign T844 = {1'h0, T817};
  assign T817 = id_sel_alu2;
  assign id_sel_alu2 = {T828, T818};
  assign T818 = T821 | T819;
  assign T819 = T820 == 32'h4050;
  assign T820 = io_dpath_inst & 32'h4058;
  assign T821 = T822 | T813;
  assign T822 = T825 | T823;
  assign T823 = T824 == 32'h10;
  assign T824 = io_dpath_inst & 32'h70;
  assign T825 = T270 | T826;
  assign T826 = T827 == 32'h4;
  assign T827 = io_dpath_inst & 32'hc;
  assign T828 = T831 | T829;
  assign T829 = T830 == 32'h4000;
  assign T830 = io_dpath_inst & 32'h4008;
  assign T831 = T799 | T158;
  assign io_dpath_ren_0 = id_renx1;
  assign io_dpath_ren_1 = id_renx2;
  assign io_dpath_killd = T832;
  assign T832 = take_pc | T833;
  assign T833 = ctrl_stalld & T834;
  assign T834 = ctrl_draind ^ 1'h1;
  assign io_dpath_sel_pc = T845;
  assign T845 = {1'h0, T835};
  assign T835 = wb_reg_xcpt ? 2'h3 : T836;
  assign T836 = wb_reg_sret ? 2'h3 : T837;
  assign T837 = replay_wb ? 2'h2 : 2'h1;

  always @(posedge clk) begin
    wb_reg_xcpt <= T1;
    if(ctrl_killm) begin
      wb_reg_sret <= 1'h0;
    end else begin
      wb_reg_sret <= T5;
    end
    mem_reg_replay <= T7;
    if(ctrl_killx) begin
      mem_reg_replay_next <= 1'h0;
    end else begin
      mem_reg_replay_next <= ex_reg_replay_next;
    end
    if(ctrl_killd) begin
      ex_reg_replay_next <= 1'h0;
    end else begin
      ex_reg_replay_next <= T10;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T88;
    end
    if(ctrl_killd) begin
      ex_reg_mem_val <= 1'h0;
    end else begin
      ex_reg_mem_val <= T97;
    end
    if(ctrl_killm) begin
      wb_reg_rocc_val <= 1'h0;
    end else begin
      wb_reg_rocc_val <= mem_reg_rocc_val;
    end
    if(ctrl_killx) begin
      mem_reg_rocc_val <= 1'h0;
    end else begin
      mem_reg_rocc_val <= ex_reg_rocc_val;
    end
    if(ctrl_killd) begin
      ex_reg_rocc_val <= 1'h0;
    end else begin
      ex_reg_rocc_val <= T103;
    end
    if(reset) begin
      R118 <= 32'h0;
    end else if(T180) begin
      R118 <= T176;
    end else if(T175) begin
      R118 <= T171;
    end else if(T125) begin
      R118 <= T122;
    end
    wb_reg_replay <= T130;
    if(ctrl_killx) begin
      mem_reg_fp_val <= 1'h0;
    end else begin
      mem_reg_fp_val <= ex_reg_fp_val;
    end
    if(ctrl_killd) begin
      ex_reg_fp_val <= 1'h0;
    end else begin
      ex_reg_fp_val <= id_fp_val;
    end
    if(ctrl_killx) begin
      mem_reg_wen <= 1'h0;
    end else begin
      mem_reg_wen <= ex_reg_wen;
    end
    if(ctrl_killd) begin
      ex_reg_wen <= 1'h0;
    end else begin
      ex_reg_wen <= id_wen;
    end
    if(ctrl_killm) begin
      wb_reg_fp_wen <= 1'h0;
    end else begin
      wb_reg_fp_wen <= mem_reg_fp_wen;
    end
    if(ctrl_killx) begin
      mem_reg_fp_wen <= 1'h0;
    end else begin
      mem_reg_fp_wen <= ex_reg_fp_wen;
    end
    if(ctrl_killd) begin
      ex_reg_fp_wen <= 1'h0;
    end else begin
      ex_reg_fp_wen <= T167;
    end
    if(ctrl_killm) begin
      wb_reg_mem_val <= 1'h0;
    end else begin
      wb_reg_mem_val <= mem_reg_mem_val;
    end
    if(ctrl_killx) begin
      mem_reg_mem_val <= 1'h0;
    end else begin
      mem_reg_mem_val <= ex_reg_mem_val;
    end
    if(reset) begin
      R226 <= 32'h0;
    end else if(T240) begin
      R226 <= T229;
    end else if(io_dpath_ll_wen) begin
      R226 <= T222;
    end
    if(ctrl_killm) begin
      wb_reg_div_mul_val <= 1'h0;
    end else begin
      wb_reg_div_mul_val <= mem_reg_div_mul_val;
    end
    mem_reg_div_mul_val <= T235;
    if(ctrl_killd) begin
      ex_reg_div_mul_val <= 1'h0;
    end else begin
      ex_reg_div_mul_val <= T237;
    end
    if(ctrl_killm) begin
      wb_reg_fp_val <= 1'h0;
    end else begin
      wb_reg_fp_val <= mem_reg_fp_val;
    end
    if(ctrl_killm) begin
      wb_reg_wen <= 1'h0;
    end else begin
      wb_reg_wen <= mem_reg_wen;
    end
    if(T380) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T348) begin
      ex_reg_mem_type <= T340;
    end
    if(T348) begin
      ex_reg_mem_cmd <= id_mem_cmd;
    end
    if(ctrl_killx) begin
      mem_reg_csr <= 2'h0;
    end else begin
      mem_reg_csr <= ex_reg_csr;
    end
    if(ctrl_killd) begin
      ex_reg_csr <= 2'h0;
    end else begin
      ex_reg_csr <= id_csr;
    end
    if(ctrl_killd) begin
      ex_reg_jalr <= 1'h0;
    end else begin
      ex_reg_jalr <= id_jalr;
    end
    if(ctrl_killx) begin
      mem_reg_jal <= 1'h0;
    end else begin
      mem_reg_jal <= ex_reg_jal;
    end
    if(ctrl_killd) begin
      ex_reg_jal <= 1'h0;
    end else begin
      ex_reg_jal <= id_jal;
    end
    if(ctrl_killx) begin
      mem_reg_jalr <= 1'h0;
    end else begin
      mem_reg_jalr <= ex_reg_jalr;
    end
    if(ctrl_killx) begin
      mem_reg_branch <= 1'h0;
    end else begin
      mem_reg_branch <= ex_reg_branch;
    end
    if(ctrl_killd) begin
      ex_reg_branch <= 1'h0;
    end else begin
      ex_reg_branch <= id_branch;
    end
    if(ctrl_killd) begin
      ex_reg_load_use <= 1'h0;
    end else begin
      ex_reg_load_use <= id_load_use;
    end
    if(ctrl_killx) begin
      mem_reg_sret <= 1'h0;
    end else begin
      mem_reg_sret <= ex_reg_sret;
    end
    if(ctrl_killd) begin
      ex_reg_sret <= 1'h0;
    end else begin
      ex_reg_sret <= id_sret;
    end
    if(ctrl_killx) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ex_reg_valid;
    end
    if(ctrl_killd) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= 1'h1;
    end
    if(ctrl_killx) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ex_xcpt;
    end
    if(ctrl_killd) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= id_xcpt;
    end
    ex_reg_xcpt_interrupt <= T608;
    mem_reg_xcpt_interrupt <= T621;
    if(ctrl_killm) begin
      wb_reg_flush_inst <= 1'h0;
    end else begin
      wb_reg_flush_inst <= mem_reg_flush_inst;
    end
    if(ctrl_killx) begin
      mem_reg_flush_inst <= 1'h0;
    end else begin
      mem_reg_flush_inst <= ex_reg_flush_inst;
    end
    if(ctrl_killd) begin
      ex_reg_flush_inst <= 1'h0;
    end else begin
      ex_reg_flush_inst <= id_fence_i;
    end
    if(T641) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T640) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(ctrl_killd) begin
      ex_reg_btb_hit <= 1'h0;
    end else begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T641) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T640) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T641) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T640) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T641) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T640) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T641) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T640) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T380) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(ctrl_killm) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= mem_reg_valid;
    end
    if(ctrl_killm) begin
      wb_reg_csr <= 2'h0;
    end else begin
      wb_reg_csr <= mem_reg_csr;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T133;
  wire cmp;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] T29;
  wire T30;
  wire[63:0] shout_l;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[62:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[61:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[59:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[55:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[47:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T134;
  wire[31:0] T55;
  wire[63:0] T56;
  wire[63:0] T135;
  wire[47:0] T57;
  wire[63:0] T58;
  wire[63:0] T136;
  wire[55:0] T59;
  wire[63:0] T60;
  wire[63:0] T137;
  wire[59:0] T61;
  wire[63:0] T62;
  wire[63:0] T138;
  wire[61:0] T63;
  wire[63:0] T64;
  wire[63:0] T139;
  wire[62:0] T65;
  wire T66;
  wire[63:0] shout_r;
  wire[64:0] T67;
  wire[5:0] shamt;
  wire[5:0] T68;
  wire[4:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[64:0] T73;
  wire[64:0] T74;
  wire[63:0] shin;
  wire[63:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[62:0] T78;
  wire[63:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[61:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[59:0] T86;
  wire[63:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[55:0] T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[47:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[31:0] T98;
  wire[63:0] T99;
  wire[63:0] T140;
  wire[31:0] T100;
  wire[63:0] T101;
  wire[63:0] T141;
  wire[47:0] T102;
  wire[63:0] T103;
  wire[63:0] T142;
  wire[55:0] T104;
  wire[63:0] T105;
  wire[63:0] T143;
  wire[59:0] T106;
  wire[63:0] T107;
  wire[63:0] T144;
  wire[61:0] T108;
  wire[63:0] T109;
  wire[63:0] T145;
  wire[62:0] T110;
  wire[63:0] shin_r;
  wire[31:0] T111;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T112;
  wire[31:0] T146;
  wire T113;
  wire T114;
  wire[31:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[31:0] out_hi;
  wire[31:0] T129;
  wire[31:0] T147;
  wire T130;
  wire[31:0] T131;
  wire T132;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T126 ? sum : T6;
  assign T6 = T123 ? shout_r : T7;
  assign T7 = T66 ? shout_l : T8;
  assign T8 = T30 ? T29 : T9;
  assign T9 = T28 ? T27 : T10;
  assign T10 = T26 ? T25 : T133;
  assign T133 = {63'h0, cmp};
  assign cmp = T24 ^ T11;
  assign T11 = T22 ? T21 : T12;
  assign T12 = T18 ? T17 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = io_in1[6'h3f:6'h3f];
  assign T15 = io_in2[6'h3f:6'h3f];
  assign T16 = io_fn[1'h1:1'h1];
  assign T17 = sum[6'h3f:6'h3f];
  assign T18 = T20 == T19;
  assign T19 = io_in2[6'h3f:6'h3f];
  assign T20 = io_in1[6'h3f:6'h3f];
  assign T21 = sum == 64'h0;
  assign T22 = T23 ^ 1'h1;
  assign T23 = io_fn[2'h2:2'h2];
  assign T24 = io_fn[1'h0:1'h0];
  assign T25 = io_in1 ^ io_in2;
  assign T26 = io_fn == 4'h4;
  assign T27 = io_in1 | io_in2;
  assign T28 = io_fn == 4'h6;
  assign T29 = io_in1 & io_in2;
  assign T30 = io_fn == 4'h7;
  assign shout_l = T64 | T31;
  assign T31 = T32 & 64'haaaaaaaaaaaaaaaa;
  assign T32 = T33 << 1'h1;
  assign T33 = T34[6'h3e:1'h0];
  assign T34 = T62 | T35;
  assign T35 = T36 & 64'hcccccccccccccccc;
  assign T36 = T37 << 2'h2;
  assign T37 = T38[6'h3d:1'h0];
  assign T38 = T60 | T39;
  assign T39 = T40 & 64'hf0f0f0f0f0f0f0f0;
  assign T40 = T41 << 3'h4;
  assign T41 = T42[6'h3b:1'h0];
  assign T42 = T58 | T43;
  assign T43 = T44 & 64'hff00ff00ff00ff00;
  assign T44 = T45 << 4'h8;
  assign T45 = T46[6'h37:1'h0];
  assign T46 = T56 | T47;
  assign T47 = T48 & 64'hffff0000ffff0000;
  assign T48 = T49 << 5'h10;
  assign T49 = T50[6'h2f:1'h0];
  assign T50 = T54 | T51;
  assign T51 = T52 & 64'hffffffff00000000;
  assign T52 = T53 << 6'h20;
  assign T53 = shout_r[5'h1f:1'h0];
  assign T54 = T134 & 64'hffffffff;
  assign T134 = {32'h0, T55};
  assign T55 = shout_r >> 6'h20;
  assign T56 = T135 & 64'hffff0000ffff;
  assign T135 = {16'h0, T57};
  assign T57 = T50 >> 5'h10;
  assign T58 = T136 & 64'hff00ff00ff00ff;
  assign T136 = {8'h0, T59};
  assign T59 = T46 >> 4'h8;
  assign T60 = T137 & 64'hf0f0f0f0f0f0f0f;
  assign T137 = {4'h0, T61};
  assign T61 = T42 >> 3'h4;
  assign T62 = T138 & 64'h3333333333333333;
  assign T138 = {2'h0, T63};
  assign T63 = T38 >> 2'h2;
  assign T64 = T139 & 64'h5555555555555555;
  assign T139 = {1'h0, T65};
  assign T65 = T34 >> 1'h1;
  assign T66 = io_fn == 4'h1;
  assign shout_r = T67[6'h3f:1'h0];
  assign T67 = $signed(T73) >>> shamt;
  assign shamt = T68;
  assign T68 = {T70, T69};
  assign T69 = io_in2[3'h4:1'h0];
  assign T70 = T72 & T71;
  assign T71 = io_dw == 1'h1;
  assign T72 = io_in2[3'h5:3'h5];
  assign T73 = T74;
  assign T74 = {T120, shin};
  assign shin = T117 ? shin_r : T75;
  assign T75 = T109 | T76;
  assign T76 = T77 & 64'haaaaaaaaaaaaaaaa;
  assign T77 = T78 << 1'h1;
  assign T78 = T79[6'h3e:1'h0];
  assign T79 = T107 | T80;
  assign T80 = T81 & 64'hcccccccccccccccc;
  assign T81 = T82 << 2'h2;
  assign T82 = T83[6'h3d:1'h0];
  assign T83 = T105 | T84;
  assign T84 = T85 & 64'hf0f0f0f0f0f0f0f0;
  assign T85 = T86 << 3'h4;
  assign T86 = T87[6'h3b:1'h0];
  assign T87 = T103 | T88;
  assign T88 = T89 & 64'hff00ff00ff00ff00;
  assign T89 = T90 << 4'h8;
  assign T90 = T91[6'h37:1'h0];
  assign T91 = T101 | T92;
  assign T92 = T93 & 64'hffff0000ffff0000;
  assign T93 = T94 << 5'h10;
  assign T94 = T95[6'h2f:1'h0];
  assign T95 = T99 | T96;
  assign T96 = T97 & 64'hffffffff00000000;
  assign T97 = T98 << 6'h20;
  assign T98 = shin_r[5'h1f:1'h0];
  assign T99 = T140 & 64'hffffffff;
  assign T140 = {32'h0, T100};
  assign T100 = shin_r >> 6'h20;
  assign T101 = T141 & 64'hffff0000ffff;
  assign T141 = {16'h0, T102};
  assign T102 = T95 >> 5'h10;
  assign T103 = T142 & 64'hff00ff00ff00ff;
  assign T142 = {8'h0, T104};
  assign T104 = T91 >> 4'h8;
  assign T105 = T143 & 64'hf0f0f0f0f0f0f0f;
  assign T143 = {4'h0, T106};
  assign T106 = T87 >> 3'h4;
  assign T107 = T144 & 64'h3333333333333333;
  assign T144 = {2'h0, T108};
  assign T108 = T83 >> 2'h2;
  assign T109 = T145 & 64'h5555555555555555;
  assign T145 = {1'h0, T110};
  assign T110 = T79 >> 1'h1;
  assign shin_r = {shin_hi, T111};
  assign T111 = io_in1[5'h1f:1'h0];
  assign shin_hi = T116 ? T115 : shin_hi_32;
  assign shin_hi_32 = T114 ? T112 : 32'h0;
  assign T112 = 32'h0 - T146;
  assign T146 = {31'h0, T113};
  assign T113 = io_in1[5'h1f:5'h1f];
  assign T114 = io_fn[2'h3:2'h3];
  assign T115 = io_in1[6'h3f:6'h20];
  assign T116 = io_dw == 1'h1;
  assign T117 = T119 | T118;
  assign T118 = io_fn == 4'hb;
  assign T119 = io_fn == 4'h5;
  assign T120 = T122 & T121;
  assign T121 = shin[6'h3f:6'h3f];
  assign T122 = io_fn[2'h3:2'h3];
  assign T123 = T125 | T124;
  assign T124 = io_fn == 4'hb;
  assign T125 = io_fn == 4'h5;
  assign T126 = T128 | T127;
  assign T127 = io_fn == 4'ha;
  assign T128 = io_fn == 4'h0;
  assign out_hi = T132 ? T131 : T129;
  assign T129 = 32'h0 - T147;
  assign T147 = {31'h0, T130};
  assign T130 = out64[5'h1f:5'h1f];
  assign T131 = out64[6'h3f:6'h20];
  assign T132 = io_dw == 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[129:0] T180;
  wire[63:0] negated_remainder;
  wire[63:0] T119;
  wire T11;
  wire T12;
  reg  isMul;
  wire T13;
  wire cmdMul;
  wire T14;
  wire[3:0] T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  reg [2:0] state;
  wire[2:0] T181;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  reg  neg_out;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  isHi;
  wire T33;
  wire cmdHi;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire T37;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T41;
  wire[64:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[64:0] T46;
  wire[63:0] rhs_in;
  wire[31:0] T47;
  wire[31:0] T48;
  wire[31:0] T49;
  wire[31:0] T182;
  wire[31:0] T50;
  wire T51;
  wire rhs_sign;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire rhsSigned;
  wire T56;
  wire[3:0] T57;
  wire[64:0] T58;
  wire T59;
  reg [6:0] count;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire[6:0] T65;
  wire[6:0] T183;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[5:0] T184;
  wire[5:0] T185;
  wire[5:0] T186;
  wire[5:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[5:0] T190;
  wire[5:0] T191;
  wire[5:0] T192;
  wire[5:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire[5:0] T196;
  wire[5:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[4:0] T216;
  wire[4:0] T217;
  wire[4:0] T218;
  wire[4:0] T219;
  wire[4:0] T220;
  wire[4:0] T221;
  wire[4:0] T222;
  wire[4:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[4:0] T226;
  wire[4:0] T227;
  wire[4:0] T228;
  wire[4:0] T229;
  wire[4:0] T230;
  wire[4:0] T231;
  wire[3:0] T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[3:0] T238;
  wire[3:0] T239;
  wire[2:0] T240;
  wire[2:0] T241;
  wire[2:0] T242;
  wire[2:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire T246;
  wire[63:0] T70;
  wire[63:0] T71;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire[5:0] T72;
  wire[5:0] T309;
  wire[5:0] T310;
  wire[5:0] T311;
  wire[5:0] T312;
  wire[5:0] T313;
  wire[5:0] T314;
  wire[5:0] T315;
  wire[5:0] T316;
  wire[5:0] T317;
  wire[5:0] T318;
  wire[5:0] T319;
  wire[5:0] T320;
  wire[5:0] T321;
  wire[5:0] T322;
  wire[5:0] T323;
  wire[5:0] T324;
  wire[5:0] T325;
  wire[5:0] T326;
  wire[5:0] T327;
  wire[5:0] T328;
  wire[5:0] T329;
  wire[5:0] T330;
  wire[5:0] T331;
  wire[5:0] T332;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[4:0] T341;
  wire[4:0] T342;
  wire[4:0] T343;
  wire[4:0] T344;
  wire[4:0] T345;
  wire[4:0] T346;
  wire[4:0] T347;
  wire[4:0] T348;
  wire[4:0] T349;
  wire[4:0] T350;
  wire[4:0] T351;
  wire[4:0] T352;
  wire[4:0] T353;
  wire[4:0] T354;
  wire[4:0] T355;
  wire[4:0] T356;
  wire[3:0] T357;
  wire[3:0] T358;
  wire[3:0] T359;
  wire[3:0] T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[2:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire T371;
  wire[63:0] T74;
  wire[63:0] T75;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire lhs_sign;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire lhsSigned;
  wire T84;
  wire[3:0] T85;
  wire T86;
  wire T87;
  wire[2:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[64:0] T97;
  wire[5:0] T98;
  wire[10:0] T99;
  wire[63:0] T100;
  wire[128:0] T101;
  wire[63:0] T102;
  wire[64:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire[129:0] T434;
  wire T120;
  wire[129:0] T435;
  wire[63:0] T121;
  wire T122;
  wire[129:0] T123;
  wire[129:0] T124;
  wire[64:0] T125;
  wire[63:0] T126;
  wire[128:0] T127;
  wire[63:0] T128;
  wire[128:0] T129;
  wire[128:0] T130;
  wire[128:0] T131;
  wire[55:0] T132;
  wire[72:0] T133;
  wire[72:0] T436;
  wire[64:0] T134;
  wire[64:0] T135;
  wire[7:0] T437;
  wire T438;
  wire[72:0] T136;
  wire[8:0] T137;
  wire[8:0] T138;
  wire[7:0] T139;
  wire[64:0] T140;
  wire[128:0] T141;
  wire[5:0] T142;
  wire[10:0] T143;
  wire[10:0] T144;
  wire[64:0] T145;
  wire[64:0] T146;
  wire T147;
  wire T148;
  wire[129:0] T439;
  wire[128:0] T149;
  wire[64:0] T150;
  wire T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[63:0] T154;
  wire[63:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[129:0] T440;
  wire[126:0] T159;
  wire[63:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire[129:0] T441;
  wire[63:0] lhs_in;
  wire[31:0] T167;
  wire[31:0] T168;
  wire[31:0] T169;
  wire[31:0] T442;
  wire[31:0] T170;
  wire T171;
  wire[63:0] T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T443;
  wire T175;
  wire T176;
  reg  req_dw;
  wire T177;
  wire T178;
  wire T179;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T176 ? T172 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T441 : T5;
  assign T5 = T161 ? T440 : T6;
  assign T6 = T156 ? T439 : T7;
  assign T7 = T147 ? T123 : T8;
  assign T8 = T122 ? T435 : T9;
  assign T9 = T120 ? T434 : T10;
  assign T10 = T11 ? T180 : remainder;
  assign T180 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T119;
  assign T119 = remainder[6'h3f:1'h0];
  assign T11 = T19 & T12;
  assign T12 = T18 | isMul;
  assign T13 = T1 ? cmdMul : isMul;
  assign cmdMul = T16 | T14;
  assign T14 = T15 == 4'h8;
  assign T15 = io_req_bits_fn & 4'h8;
  assign T16 = T17 == 4'h0;
  assign T17 = io_req_bits_fn & 4'h4;
  assign T18 = remainder[6'h3f:6'h3f];
  assign T19 = state == 3'h1;
  assign T181 = reset ? 3'h0 : T20;
  assign T20 = T1 ? T115 : T21;
  assign T21 = T113 ? 3'h0 : T22;
  assign T22 = T111 ? T109 : T23;
  assign T23 = T89 ? T88 : T24;
  assign T24 = T122 ? T27 : T25;
  assign T25 = T120 ? 3'h5 : T26;
  assign T26 = T19 ? 3'h2 : state;
  assign T27 = neg_out ? 3'h4 : 3'h5;
  assign T28 = T1 ? T77 : T29;
  assign T29 = T30 ? 1'h0 : neg_out;
  assign T30 = T156 & T31;
  assign T31 = T39 & T32;
  assign T32 = isHi ^ 1'h1;
  assign T33 = T1 ? cmdHi : isHi;
  assign cmdHi = T34 | T14;
  assign T34 = T37 | T35;
  assign T35 = T36 == 4'h2;
  assign T36 = io_req_bits_fn & 4'h2;
  assign T37 = T38 == 4'h1;
  assign T38 = io_req_bits_fn & 4'h5;
  assign T39 = T59 & T40;
  assign T40 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T58 - divisor;
  assign T41 = T1 ? T46 : T42;
  assign T42 = T43 ? subtractor : divisor;
  assign T43 = T19 & T44;
  assign T44 = T45 | isMul;
  assign T45 = divisor[6'h3f:6'h3f];
  assign T46 = {rhs_sign, rhs_in};
  assign rhs_in = {T48, T47};
  assign T47 = io_req_bits_in2[5'h1f:1'h0];
  assign T48 = T51 ? T50 : T49;
  assign T49 = 32'h0 - T182;
  assign T182 = {31'h0, rhs_sign};
  assign T50 = io_req_bits_in2[6'h3f:6'h20];
  assign T51 = io_req_bits_dw == 1'h1;
  assign rhs_sign = rhsSigned & T52;
  assign T52 = T55 ? T54 : T53;
  assign T53 = io_req_bits_in2[5'h1f:5'h1f];
  assign T54 = io_req_bits_in2[6'h3f:6'h3f];
  assign T55 = io_req_bits_dw == 1'h1;
  assign rhsSigned = T56 | T16;
  assign T56 = T57 == 4'h0;
  assign T57 = io_req_bits_fn & 4'h9;
  assign T58 = remainder[8'h80:7'h40];
  assign T59 = count == 7'h0;
  assign T60 = T1 ? 7'h0 : T61;
  assign T61 = T161 ? T183 : T62;
  assign T62 = T156 ? T65 : T63;
  assign T63 = T147 ? T64 : count;
  assign T64 = count + 7'h1;
  assign T65 = count + 7'h1;
  assign T183 = {1'h0, T66};
  assign T66 = T76 ? 6'h3f : T67;
  assign T67 = T68[3'h5:1'h0];
  assign T68 = T72 - T184;
  assign T184 = T308 ? 6'h3f : T185;
  assign T185 = T307 ? 6'h3e : T186;
  assign T186 = T306 ? 6'h3d : T187;
  assign T187 = T305 ? 6'h3c : T188;
  assign T188 = T304 ? 6'h3b : T189;
  assign T189 = T303 ? 6'h3a : T190;
  assign T190 = T302 ? 6'h39 : T191;
  assign T191 = T301 ? 6'h38 : T192;
  assign T192 = T300 ? 6'h37 : T193;
  assign T193 = T299 ? 6'h36 : T194;
  assign T194 = T298 ? 6'h35 : T195;
  assign T195 = T297 ? 6'h34 : T196;
  assign T196 = T296 ? 6'h33 : T197;
  assign T197 = T295 ? 6'h32 : T198;
  assign T198 = T294 ? 6'h31 : T199;
  assign T199 = T293 ? 6'h30 : T200;
  assign T200 = T292 ? 6'h2f : T201;
  assign T201 = T291 ? 6'h2e : T202;
  assign T202 = T290 ? 6'h2d : T203;
  assign T203 = T289 ? 6'h2c : T204;
  assign T204 = T288 ? 6'h2b : T205;
  assign T205 = T287 ? 6'h2a : T206;
  assign T206 = T286 ? 6'h29 : T207;
  assign T207 = T285 ? 6'h28 : T208;
  assign T208 = T284 ? 6'h27 : T209;
  assign T209 = T283 ? 6'h26 : T210;
  assign T210 = T282 ? 6'h25 : T211;
  assign T211 = T281 ? 6'h24 : T212;
  assign T212 = T280 ? 6'h23 : T213;
  assign T213 = T279 ? 6'h22 : T214;
  assign T214 = T278 ? 6'h21 : T215;
  assign T215 = T277 ? 6'h20 : T216;
  assign T216 = T276 ? 5'h1f : T217;
  assign T217 = T275 ? 5'h1e : T218;
  assign T218 = T274 ? 5'h1d : T219;
  assign T219 = T273 ? 5'h1c : T220;
  assign T220 = T272 ? 5'h1b : T221;
  assign T221 = T271 ? 5'h1a : T222;
  assign T222 = T270 ? 5'h19 : T223;
  assign T223 = T269 ? 5'h18 : T224;
  assign T224 = T268 ? 5'h17 : T225;
  assign T225 = T267 ? 5'h16 : T226;
  assign T226 = T266 ? 5'h15 : T227;
  assign T227 = T265 ? 5'h14 : T228;
  assign T228 = T264 ? 5'h13 : T229;
  assign T229 = T263 ? 5'h12 : T230;
  assign T230 = T262 ? 5'h11 : T231;
  assign T231 = T261 ? 5'h10 : T232;
  assign T232 = T260 ? 4'hf : T233;
  assign T233 = T259 ? 4'he : T234;
  assign T234 = T258 ? 4'hd : T235;
  assign T235 = T257 ? 4'hc : T236;
  assign T236 = T256 ? 4'hb : T237;
  assign T237 = T255 ? 4'ha : T238;
  assign T238 = T254 ? 4'h9 : T239;
  assign T239 = T253 ? 4'h8 : T240;
  assign T240 = T252 ? 3'h7 : T241;
  assign T241 = T251 ? 3'h6 : T242;
  assign T242 = T250 ? 3'h5 : T243;
  assign T243 = T249 ? 3'h4 : T244;
  assign T244 = T248 ? 2'h3 : T245;
  assign T245 = T247 ? 2'h2 : T246;
  assign T246 = T70[1'h1:1'h1];
  assign T70 = T71[6'h3f:1'h0];
  assign T71 = remainder[6'h3f:1'h0];
  assign T247 = T70[2'h2:2'h2];
  assign T248 = T70[2'h3:2'h3];
  assign T249 = T70[3'h4:3'h4];
  assign T250 = T70[3'h5:3'h5];
  assign T251 = T70[3'h6:3'h6];
  assign T252 = T70[3'h7:3'h7];
  assign T253 = T70[4'h8:4'h8];
  assign T254 = T70[4'h9:4'h9];
  assign T255 = T70[4'ha:4'ha];
  assign T256 = T70[4'hb:4'hb];
  assign T257 = T70[4'hc:4'hc];
  assign T258 = T70[4'hd:4'hd];
  assign T259 = T70[4'he:4'he];
  assign T260 = T70[4'hf:4'hf];
  assign T261 = T70[5'h10:5'h10];
  assign T262 = T70[5'h11:5'h11];
  assign T263 = T70[5'h12:5'h12];
  assign T264 = T70[5'h13:5'h13];
  assign T265 = T70[5'h14:5'h14];
  assign T266 = T70[5'h15:5'h15];
  assign T267 = T70[5'h16:5'h16];
  assign T268 = T70[5'h17:5'h17];
  assign T269 = T70[5'h18:5'h18];
  assign T270 = T70[5'h19:5'h19];
  assign T271 = T70[5'h1a:5'h1a];
  assign T272 = T70[5'h1b:5'h1b];
  assign T273 = T70[5'h1c:5'h1c];
  assign T274 = T70[5'h1d:5'h1d];
  assign T275 = T70[5'h1e:5'h1e];
  assign T276 = T70[5'h1f:5'h1f];
  assign T277 = T70[6'h20:6'h20];
  assign T278 = T70[6'h21:6'h21];
  assign T279 = T70[6'h22:6'h22];
  assign T280 = T70[6'h23:6'h23];
  assign T281 = T70[6'h24:6'h24];
  assign T282 = T70[6'h25:6'h25];
  assign T283 = T70[6'h26:6'h26];
  assign T284 = T70[6'h27:6'h27];
  assign T285 = T70[6'h28:6'h28];
  assign T286 = T70[6'h29:6'h29];
  assign T287 = T70[6'h2a:6'h2a];
  assign T288 = T70[6'h2b:6'h2b];
  assign T289 = T70[6'h2c:6'h2c];
  assign T290 = T70[6'h2d:6'h2d];
  assign T291 = T70[6'h2e:6'h2e];
  assign T292 = T70[6'h2f:6'h2f];
  assign T293 = T70[6'h30:6'h30];
  assign T294 = T70[6'h31:6'h31];
  assign T295 = T70[6'h32:6'h32];
  assign T296 = T70[6'h33:6'h33];
  assign T297 = T70[6'h34:6'h34];
  assign T298 = T70[6'h35:6'h35];
  assign T299 = T70[6'h36:6'h36];
  assign T300 = T70[6'h37:6'h37];
  assign T301 = T70[6'h38:6'h38];
  assign T302 = T70[6'h39:6'h39];
  assign T303 = T70[6'h3a:6'h3a];
  assign T304 = T70[6'h3b:6'h3b];
  assign T305 = T70[6'h3c:6'h3c];
  assign T306 = T70[6'h3d:6'h3d];
  assign T307 = T70[6'h3e:6'h3e];
  assign T308 = T70[6'h3f:6'h3f];
  assign T72 = 6'h3f + T309;
  assign T309 = T433 ? 6'h3f : T310;
  assign T310 = T432 ? 6'h3e : T311;
  assign T311 = T431 ? 6'h3d : T312;
  assign T312 = T430 ? 6'h3c : T313;
  assign T313 = T429 ? 6'h3b : T314;
  assign T314 = T428 ? 6'h3a : T315;
  assign T315 = T427 ? 6'h39 : T316;
  assign T316 = T426 ? 6'h38 : T317;
  assign T317 = T425 ? 6'h37 : T318;
  assign T318 = T424 ? 6'h36 : T319;
  assign T319 = T423 ? 6'h35 : T320;
  assign T320 = T422 ? 6'h34 : T321;
  assign T321 = T421 ? 6'h33 : T322;
  assign T322 = T420 ? 6'h32 : T323;
  assign T323 = T419 ? 6'h31 : T324;
  assign T324 = T418 ? 6'h30 : T325;
  assign T325 = T417 ? 6'h2f : T326;
  assign T326 = T416 ? 6'h2e : T327;
  assign T327 = T415 ? 6'h2d : T328;
  assign T328 = T414 ? 6'h2c : T329;
  assign T329 = T413 ? 6'h2b : T330;
  assign T330 = T412 ? 6'h2a : T331;
  assign T331 = T411 ? 6'h29 : T332;
  assign T332 = T410 ? 6'h28 : T333;
  assign T333 = T409 ? 6'h27 : T334;
  assign T334 = T408 ? 6'h26 : T335;
  assign T335 = T407 ? 6'h25 : T336;
  assign T336 = T406 ? 6'h24 : T337;
  assign T337 = T405 ? 6'h23 : T338;
  assign T338 = T404 ? 6'h22 : T339;
  assign T339 = T403 ? 6'h21 : T340;
  assign T340 = T402 ? 6'h20 : T341;
  assign T341 = T401 ? 5'h1f : T342;
  assign T342 = T400 ? 5'h1e : T343;
  assign T343 = T399 ? 5'h1d : T344;
  assign T344 = T398 ? 5'h1c : T345;
  assign T345 = T397 ? 5'h1b : T346;
  assign T346 = T396 ? 5'h1a : T347;
  assign T347 = T395 ? 5'h19 : T348;
  assign T348 = T394 ? 5'h18 : T349;
  assign T349 = T393 ? 5'h17 : T350;
  assign T350 = T392 ? 5'h16 : T351;
  assign T351 = T391 ? 5'h15 : T352;
  assign T352 = T390 ? 5'h14 : T353;
  assign T353 = T389 ? 5'h13 : T354;
  assign T354 = T388 ? 5'h12 : T355;
  assign T355 = T387 ? 5'h11 : T356;
  assign T356 = T386 ? 5'h10 : T357;
  assign T357 = T385 ? 4'hf : T358;
  assign T358 = T384 ? 4'he : T359;
  assign T359 = T383 ? 4'hd : T360;
  assign T360 = T382 ? 4'hc : T361;
  assign T361 = T381 ? 4'hb : T362;
  assign T362 = T380 ? 4'ha : T363;
  assign T363 = T379 ? 4'h9 : T364;
  assign T364 = T378 ? 4'h8 : T365;
  assign T365 = T377 ? 3'h7 : T366;
  assign T366 = T376 ? 3'h6 : T367;
  assign T367 = T375 ? 3'h5 : T368;
  assign T368 = T374 ? 3'h4 : T369;
  assign T369 = T373 ? 2'h3 : T370;
  assign T370 = T372 ? 2'h2 : T371;
  assign T371 = T74[1'h1:1'h1];
  assign T74 = T75[6'h3f:1'h0];
  assign T75 = divisor[6'h3f:1'h0];
  assign T372 = T74[2'h2:2'h2];
  assign T373 = T74[2'h3:2'h3];
  assign T374 = T74[3'h4:3'h4];
  assign T375 = T74[3'h5:3'h5];
  assign T376 = T74[3'h6:3'h6];
  assign T377 = T74[3'h7:3'h7];
  assign T378 = T74[4'h8:4'h8];
  assign T379 = T74[4'h9:4'h9];
  assign T380 = T74[4'ha:4'ha];
  assign T381 = T74[4'hb:4'hb];
  assign T382 = T74[4'hc:4'hc];
  assign T383 = T74[4'hd:4'hd];
  assign T384 = T74[4'he:4'he];
  assign T385 = T74[4'hf:4'hf];
  assign T386 = T74[5'h10:5'h10];
  assign T387 = T74[5'h11:5'h11];
  assign T388 = T74[5'h12:5'h12];
  assign T389 = T74[5'h13:5'h13];
  assign T390 = T74[5'h14:5'h14];
  assign T391 = T74[5'h15:5'h15];
  assign T392 = T74[5'h16:5'h16];
  assign T393 = T74[5'h17:5'h17];
  assign T394 = T74[5'h18:5'h18];
  assign T395 = T74[5'h19:5'h19];
  assign T396 = T74[5'h1a:5'h1a];
  assign T397 = T74[5'h1b:5'h1b];
  assign T398 = T74[5'h1c:5'h1c];
  assign T399 = T74[5'h1d:5'h1d];
  assign T400 = T74[5'h1e:5'h1e];
  assign T401 = T74[5'h1f:5'h1f];
  assign T402 = T74[6'h20:6'h20];
  assign T403 = T74[6'h21:6'h21];
  assign T404 = T74[6'h22:6'h22];
  assign T405 = T74[6'h23:6'h23];
  assign T406 = T74[6'h24:6'h24];
  assign T407 = T74[6'h25:6'h25];
  assign T408 = T74[6'h26:6'h26];
  assign T409 = T74[6'h27:6'h27];
  assign T410 = T74[6'h28:6'h28];
  assign T411 = T74[6'h29:6'h29];
  assign T412 = T74[6'h2a:6'h2a];
  assign T413 = T74[6'h2b:6'h2b];
  assign T414 = T74[6'h2c:6'h2c];
  assign T415 = T74[6'h2d:6'h2d];
  assign T416 = T74[6'h2e:6'h2e];
  assign T417 = T74[6'h2f:6'h2f];
  assign T418 = T74[6'h30:6'h30];
  assign T419 = T74[6'h31:6'h31];
  assign T420 = T74[6'h32:6'h32];
  assign T421 = T74[6'h33:6'h33];
  assign T422 = T74[6'h34:6'h34];
  assign T423 = T74[6'h35:6'h35];
  assign T424 = T74[6'h36:6'h36];
  assign T425 = T74[6'h37:6'h37];
  assign T426 = T74[6'h38:6'h38];
  assign T427 = T74[6'h39:6'h39];
  assign T428 = T74[6'h3a:6'h3a];
  assign T429 = T74[6'h3b:6'h3b];
  assign T430 = T74[6'h3c:6'h3c];
  assign T431 = T74[6'h3d:6'h3d];
  assign T432 = T74[6'h3e:6'h3e];
  assign T433 = T74[6'h3f:6'h3f];
  assign T76 = T184 < T309;
  assign T77 = T87 & T78;
  assign T78 = cmdHi ? lhs_sign : T79;
  assign T79 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T80;
  assign T80 = T83 ? T82 : T81;
  assign T81 = io_req_bits_in1[5'h1f:5'h1f];
  assign T82 = io_req_bits_in1[6'h3f:6'h3f];
  assign T83 = io_req_bits_dw == 1'h1;
  assign lhsSigned = T86 | T84;
  assign T84 = T85 == 4'h0;
  assign T85 = io_req_bits_fn & 4'h3;
  assign T86 = T56 | T16;
  assign T87 = cmdMul ^ 1'h1;
  assign T88 = isHi ? 3'h3 : 3'h5;
  assign T89 = T147 & T90;
  assign T90 = T92 | T91;
  assign T91 = count == 7'h7;
  assign T92 = T104 & T93;
  assign T93 = T94 == 64'h0;
  assign T94 = T100 & T95;
  assign T95 = ~ T96;
  assign T96 = T97[6'h3f:1'h0];
  assign T97 = $signed(65'h10000000000000000) >>> T98;
  assign T98 = T99[3'h5:1'h0];
  assign T99 = count * 4'h8;
  assign T100 = T101[6'h3f:1'h0];
  assign T101 = {T103, T102};
  assign T102 = remainder[6'h3f:1'h0];
  assign T103 = remainder[8'h81:7'h41];
  assign T104 = T106 & T105;
  assign T105 = isHi ^ 1'h1;
  assign T106 = T108 & T107;
  assign T107 = count != 7'h0;
  assign T108 = count != 7'h7;
  assign T109 = isHi ? 3'h3 : T110;
  assign T110 = neg_out ? 3'h4 : 3'h5;
  assign T111 = T156 & T112;
  assign T112 = count == 7'h40;
  assign T113 = T114 | io_kill;
  assign T114 = io_resp_ready & io_resp_valid;
  assign T115 = T116 ? 3'h1 : 3'h2;
  assign T116 = lhs_sign | T117;
  assign T117 = rhs_sign & T118;
  assign T118 = cmdMul ^ 1'h1;
  assign T434 = {66'h0, negated_remainder};
  assign T120 = state == 3'h4;
  assign T435 = {66'h0, T121};
  assign T121 = remainder[8'h80:7'h41];
  assign T122 = state == 3'h3;
  assign T123 = T124;
  assign T124 = {T146, T125};
  assign T125 = {1'h0, T126};
  assign T126 = T127[6'h3f:1'h0];
  assign T127 = {T145, T128};
  assign T128 = T129[6'h3f:1'h0];
  assign T129 = T92 ? T141 : T130;
  assign T130 = T131;
  assign T131 = {T133, T132};
  assign T132 = T100[6'h3f:4'h8];
  assign T133 = T136 + T436;
  assign T436 = {T437, T134};
  assign T134 = T135;
  assign T135 = T101[8'h80:7'h40];
  assign T437 = T438 ? 8'hff : 8'h0;
  assign T438 = T134[7'h40:7'h40];
  assign T136 = $signed(T140) * $signed(T137);
  assign T137 = T138;
  assign T138 = {1'h0, T139};
  assign T139 = T100[3'h7:1'h0];
  assign T140 = divisor;
  assign T141 = T101 >> T142;
  assign T142 = T143[3'h5:1'h0];
  assign T143 = 11'h40 - T144;
  assign T144 = count * 4'h8;
  assign T145 = T130[8'h80:7'h40];
  assign T146 = T127 >> 7'h40;
  assign T147 = T148 & isMul;
  assign T148 = state == 3'h2;
  assign T439 = {1'h0, T149};
  assign T149 = {T153, T150};
  assign T150 = {T152, T151};
  assign T151 = less ^ 1'h1;
  assign T152 = remainder[6'h3f:1'h0];
  assign T153 = less ? T155 : T154;
  assign T154 = subtractor[6'h3f:1'h0];
  assign T155 = remainder[7'h7f:7'h40];
  assign T156 = T158 & T157;
  assign T157 = isMul ^ 1'h1;
  assign T158 = state == 3'h2;
  assign T440 = {3'h0, T159};
  assign T159 = T160 << T66;
  assign T160 = remainder[6'h3f:1'h0];
  assign T161 = T156 & T162;
  assign T162 = T165 & T163;
  assign T163 = T164 | T76;
  assign T164 = 6'h0 < T68;
  assign T165 = T166 & less;
  assign T166 = count == 7'h0;
  assign T441 = {66'h0, lhs_in};
  assign lhs_in = {T168, T167};
  assign T167 = io_req_bits_in1[5'h1f:1'h0];
  assign T168 = T171 ? T170 : T169;
  assign T169 = 32'h0 - T442;
  assign T442 = {31'h0, lhs_sign};
  assign T170 = io_req_bits_in1[6'h3f:6'h20];
  assign T171 = io_req_bits_dw == 1'h1;
  assign T172 = {T174, T173};
  assign T173 = remainder[5'h1f:1'h0];
  assign T174 = 32'h0 - T443;
  assign T443 = {31'h0, T175};
  assign T175 = remainder[5'h1f:5'h1f];
  assign T176 = req_dw == 1'h0;
  assign T177 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T178;
  assign T178 = state == 3'h5;
  assign io_req_ready = T179;
  assign T179 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T441;
    end else if(T161) begin
      remainder <= T440;
    end else if(T156) begin
      remainder <= T439;
    end else if(T147) begin
      remainder <= T123;
    end else if(T122) begin
      remainder <= T435;
    end else if(T120) begin
      remainder <= T434;
    end else if(T11) begin
      remainder <= T180;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T115;
    end else if(T113) begin
      state <= 3'h0;
    end else if(T111) begin
      state <= T109;
    end else if(T89) begin
      state <= T88;
    end else if(T122) begin
      state <= T27;
    end else if(T120) begin
      state <= 3'h5;
    end else if(T19) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T77;
    end else if(T30) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T46;
    end else if(T43) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T161) begin
      count <= T183;
    end else if(T156) begin
      count <= T65;
    end else if(T147) begin
      count <= T64;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module ManagementMachine(input clk, input reset,
    output io_stall_out,
    input  io_write_to_cfga,
    input [63:0] io_cfgd_in,
    output io_s_axi_awvalid,
    input  io_s_axi_awready,
    output io_s_axi_wvalid,
    input  io_s_axi_wready,
    input [1:0] io_s_axi_bresp,
    input  io_s_axi_bvalid,
    output io_s_axi_bready,
    output io_s_axi_arvalid,
    input  io_s_axi_arready,
    input [31:0] io_s_axi_rdata,
    input [1:0] io_s_axi_rresp,
    input  io_s_axi_rvalid,
    output io_s_axi_rready,
    output io_sfp_tx_disable
);

  wire T0;
  reg [31:0] bringup_sfp_tx_disable;
  wire[31:0] T66;
  wire[31:0] T1;
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  reg [2:0] state;
  wire[2:0] T67;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  reg  handled;
  wire T68;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    bringup_sfp_tx_disable = {1{$random}};
    state = {1{$random}};
    handled = {1{$random}};
  end
`endif

  assign io_sfp_tx_disable = T0;
  assign T0 = bringup_sfp_tx_disable < 32'h2faf080;
  assign T66 = reset ? 32'h0 : T1;
  assign T1 = T9 ? 32'h1 : T2;
  assign T2 = T6 ? 32'h0 : T3;
  assign T3 = T5 ? bringup_sfp_tx_disable : T4;
  assign T4 = bringup_sfp_tx_disable + 32'h1;
  assign T5 = bringup_sfp_tx_disable == 32'h0;
  assign T6 = T8 & T7;
  assign T7 = bringup_sfp_tx_disable == 32'h5f5e100;
  assign T8 = T5 ^ 1'h1;
  assign T9 = T11 & T10;
  assign T10 = io_cfgd_in[6'h21:6'h21];
  assign T11 = T12 & io_s_axi_bvalid;
  assign T12 = T48 & T13;
  assign T13 = state == 3'h4;
  assign T67 = reset ? 3'h0 : T14;
  assign T14 = T45 ? 3'h0 : T15;
  assign T15 = T11 ? 3'h0 : T16;
  assign T16 = T40 ? 3'h0 : T17;
  assign T17 = T35 ? 3'h4 : T18;
  assign T18 = T29 ? 3'h3 : T19;
  assign T19 = T23 ? 3'h2 : T20;
  assign T20 = T21 ? 3'h1 : state;
  assign T21 = T22 & io_write_to_cfga;
  assign T22 = state == 3'h0;
  assign T23 = T26 & T24;
  assign T24 = T25 & io_s_axi_awready;
  assign T25 = io_cfgd_in[6'h20:6'h20];
  assign T26 = T28 & T27;
  assign T27 = state == 3'h1;
  assign T28 = T22 ^ 1'h1;
  assign T29 = T26 & T30;
  assign T30 = T34 & T31;
  assign T31 = T32 & io_s_axi_arready;
  assign T32 = T33 == 1'h0;
  assign T33 = io_cfgd_in[6'h20:6'h20];
  assign T34 = T24 ^ 1'h1;
  assign T35 = T36 & io_s_axi_wready;
  assign T36 = T38 & T37;
  assign T37 = state == 3'h2;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T22 | T27;
  assign T40 = T41 & io_s_axi_rvalid;
  assign T41 = T43 & T42;
  assign T42 = state == 3'h3;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T39 | T37;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 | T13;
  assign T47 = T44 | T42;
  assign T48 = T47 ^ 1'h1;
  assign io_s_axi_rready = T49;
  assign T49 = state == 3'h3;
  assign io_s_axi_arvalid = T50;
  assign T50 = T53 & T51;
  assign T51 = T52 == 1'h0;
  assign T52 = io_cfgd_in[6'h20:6'h20];
  assign T53 = state == 3'h1;
  assign io_s_axi_bready = T54;
  assign T54 = state == 3'h4;
  assign io_s_axi_wvalid = T55;
  assign T55 = state == 3'h2;
  assign io_s_axi_awvalid = T56;
  assign T56 = T58 & T57;
  assign T57 = io_cfgd_in[6'h20:6'h20];
  assign T58 = state == 3'h1;
  assign io_stall_out = T59;
  assign T59 = T64 & T60;
  assign T60 = handled == 1'h0;
  assign T68 = reset ? 1'h0 : T61;
  assign T61 = T11 ? 1'h1 : T62;
  assign T62 = T40 ? 1'h1 : T63;
  assign T63 = T22 ? 1'h0 : handled;
  assign T64 = T65 | io_write_to_cfga;
  assign T65 = state != 3'h0;

  always @(posedge clk) begin
    if(reset) begin
      bringup_sfp_tx_disable <= 32'h0;
    end else if(T9) begin
      bringup_sfp_tx_disable <= 32'h1;
    end else if(T6) begin
      bringup_sfp_tx_disable <= 32'h0;
    end else if(T5) begin
      bringup_sfp_tx_disable <= bringup_sfp_tx_disable;
    end else begin
      bringup_sfp_tx_disable <= T4;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T45) begin
      state <= 3'h0;
    end else if(T11) begin
      state <= 3'h0;
    end else if(T40) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h4;
    end else if(T29) begin
      state <= 3'h3;
    end else if(T23) begin
      state <= 3'h2;
    end else if(T21) begin
      state <= 3'h1;
    end
    if(reset) begin
      handled <= 1'h0;
    end else if(T11) begin
      handled <= 1'h1;
    end else if(T40) begin
      handled <= 1'h1;
    end else if(T22) begin
      handled <= 1'h0;
    end
  end
endmodule

module TransmitMachine(input clk, input reset,
    output[7:0] io_tx_axis_fifo_tdata,
    output io_tx_axis_fifo_tvalid,
    input  io_tx_axis_fifo_tready,
    output io_tx_axis_fifo_tlast,
    input [63:0] io_txd_in,
    input  io_write_to_txd
);

  wire T0;
  wire T1;
  reg  state;
  wire T11;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[7:0] T10;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
  end
`endif

  assign io_tx_axis_fifo_tlast = T0;
  assign T0 = io_txd_in[4'h9:4'h9];
  assign io_tx_axis_fifo_tvalid = T1;
  assign T1 = state == 1'h1;
  assign T11 = reset ? 1'h0 : T2;
  assign T2 = T6 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : state;
  assign T4 = T5 & io_write_to_txd;
  assign T5 = state == 1'h0;
  assign T6 = T7 & io_tx_axis_fifo_tready;
  assign T7 = T9 & T8;
  assign T8 = state == 1'h1;
  assign T9 = T5 ^ 1'h1;
  assign io_tx_axis_fifo_tdata = T10;
  assign T10 = io_txd_in[3'h7:1'h0];

  always @(posedge clk) begin
    if(reset) begin
      state <= 1'h0;
    end else if(T6) begin
      state <= 1'h0;
    end else if(T4) begin
      state <= 1'h1;
    end
  end
endmodule

module ReceiveMachine(input clk, input reset,
    input [7:0] io_rx_axis_fifo_tdata,
    input  io_rx_axis_fifo_tvalid,
    output io_rx_axis_fifo_tready,
    input  io_rx_axis_fifo_tlast,
    output[63:0] io_rxd_val,
    input [63:0] io_rxd_val_in,
    input  io_rxd_val_in_valid
);

  reg [63:0] rxd_reg;
  wire[63:0] T11;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T12;
  wire[9:0] T2;
  wire[8:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    rxd_reg = {2{$random}};
  end
`endif

  assign io_rxd_val = rxd_reg;
  assign T11 = reset ? 64'h0 : T0;
  assign T0 = T4 ? T12 : T1;
  assign T1 = io_rxd_val_in_valid ? io_rxd_val_in : rxd_reg;
  assign T12 = {54'h0, T2};
  assign T2 = {io_rx_axis_fifo_tlast, T3};
  assign T3 = {1'h1, io_rx_axis_fifo_tdata};
  assign T4 = T8 & T5;
  assign T5 = T6 & io_rx_axis_fifo_tvalid;
  assign T6 = T7 == 1'h0;
  assign T7 = rxd_reg[4'h8:4'h8];
  assign T8 = io_rxd_val_in_valid ^ 1'h1;
  assign io_rx_axis_fifo_tready = T9;
  assign T9 = T10 == 1'h0;
  assign T10 = rxd_reg[4'h8:4'h8];

  always @(posedge clk) begin
    if(reset) begin
      rxd_reg <= 64'h0;
    end else if(T4) begin
      rxd_reg <= T12;
    end else if(io_rxd_val_in_valid) begin
      rxd_reg <= io_rxd_val_in;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [1:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready,
    output io_temac_sfp_tx_disable,
    output[7:0] io_status_ip,
    output[7:0] io_status_im,
    output[6:0] io_status_zero,
    output io_status_er,
    output io_status_vm,
    output io_status_s64,
    output io_status_u64,
    output io_status_ef,
    output io_status_pei,
    output io_status_ei,
    output io_status_ps,
    output io_status_s,
    output[31:0] io_ptbr,
    output[43:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input  io_badvaddr_wen,
    input [43:0] io_pc,
    input  io_sret,
    output io_fatc,
    output io_replay,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [2:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [511:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[2:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  wire T593;
  wire T367;
  reg [45:0] T10;
  wire[11:0] addr;
  wire[11:0] T504;
  wire[10:0] T12;
  wire[10:0] T505;
  reg [4:0] host_pcr_bits_addr;
  wire[4:0] T13;
  wire T4;
  wire cpu_req_valid;
  wire wen;
  wire T14;
  reg  host_pcr_bits_rw;
  wire T15;
  wire host_pcr_req_fire;
  wire T5;
  reg  host_pcr_req_valid;
  wire T6;
  wire T7;
  wire[63:0] T594;
  wire[63:0] wdata;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T2;
  wire[63:0] T3;
  wire T371;
  wire T372;
  reg [63:0] reg_txd;
  wire[63:0] T567;
  wire[63:0] T370;
  reg [63:0] reg_cfgd;
  wire[63:0] T517;
  wire[63:0] T136;
  wire[63:0] T137;
  wire[63:0] T518;
  wire T138;
  wire T139;
  wire T133;
  wire T134;
  reg [2:0] reg_frm;
  wire[2:0] T502;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T503;
  wire T8;
  wire T9;
  wire[63:0] T506;
  wire[58:0] T16;
  wire T17;
  wire T18;
  wire[63:0] T19;
  reg [5:0] R20;
  wire[5:0] T507;
  wire[5:0] T21;
  wire[5:0] T22;
  wire[6:0] T23;
  wire[6:0] T508;
  wire[5:0] T24;
  wire[63:0] T25;
  wire T26;
  wire T27;
  reg [57:0] R28;
  wire[57:0] T509;
  wire[57:0] T29;
  wire[57:0] T30;
  wire[57:0] T31;
  wire T32;
  wire[57:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[43:0] T38;
  wire[43:0] T39;
  reg [43:0] reg_epc;
  wire[43:0] T40;
  wire[43:0] T41;
  wire[43:0] T42;
  wire[43:0] T43;
  wire[43:0] T44;
  wire T45;
  wire T46;
  wire[43:0] T510;
  wire[42:0] T47;
  reg [42:0] reg_evec;
  wire[42:0] T48;
  wire[42:0] T49;
  wire[42:0] T50;
  wire T51;
  wire T52;
  wire T511;
  reg [31:0] reg_ptbr;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[18:0] T56;
  wire T57;
  wire T58;
  reg  reg_status_s;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  reg_status_ps;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg  reg_status_ei;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  reg_status_pei;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg  reg_status_ef;
  wire T79;
  wire T80;
  wire T81;
  reg  reg_status_u64;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  reg  reg_status_s64;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  reg_status_vm;
  wire T90;
  wire T91;
  wire T92;
  reg  reg_status_er;
  wire T93;
  wire T94;
  wire T95;
  reg [6:0] reg_status_zero;
  wire[6:0] T96;
  wire[6:0] T97;
  wire[6:0] T98;
  wire[6:0] T99;
  reg [7:0] reg_status_im;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[3:0] T104;
  wire[1:0] T105;
  wire[3:0] T106;
  wire[1:0] T107;
  reg  r_rx_axis_fifo_tvalid;
  wire T512;
  reg  r_irq_ipi;
  wire T513;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[1:0] T113;
  wire T114;
  reg [63:0] reg_fromhost;
  wire[63:0] T514;
  wire[63:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  reg  r_irq_timer;
  wire T515;
  wire T122;
  wire T123;
  wire T124;
  reg [31:0] reg_compare;
  wire[31:0] T125;
  wire[31:0] T126;
  wire[31:0] T127;
  wire[31:0] T128;
  wire T129;
  wire T130;
  wire[11:0] T131;
  reg [63:0] reg_cfga;
  wire[63:0] T516;
  wire[63:0] T132;
  wire[31:0] T135;
  wire[11:0] T140;
  wire[63:0] T141;
  wire[63:0] T142;
  wire[63:0] T143;
  reg [5:0] R144;
  wire[5:0] T519;
  wire[5:0] T145;
  wire[5:0] T146;
  wire[6:0] T147;
  wire[6:0] T520;
  wire T148;
  reg [57:0] R149;
  wire[57:0] T521;
  wire[57:0] T150;
  wire[57:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire[63:0] T155;
  wire[63:0] T156;
  wire[63:0] T157;
  reg [5:0] R158;
  wire[5:0] T522;
  wire[5:0] T159;
  wire[5:0] T160;
  wire[6:0] T161;
  wire[6:0] T523;
  wire T162;
  reg [57:0] R163;
  wire[57:0] T524;
  wire[57:0] T164;
  wire[57:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[63:0] T169;
  wire[63:0] T170;
  wire[63:0] T171;
  reg [5:0] R172;
  wire[5:0] T525;
  wire[5:0] T173;
  wire[5:0] T174;
  wire[6:0] T175;
  wire[6:0] T526;
  wire T176;
  reg [57:0] R177;
  wire[57:0] T527;
  wire[57:0] T178;
  wire[57:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[63:0] T183;
  wire[63:0] T184;
  wire[63:0] T185;
  reg [5:0] R186;
  wire[5:0] T528;
  wire[5:0] T187;
  wire[5:0] T188;
  wire[6:0] T189;
  wire[6:0] T529;
  wire T190;
  reg [57:0] R191;
  wire[57:0] T530;
  wire[57:0] T192;
  wire[57:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T199;
  reg [5:0] R200;
  wire[5:0] T531;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[6:0] T203;
  wire[6:0] T532;
  wire T204;
  reg [57:0] R205;
  wire[57:0] T533;
  wire[57:0] T206;
  wire[57:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[63:0] T211;
  wire[63:0] T212;
  wire[63:0] T213;
  reg [5:0] R214;
  wire[5:0] T534;
  wire[5:0] T215;
  wire[5:0] T216;
  wire[6:0] T217;
  wire[6:0] T535;
  wire T218;
  reg [57:0] R219;
  wire[57:0] T536;
  wire[57:0] T220;
  wire[57:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire[63:0] T225;
  wire[63:0] T226;
  wire[63:0] T227;
  reg [5:0] R228;
  wire[5:0] T537;
  wire[5:0] T229;
  wire[5:0] T230;
  wire[6:0] T231;
  wire[6:0] T538;
  wire T232;
  reg [57:0] R233;
  wire[57:0] T539;
  wire[57:0] T234;
  wire[57:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire[63:0] T239;
  wire[63:0] T240;
  wire[63:0] T241;
  reg [5:0] R242;
  wire[5:0] T540;
  wire[5:0] T243;
  wire[5:0] T244;
  wire[6:0] T245;
  wire[6:0] T541;
  wire T246;
  reg [57:0] R247;
  wire[57:0] T542;
  wire[57:0] T248;
  wire[57:0] T249;
  wire T250;
  wire T251;
  wire T252;
  wire[63:0] T253;
  wire[63:0] T254;
  wire[63:0] T255;
  reg [5:0] R256;
  wire[5:0] T543;
  wire[5:0] T257;
  wire[5:0] T258;
  wire[6:0] T259;
  wire[6:0] T544;
  wire T260;
  reg [57:0] R261;
  wire[57:0] T545;
  wire[57:0] T262;
  wire[57:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[63:0] T267;
  wire[63:0] T268;
  wire[63:0] T269;
  reg [5:0] R270;
  wire[5:0] T546;
  wire[5:0] T271;
  wire[5:0] T272;
  wire[6:0] T273;
  wire[6:0] T547;
  wire T274;
  reg [57:0] R275;
  wire[57:0] T548;
  wire[57:0] T276;
  wire[57:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[63:0] T281;
  wire[63:0] T282;
  wire[63:0] T283;
  reg [5:0] R284;
  wire[5:0] T549;
  wire[5:0] T285;
  wire[5:0] T286;
  wire[6:0] T287;
  wire[6:0] T550;
  wire T288;
  reg [57:0] R289;
  wire[57:0] T551;
  wire[57:0] T290;
  wire[57:0] T291;
  wire T292;
  wire T293;
  wire T294;
  wire[63:0] T295;
  wire[63:0] T296;
  wire[63:0] T297;
  reg [5:0] R298;
  wire[5:0] T552;
  wire[5:0] T299;
  wire[5:0] T300;
  wire[6:0] T301;
  wire[6:0] T553;
  wire T302;
  reg [57:0] R303;
  wire[57:0] T554;
  wire[57:0] T304;
  wire[57:0] T305;
  wire T306;
  wire T307;
  wire T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[63:0] T311;
  reg [5:0] R312;
  wire[5:0] T555;
  wire[5:0] T313;
  wire[5:0] T314;
  wire[6:0] T315;
  wire[6:0] T556;
  wire T316;
  reg [57:0] R317;
  wire[57:0] T557;
  wire[57:0] T318;
  wire[57:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[63:0] T323;
  wire[63:0] T324;
  wire[63:0] T325;
  reg [5:0] R326;
  wire[5:0] T558;
  wire[5:0] T327;
  wire[5:0] T328;
  wire[6:0] T329;
  wire[6:0] T559;
  wire T330;
  reg [57:0] R331;
  wire[57:0] T560;
  wire[57:0] T332;
  wire[57:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[63:0] T337;
  wire[63:0] T338;
  wire[63:0] T339;
  reg [5:0] R340;
  wire[5:0] T561;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[6:0] T343;
  wire[6:0] T562;
  wire T344;
  reg [57:0] R345;
  wire[57:0] T563;
  wire[57:0] T346;
  wire[57:0] T347;
  wire T348;
  wire T349;
  wire T350;
  wire[63:0] T351;
  wire[63:0] T352;
  wire[63:0] T353;
  reg [5:0] R354;
  wire[5:0] T564;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[6:0] T357;
  wire[6:0] T565;
  wire T358;
  reg [57:0] R359;
  wire[57:0] T566;
  wire[57:0] T360;
  wire[57:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire[63:0] T365;
  wire[63:0] T366;
  wire[63:0] T368;
  wire[63:0] T369;
  wire[63:0] T373;
  wire[63:0] T374;
  wire[63:0] T375;
  wire[63:0] T376;
  wire[63:0] T377;
  wire[63:0] T378;
  wire[63:0] T379;
  wire[63:0] T380;
  reg [63:0] reg_tohost;
  wire[63:0] T568;
  wire[63:0] T381;
  wire[63:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire[63:0] T391;
  wire[63:0] T569;
  wire T392;
  reg  reg_stats;
  wire T570;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire[63:0] T397;
  wire[63:0] T571;
  wire[1:0] T398;
  wire[63:0] T399;
  wire[63:0] T572;
  wire[1:0] T400;
  wire T401;
  wire[63:0] T402;
  wire[63:0] T573;
  wire[1:0] T403;
  wire[63:0] T404;
  wire[63:0] T574;
  wire[1:0] T405;
  wire T406;
  wire[63:0] T407;
  wire[63:0] T575;
  wire T408;
  wire T409;
  wire[63:0] T410;
  wire[63:0] T576;
  wire[31:0] T411;
  wire[31:0] T412;
  wire[31:0] T413;
  wire[5:0] T414;
  wire[2:0] T415;
  wire[1:0] T416;
  wire[2:0] T417;
  wire[1:0] T418;
  wire[25:0] T419;
  wire[2:0] T420;
  wire[1:0] T421;
  wire[22:0] T422;
  wire[14:0] T423;
  wire[63:0] T424;
  wire[63:0] T425;
  reg [63:0] reg_cause;
  wire[63:0] T426;
  wire T427;
  wire[63:0] T428;
  wire[63:0] T577;
  wire[42:0] T429;
  wire[63:0] T430;
  wire[63:0] T578;
  wire[31:0] T431;
  wire[63:0] T432;
  wire[63:0] T433;
  wire[63:0] T434;
  wire[63:0] T435;
  wire[63:0] T579;
  wire[31:0] T436;
  wire[31:0] read_ptbr;
  wire[18:0] T437;
  wire[63:0] T438;
  wire[63:0] T580;
  wire[42:0] T439;
  reg [42:0] reg_badvaddr;
  wire[42:0] T581;
  wire[43:0] T440;
  wire[43:0] T582;
  wire[43:0] T441;
  wire[43:0] T442;
  wire[42:0] T443;
  wire T444;
  wire T445;
  wire[20:0] T446;
  wire T447;
  wire T448;
  wire[42:0] T449;
  wire T450;
  wire[63:0] T451;
  wire[63:0] T583;
  wire[43:0] T452;
  wire[63:0] T453;
  wire[63:0] T454;
  reg [63:0] reg_sup1;
  wire[63:0] T455;
  wire T456;
  wire T457;
  wire[63:0] T458;
  wire[63:0] T459;
  reg [63:0] reg_sup0;
  wire[63:0] T460;
  wire T461;
  wire T462;
  wire[63:0] T463;
  wire[63:0] T464;
  wire[63:0] T465;
  reg [5:0] R466;
  wire[5:0] T584;
  wire[5:0] T467;
  wire[5:0] T468;
  wire[6:0] T469;
  wire[6:0] T585;
  wire T470;
  reg [57:0] R471;
  wire[57:0] T586;
  wire[57:0] T472;
  wire[57:0] T473;
  wire T474;
  wire T475;
  wire T476;
  wire[63:0] T477;
  wire[63:0] T478;
  wire T479;
  wire[63:0] T480;
  wire[63:0] T481;
  wire T482;
  wire[63:0] T587;
  wire[7:0] T483;
  wire[7:0] T484;
  wire[7:0] T485;
  reg [4:0] reg_fflags;
  wire[4:0] T588;
  wire[63:0] T486;
  wire[63:0] T487;
  wire[63:0] T589;
  wire[4:0] T488;
  wire[4:0] T489;
  wire T490;
  wire T491;
  wire[7:0] T590;
  wire[4:0] T492;
  wire[4:0] T591;
  wire[2:0] T493;
  wire[4:0] T494;
  wire T592;
  wire T495;
  reg  host_pcr_rep_valid;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire temac_manage_io_s_axi_awvalid;
  wire temac_manage_io_s_axi_wvalid;
  wire temac_manage_io_s_axi_bready;
  wire temac_manage_io_s_axi_arvalid;
  wire temac_manage_io_s_axi_rready;
  wire temac_manage_io_sfp_tx_disable;
  wire[7:0] temac_transmit_io_tx_axis_fifo_tdata;
  wire temac_transmit_io_tx_axis_fifo_tvalid;
  wire temac_transmit_io_tx_axis_fifo_tlast;
  wire temac_receive_io_rx_axis_fifo_tready;
  wire[63:0] temac_receive_io_rxd_val;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_data = {2{$random}};
    reg_txd = {2{$random}};
    reg_cfgd = {2{$random}};
    reg_frm = {1{$random}};
    R20 = {1{$random}};
    R28 = {2{$random}};
    reg_epc = {2{$random}};
    reg_evec = {2{$random}};
    reg_ptbr = {1{$random}};
    reg_status_s = {1{$random}};
    reg_status_ps = {1{$random}};
    reg_status_ei = {1{$random}};
    reg_status_pei = {1{$random}};
    reg_status_ef = {1{$random}};
    reg_status_u64 = {1{$random}};
    reg_status_s64 = {1{$random}};
    reg_status_vm = {1{$random}};
    reg_status_er = {1{$random}};
    reg_status_zero = {1{$random}};
    reg_status_im = {1{$random}};
    r_rx_axis_fifo_tvalid = {1{$random}};
    r_irq_ipi = {1{$random}};
    reg_fromhost = {2{$random}};
    r_irq_timer = {1{$random}};
    reg_compare = {1{$random}};
    reg_cfga = {2{$random}};
    R144 = {1{$random}};
    R149 = {2{$random}};
    R158 = {1{$random}};
    R163 = {2{$random}};
    R172 = {1{$random}};
    R177 = {2{$random}};
    R186 = {1{$random}};
    R191 = {2{$random}};
    R200 = {1{$random}};
    R205 = {2{$random}};
    R214 = {1{$random}};
    R219 = {2{$random}};
    R228 = {1{$random}};
    R233 = {2{$random}};
    R242 = {1{$random}};
    R247 = {2{$random}};
    R256 = {1{$random}};
    R261 = {2{$random}};
    R270 = {1{$random}};
    R275 = {2{$random}};
    R284 = {1{$random}};
    R289 = {2{$random}};
    R298 = {1{$random}};
    R303 = {2{$random}};
    R312 = {1{$random}};
    R317 = {2{$random}};
    R326 = {1{$random}};
    R331 = {2{$random}};
    R340 = {1{$random}};
    R345 = {2{$random}};
    R354 = {1{$random}};
    R359 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_cause = {2{$random}};
    reg_badvaddr = {2{$random}};
    reg_sup1 = {2{$random}};
    reg_sup0 = {2{$random}};
    R466 = {1{$random}};
    R471 = {2{$random}};
    reg_fflags = {1{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
`endif

  assign T593 = wen & T367;
  assign T367 = T10[5'h18:5'h18];
  always @(*) case (addr)
    1: T10 = 46'h1;
    2: T10 = 46'h2;
    3: T10 = 46'h4;
    192: T10 = 46'h8;
    1280: T10 = 46'h10;
    1281: T10 = 46'h20;
    1282: T10 = 46'h40;
    1283: T10 = 46'h80;
    1284: T10 = 46'h100;
    1285: T10 = 46'h200;
    1286: T10 = 46'h400;
    1287: T10 = 46'h800;
    1288: T10 = 46'h1000;
    1289: T10 = 46'h2000;
    1290: T10 = 46'h4000;
    1291: T10 = 46'h8000;
    1292: T10 = 46'h10000;
    1293: T10 = 46'h20000;
    1294: T10 = 46'h40000;
    1295: T10 = 46'h80000;
    1309: T10 = 46'h100000;
    1310: T10 = 46'h200000;
    1311: T10 = 46'h400000;
    1312: T10 = 46'h800000;
    1313: T10 = 46'h1000000;
    1314: T10 = 46'h2000000;
    1315: T10 = 46'h4000000;
    3072: T10 = 46'h8000000;
    3073: T10 = 46'h10000000;
    3074: T10 = 46'h20000000;
    3264: T10 = 46'h40000000;
    3265: T10 = 46'h80000000;
    3266: T10 = 46'h100000000;
    3267: T10 = 46'h200000000;
    3268: T10 = 46'h400000000;
    3269: T10 = 46'h800000000;
    3270: T10 = 46'h1000000000;
    3271: T10 = 46'h2000000000;
    3272: T10 = 46'h4000000000;
    3273: T10 = 46'h8000000000;
    3274: T10 = 46'h10000000000;
    3275: T10 = 46'h20000000000;
    3276: T10 = 46'h40000000000;
    3277: T10 = 46'h80000000000;
    3278: T10 = 46'h100000000000;
    3279: T10 = 46'h200000000000;
`ifndef SYNTHESIS
    default: T10 = {2{$random}};
`else
    default: T10 = 46'bx;
`endif
  endcase
  assign addr = cpu_req_valid ? io_rw_addr : T504;
  assign T504 = {1'h0, T12};
  assign T12 = T505 | 11'h500;
  assign T505 = {6'h0, host_pcr_bits_addr};
  assign T13 = T4 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign T4 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign cpu_req_valid = io_rw_cmd != 2'h0;
  assign wen = cpu_req_valid | T14;
  assign T14 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T15 = T4 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign host_pcr_req_fire = host_pcr_req_valid & T5;
  assign T5 = cpu_req_valid ^ 1'h1;
  assign T6 = host_pcr_req_fire ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : host_pcr_req_valid;
  assign T594 = T593 ? wdata : 64'h0;
  assign wdata = cpu_req_valid ? io_rw_wdata : host_pcr_bits_data;
  assign T2 = host_pcr_req_fire ? io_rw_rdata : T3;
  assign T3 = T4 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T371 = wen & T372;
  assign T372 = T10[5'h17:5'h17];
  assign T567 = reset ? 64'h0 : T370;
  assign T370 = T371 ? wdata : reg_txd;
  assign T517 = reset ? 64'h0 : T136;
  assign T136 = T138 ? wdata : T137;
  assign T137 = io_temac_s_axi_rvalid ? T518 : reg_cfgd;
  assign T518 = {32'h0, io_temac_s_axi_rdata};
  assign T138 = wen & T139;
  assign T139 = T10[5'h1a:5'h1a];
  assign T133 = wen & T134;
  assign T134 = T10[5'h19:5'h19];
  assign io_fcsr_rm = reg_frm;
  assign T502 = T0[2'h2:1'h0];
  assign T0 = T17 ? T506 : T1;
  assign T1 = T8 ? wdata : T503;
  assign T503 = {61'h0, reg_frm};
  assign T8 = wen & T9;
  assign T9 = T10[1'h1:1'h1];
  assign T506 = {5'h0, T16};
  assign T16 = wdata >> 3'h5;
  assign T17 = wen & T18;
  assign T18 = T10[2'h2:2'h2];
  assign io_time = T19;
  assign T19 = {R28, R20};
  assign T507 = reset ? 6'h0 : T21;
  assign T21 = T26 ? T24 : T22;
  assign T22 = T23[3'h5:1'h0];
  assign T23 = T508 + 7'h1;
  assign T508 = {1'h0, R20};
  assign T24 = T25[3'h5:1'h0];
  assign T25 = wdata;
  assign T26 = wen & T27;
  assign T27 = T10[4'ha:4'ha];
  assign T509 = reset ? 58'h0 : T29;
  assign T29 = T26 ? T33 : T30;
  assign T30 = T32 ? T31 : R28;
  assign T31 = R28 + 58'h1;
  assign T32 = T23[3'h6:3'h6];
  assign T33 = T25[6'h3f:3'h6];
  assign io_replay = T34;
  assign T34 = io_host_ipi_req_valid & T35;
  assign T35 = io_host_ipi_req_ready ^ 1'h1;
  assign io_fatc = T36;
  assign T36 = wen & T37;
  assign T37 = T10[5'h11:5'h11];
  assign io_evec = T38;
  assign T38 = T39;
  assign T39 = io_exception ? T510 : reg_epc;
  assign T40 = T45 ? T43 : T41;
  assign T41 = io_exception ? T42 : reg_epc;
  assign T42 = io_pc;
  assign T43 = T44;
  assign T44 = wdata[6'h2b:1'h0];
  assign T45 = wen & T46;
  assign T46 = T10[3'h6:3'h6];
  assign T510 = {T511, T47};
  assign T47 = reg_evec;
  assign T48 = T51 ? T49 : reg_evec;
  assign T49 = T50;
  assign T50 = wdata[6'h2a:1'h0];
  assign T51 = wen & T52;
  assign T52 = T10[4'hc:4'hc];
  assign T511 = T47[6'h2a:6'h2a];
  assign io_ptbr = reg_ptbr;
  assign T53 = T57 ? T54 : reg_ptbr;
  assign T54 = T55;
  assign T55 = {T56, 13'h0};
  assign T56 = wdata[5'h1f:4'hd];
  assign T57 = wen & T58;
  assign T58 = T10[4'h8:4'h8];
  assign io_status_s = reg_status_s;
  assign T59 = reset ? 1'h1 : T60;
  assign T60 = T68 ? T67 : T61;
  assign T61 = io_sret ? reg_status_ps : T62;
  assign T62 = io_exception ? 1'h1 : reg_status_s;
  assign T63 = reset ? 1'h0 : T64;
  assign T64 = T68 ? T66 : T65;
  assign T65 = io_exception ? reg_status_s : reg_status_ps;
  assign T66 = wdata[1'h1:1'h1];
  assign T67 = wdata[1'h0:1'h0];
  assign T68 = wen & T69;
  assign T69 = T10[4'he:4'he];
  assign io_status_ps = reg_status_ps;
  assign io_status_ei = reg_status_ei;
  assign T70 = reset ? 1'h0 : T71;
  assign T71 = T68 ? T78 : T72;
  assign T72 = io_sret ? reg_status_pei : T73;
  assign T73 = io_exception ? 1'h0 : reg_status_ei;
  assign T74 = reset ? 1'h0 : T75;
  assign T75 = T68 ? T77 : T76;
  assign T76 = io_exception ? reg_status_ei : reg_status_pei;
  assign T77 = wdata[2'h3:2'h3];
  assign T78 = wdata[2'h2:2'h2];
  assign io_status_pei = reg_status_pei;
  assign io_status_ef = reg_status_ef;
  assign T79 = reset ? 1'h0 : T80;
  assign T80 = T68 ? T81 : reg_status_ef;
  assign T81 = wdata[3'h4:3'h4];
  assign io_status_u64 = reg_status_u64;
  assign T82 = reset ? 1'h1 : T83;
  assign T83 = T68 ? 1'h1 : T84;
  assign T84 = T68 ? T85 : reg_status_u64;
  assign T85 = wdata[3'h5:3'h5];
  assign io_status_s64 = reg_status_s64;
  assign T86 = reset ? 1'h1 : T87;
  assign T87 = T68 ? 1'h1 : T88;
  assign T88 = T68 ? T89 : reg_status_s64;
  assign T89 = wdata[3'h6:3'h6];
  assign io_status_vm = reg_status_vm;
  assign T90 = reset ? 1'h0 : T91;
  assign T91 = T68 ? T92 : reg_status_vm;
  assign T92 = wdata[3'h7:3'h7];
  assign io_status_er = reg_status_er;
  assign T93 = reset ? 1'h0 : T94;
  assign T94 = T68 ? T95 : reg_status_er;
  assign T95 = wdata[4'h8:4'h8];
  assign io_status_zero = reg_status_zero;
  assign T96 = reset ? 7'h0 : T97;
  assign T97 = T68 ? 7'h0 : T98;
  assign T98 = T68 ? T99 : reg_status_zero;
  assign T99 = wdata[4'hf:4'h9];
  assign io_status_im = reg_status_im;
  assign T100 = reset ? 8'h0 : T101;
  assign T101 = T68 ? T102 : reg_status_im;
  assign T102 = wdata[5'h17:5'h10];
  assign io_status_ip = T103;
  assign T103 = {T106, T104};
  assign T104 = {T105, 2'h0};
  assign T105 = {1'h0, io_rocc_interrupt};
  assign T106 = {T113, T107};
  assign T107 = {r_irq_ipi, r_rx_axis_fifo_tvalid};
  assign T512 = reset ? 1'h0 : io_temac_rx_axis_fifo_tvalid;
  assign T513 = reset ? 1'h1 : T108;
  assign T108 = io_host_ipi_rep_valid ? 1'h1 : T109;
  assign T109 = T111 ? T110 : r_irq_ipi;
  assign T110 = wdata[1'h0:1'h0];
  assign T111 = wen & T112;
  assign T112 = T10[5'h13:5'h13];
  assign T113 = {r_irq_timer, T114};
  assign T114 = reg_fromhost != 64'h0;
  assign T514 = reset ? 64'h0 : T115;
  assign T115 = T116 ? wdata : reg_fromhost;
  assign T116 = T120 & T117;
  assign T117 = T119 | T118;
  assign T118 = host_pcr_req_fire ^ 1'h1;
  assign T119 = reg_fromhost == 64'h0;
  assign T120 = wen & T121;
  assign T121 = T10[5'h16:5'h16];
  assign T515 = reset ? 1'h0 : T122;
  assign T122 = T129 ? 1'h0 : T123;
  assign T123 = T124 ? 1'h1 : r_irq_timer;
  assign T124 = T128 == reg_compare;
  assign T125 = T129 ? T126 : reg_compare;
  assign T126 = T127;
  assign T127 = wdata[5'h1f:1'h0];
  assign T128 = T19[5'h1f:1'h0];
  assign T129 = wen & T130;
  assign T130 = T10[4'hb:4'hb];
  assign io_temac_sfp_tx_disable = temac_manage_io_sfp_tx_disable;
  assign io_temac_s_axi_rready = temac_manage_io_s_axi_rready;
  assign io_temac_s_axi_arvalid = temac_manage_io_s_axi_arvalid;
  assign io_temac_s_axi_araddr = T131;
  assign T131 = reg_cfga[4'hb:1'h0];
  assign T516 = reset ? 64'h0 : T132;
  assign T132 = T133 ? wdata : reg_cfga;
  assign io_temac_s_axi_bready = temac_manage_io_s_axi_bready;
  assign io_temac_s_axi_wvalid = temac_manage_io_s_axi_wvalid;
  assign io_temac_s_axi_wdata = T135;
  assign T135 = reg_cfgd[5'h1f:1'h0];
  assign io_temac_s_axi_awvalid = temac_manage_io_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = T140;
  assign T140 = reg_cfga[4'hb:1'h0];
  assign io_temac_tx_axis_fifo_tlast = temac_transmit_io_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = temac_transmit_io_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = temac_transmit_io_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = temac_receive_io_rx_axis_fifo_tready;
  assign io_rw_rdata = T141;
  assign T141 = T155 | T142;
  assign T142 = T154 ? T143 : 64'h0;
  assign T143 = {R149, R144};
  assign T519 = reset ? 6'h0 : T145;
  assign T145 = T148 ? T146 : R144;
  assign T146 = T147[3'h5:1'h0];
  assign T147 = T520 + 7'h1;
  assign T520 = {1'h0, R144};
  assign T148 = io_uarch_counters_15 != 1'h0;
  assign T521 = reset ? 58'h0 : T150;
  assign T150 = T152 ? T151 : R149;
  assign T151 = R149 + 58'h1;
  assign T152 = T148 & T153;
  assign T153 = T147[3'h6:3'h6];
  assign T154 = T10[6'h2d:6'h2d];
  assign T155 = T169 | T156;
  assign T156 = T168 ? T157 : 64'h0;
  assign T157 = {R163, R158};
  assign T522 = reset ? 6'h0 : T159;
  assign T159 = T162 ? T160 : R158;
  assign T160 = T161[3'h5:1'h0];
  assign T161 = T523 + 7'h1;
  assign T523 = {1'h0, R158};
  assign T162 = io_uarch_counters_14 != 1'h0;
  assign T524 = reset ? 58'h0 : T164;
  assign T164 = T166 ? T165 : R163;
  assign T165 = R163 + 58'h1;
  assign T166 = T162 & T167;
  assign T167 = T161[3'h6:3'h6];
  assign T168 = T10[6'h2c:6'h2c];
  assign T169 = T183 | T170;
  assign T170 = T182 ? T171 : 64'h0;
  assign T171 = {R177, R172};
  assign T525 = reset ? 6'h0 : T173;
  assign T173 = T176 ? T174 : R172;
  assign T174 = T175[3'h5:1'h0];
  assign T175 = T526 + 7'h1;
  assign T526 = {1'h0, R172};
  assign T176 = io_uarch_counters_13 != 1'h0;
  assign T527 = reset ? 58'h0 : T178;
  assign T178 = T180 ? T179 : R177;
  assign T179 = R177 + 58'h1;
  assign T180 = T176 & T181;
  assign T181 = T175[3'h6:3'h6];
  assign T182 = T10[6'h2b:6'h2b];
  assign T183 = T197 | T184;
  assign T184 = T196 ? T185 : 64'h0;
  assign T185 = {R191, R186};
  assign T528 = reset ? 6'h0 : T187;
  assign T187 = T190 ? T188 : R186;
  assign T188 = T189[3'h5:1'h0];
  assign T189 = T529 + 7'h1;
  assign T529 = {1'h0, R186};
  assign T190 = io_uarch_counters_12 != 1'h0;
  assign T530 = reset ? 58'h0 : T192;
  assign T192 = T194 ? T193 : R191;
  assign T193 = R191 + 58'h1;
  assign T194 = T190 & T195;
  assign T195 = T189[3'h6:3'h6];
  assign T196 = T10[6'h2a:6'h2a];
  assign T197 = T211 | T198;
  assign T198 = T210 ? T199 : 64'h0;
  assign T199 = {R205, R200};
  assign T531 = reset ? 6'h0 : T201;
  assign T201 = T204 ? T202 : R200;
  assign T202 = T203[3'h5:1'h0];
  assign T203 = T532 + 7'h1;
  assign T532 = {1'h0, R200};
  assign T204 = io_uarch_counters_11 != 1'h0;
  assign T533 = reset ? 58'h0 : T206;
  assign T206 = T208 ? T207 : R205;
  assign T207 = R205 + 58'h1;
  assign T208 = T204 & T209;
  assign T209 = T203[3'h6:3'h6];
  assign T210 = T10[6'h29:6'h29];
  assign T211 = T225 | T212;
  assign T212 = T224 ? T213 : 64'h0;
  assign T213 = {R219, R214};
  assign T534 = reset ? 6'h0 : T215;
  assign T215 = T218 ? T216 : R214;
  assign T216 = T217[3'h5:1'h0];
  assign T217 = T535 + 7'h1;
  assign T535 = {1'h0, R214};
  assign T218 = io_uarch_counters_10 != 1'h0;
  assign T536 = reset ? 58'h0 : T220;
  assign T220 = T222 ? T221 : R219;
  assign T221 = R219 + 58'h1;
  assign T222 = T218 & T223;
  assign T223 = T217[3'h6:3'h6];
  assign T224 = T10[6'h28:6'h28];
  assign T225 = T239 | T226;
  assign T226 = T238 ? T227 : 64'h0;
  assign T227 = {R233, R228};
  assign T537 = reset ? 6'h0 : T229;
  assign T229 = T232 ? T230 : R228;
  assign T230 = T231[3'h5:1'h0];
  assign T231 = T538 + 7'h1;
  assign T538 = {1'h0, R228};
  assign T232 = io_uarch_counters_9 != 1'h0;
  assign T539 = reset ? 58'h0 : T234;
  assign T234 = T236 ? T235 : R233;
  assign T235 = R233 + 58'h1;
  assign T236 = T232 & T237;
  assign T237 = T231[3'h6:3'h6];
  assign T238 = T10[6'h27:6'h27];
  assign T239 = T253 | T240;
  assign T240 = T252 ? T241 : 64'h0;
  assign T241 = {R247, R242};
  assign T540 = reset ? 6'h0 : T243;
  assign T243 = T246 ? T244 : R242;
  assign T244 = T245[3'h5:1'h0];
  assign T245 = T541 + 7'h1;
  assign T541 = {1'h0, R242};
  assign T246 = io_uarch_counters_8 != 1'h0;
  assign T542 = reset ? 58'h0 : T248;
  assign T248 = T250 ? T249 : R247;
  assign T249 = R247 + 58'h1;
  assign T250 = T246 & T251;
  assign T251 = T245[3'h6:3'h6];
  assign T252 = T10[6'h26:6'h26];
  assign T253 = T267 | T254;
  assign T254 = T266 ? T255 : 64'h0;
  assign T255 = {R261, R256};
  assign T543 = reset ? 6'h0 : T257;
  assign T257 = T260 ? T258 : R256;
  assign T258 = T259[3'h5:1'h0];
  assign T259 = T544 + 7'h1;
  assign T544 = {1'h0, R256};
  assign T260 = io_uarch_counters_7 != 1'h0;
  assign T545 = reset ? 58'h0 : T262;
  assign T262 = T264 ? T263 : R261;
  assign T263 = R261 + 58'h1;
  assign T264 = T260 & T265;
  assign T265 = T259[3'h6:3'h6];
  assign T266 = T10[6'h25:6'h25];
  assign T267 = T281 | T268;
  assign T268 = T280 ? T269 : 64'h0;
  assign T269 = {R275, R270};
  assign T546 = reset ? 6'h0 : T271;
  assign T271 = T274 ? T272 : R270;
  assign T272 = T273[3'h5:1'h0];
  assign T273 = T547 + 7'h1;
  assign T547 = {1'h0, R270};
  assign T274 = io_uarch_counters_6 != 1'h0;
  assign T548 = reset ? 58'h0 : T276;
  assign T276 = T278 ? T277 : R275;
  assign T277 = R275 + 58'h1;
  assign T278 = T274 & T279;
  assign T279 = T273[3'h6:3'h6];
  assign T280 = T10[6'h24:6'h24];
  assign T281 = T295 | T282;
  assign T282 = T294 ? T283 : 64'h0;
  assign T283 = {R289, R284};
  assign T549 = reset ? 6'h0 : T285;
  assign T285 = T288 ? T286 : R284;
  assign T286 = T287[3'h5:1'h0];
  assign T287 = T550 + 7'h1;
  assign T550 = {1'h0, R284};
  assign T288 = io_uarch_counters_5 != 1'h0;
  assign T551 = reset ? 58'h0 : T290;
  assign T290 = T292 ? T291 : R289;
  assign T291 = R289 + 58'h1;
  assign T292 = T288 & T293;
  assign T293 = T287[3'h6:3'h6];
  assign T294 = T10[6'h23:6'h23];
  assign T295 = T309 | T296;
  assign T296 = T308 ? T297 : 64'h0;
  assign T297 = {R303, R298};
  assign T552 = reset ? 6'h0 : T299;
  assign T299 = T302 ? T300 : R298;
  assign T300 = T301[3'h5:1'h0];
  assign T301 = T553 + 7'h1;
  assign T553 = {1'h0, R298};
  assign T302 = io_uarch_counters_4 != 1'h0;
  assign T554 = reset ? 58'h0 : T304;
  assign T304 = T306 ? T305 : R303;
  assign T305 = R303 + 58'h1;
  assign T306 = T302 & T307;
  assign T307 = T301[3'h6:3'h6];
  assign T308 = T10[6'h22:6'h22];
  assign T309 = T323 | T310;
  assign T310 = T322 ? T311 : 64'h0;
  assign T311 = {R317, R312};
  assign T555 = reset ? 6'h0 : T313;
  assign T313 = T316 ? T314 : R312;
  assign T314 = T315[3'h5:1'h0];
  assign T315 = T556 + 7'h1;
  assign T556 = {1'h0, R312};
  assign T316 = io_uarch_counters_3 != 1'h0;
  assign T557 = reset ? 58'h0 : T318;
  assign T318 = T320 ? T319 : R317;
  assign T319 = R317 + 58'h1;
  assign T320 = T316 & T321;
  assign T321 = T315[3'h6:3'h6];
  assign T322 = T10[6'h21:6'h21];
  assign T323 = T337 | T324;
  assign T324 = T336 ? T325 : 64'h0;
  assign T325 = {R331, R326};
  assign T558 = reset ? 6'h0 : T327;
  assign T327 = T330 ? T328 : R326;
  assign T328 = T329[3'h5:1'h0];
  assign T329 = T559 + 7'h1;
  assign T559 = {1'h0, R326};
  assign T330 = io_uarch_counters_2 != 1'h0;
  assign T560 = reset ? 58'h0 : T332;
  assign T332 = T334 ? T333 : R331;
  assign T333 = R331 + 58'h1;
  assign T334 = T330 & T335;
  assign T335 = T329[3'h6:3'h6];
  assign T336 = T10[6'h20:6'h20];
  assign T337 = T351 | T338;
  assign T338 = T350 ? T339 : 64'h0;
  assign T339 = {R345, R340};
  assign T561 = reset ? 6'h0 : T341;
  assign T341 = T344 ? T342 : R340;
  assign T342 = T343[3'h5:1'h0];
  assign T343 = T562 + 7'h1;
  assign T562 = {1'h0, R340};
  assign T344 = io_uarch_counters_1 != 1'h0;
  assign T563 = reset ? 58'h0 : T346;
  assign T346 = T348 ? T347 : R345;
  assign T347 = R345 + 58'h1;
  assign T348 = T344 & T349;
  assign T349 = T343[3'h6:3'h6];
  assign T350 = T10[5'h1f:5'h1f];
  assign T351 = T365 | T352;
  assign T352 = T364 ? T353 : 64'h0;
  assign T353 = {R359, R354};
  assign T564 = reset ? 6'h0 : T355;
  assign T355 = T358 ? T356 : R354;
  assign T356 = T357[3'h5:1'h0];
  assign T357 = T565 + 7'h1;
  assign T565 = {1'h0, R354};
  assign T358 = io_uarch_counters_0 != 1'h0;
  assign T566 = reset ? 58'h0 : T360;
  assign T360 = T362 ? T361 : R359;
  assign T361 = R359 + 58'h1;
  assign T362 = T358 & T363;
  assign T363 = T357[3'h6:3'h6];
  assign T364 = T10[5'h1e:5'h1e];
  assign T365 = T368 | T366;
  assign T366 = T367 ? temac_receive_io_rxd_val : 64'h0;
  assign T368 = T373 | T369;
  assign T369 = T372 ? reg_txd : 64'h0;
  assign T373 = T375 | T374;
  assign T374 = T139 ? reg_cfgd : 64'h0;
  assign T375 = T377 | T376;
  assign T376 = T134 ? reg_cfga : 64'h0;
  assign T377 = T379 | T378;
  assign T378 = T121 ? reg_fromhost : 64'h0;
  assign T379 = T391 | T380;
  assign T380 = T390 ? reg_tohost : 64'h0;
  assign T568 = reset ? 64'h0 : T381;
  assign T381 = T386 ? wdata : T382;
  assign T382 = T383 ? 64'h0 : reg_tohost;
  assign T383 = T384 & T390;
  assign T384 = host_pcr_req_fire & T385;
  assign T385 = host_pcr_bits_rw ^ 1'h1;
  assign T386 = T389 & T387;
  assign T387 = T388 | host_pcr_req_fire;
  assign T388 = reg_tohost == 64'h0;
  assign T389 = wen & T390;
  assign T390 = T10[5'h15:5'h15];
  assign T391 = T397 | T569;
  assign T569 = {63'h0, T392};
  assign T392 = T396 ? reg_stats : 1'h0;
  assign T570 = reset ? 1'h0 : T393;
  assign T393 = T395 ? T394 : reg_stats;
  assign T394 = wdata[1'h0:1'h0];
  assign T395 = wen & T396;
  assign T396 = T10[2'h3:2'h3];
  assign T397 = T399 | T571;
  assign T571 = {62'h0, T398};
  assign T398 = T112 ? 2'h2 : 2'h0;
  assign T399 = T402 | T572;
  assign T572 = {62'h0, T400};
  assign T400 = T401 ? 2'h2 : 2'h0;
  assign T401 = T10[5'h12:5'h12];
  assign T402 = T404 | T573;
  assign T573 = {62'h0, T403};
  assign T403 = T37 ? 2'h2 : 2'h0;
  assign T404 = T407 | T574;
  assign T574 = {62'h0, T405};
  assign T405 = T406 ? 2'h2 : 2'h0;
  assign T406 = T10[5'h10:5'h10];
  assign T407 = T410 | T575;
  assign T575 = {63'h0, T408};
  assign T408 = T409 ? io_host_id : 1'h0;
  assign T409 = T10[4'hf:4'hf];
  assign T410 = T424 | T576;
  assign T576 = {32'h0, T411};
  assign T411 = T69 ? T412 : 32'h0;
  assign T412 = T413;
  assign T413 = {T419, T414};
  assign T414 = {T417, T415};
  assign T415 = {io_status_ei, T416};
  assign T416 = {io_status_ps, io_status_s};
  assign T417 = {io_status_u64, T418};
  assign T418 = {io_status_ef, io_status_pei};
  assign T419 = {T422, T420};
  assign T420 = {io_status_er, T421};
  assign T421 = {io_status_vm, io_status_s64};
  assign T422 = {io_status_ip, T423};
  assign T423 = {io_status_im, io_status_zero};
  assign T424 = T428 | T425;
  assign T425 = T427 ? reg_cause : 64'h0;
  assign T426 = io_exception ? io_cause : reg_cause;
  assign T427 = T10[4'hd:4'hd];
  assign T428 = T430 | T577;
  assign T577 = {21'h0, T429};
  assign T429 = T52 ? reg_evec : 43'h0;
  assign T430 = T432 | T578;
  assign T578 = {32'h0, T431};
  assign T431 = T130 ? reg_compare : 32'h0;
  assign T432 = T434 | T433;
  assign T433 = T27 ? T19 : 64'h0;
  assign T434 = T435 | 64'h0;
  assign T435 = T438 | T579;
  assign T579 = {32'h0, T436};
  assign T436 = T58 ? read_ptbr : 32'h0;
  assign read_ptbr = T437 << 4'hd;
  assign T437 = reg_ptbr[5'h1f:4'hd];
  assign T438 = T451 | T580;
  assign T580 = {21'h0, T439};
  assign T439 = T450 ? reg_badvaddr : 43'h0;
  assign T581 = T440[6'h2a:1'h0];
  assign T440 = io_badvaddr_wen ? T441 : T582;
  assign T582 = {1'h0, reg_badvaddr};
  assign T441 = T442;
  assign T442 = {T444, T443};
  assign T443 = io_rw_wdata[6'h2a:1'h0];
  assign T444 = T448 ? T447 : T445;
  assign T445 = T446 != 21'h0;
  assign T446 = io_rw_wdata[6'h3f:6'h2b];
  assign T447 = T446 == 21'h1fffff;
  assign T448 = $signed(T449) < $signed(1'h0);
  assign T449 = T443;
  assign T450 = T10[3'h7:3'h7];
  assign T451 = T453 | T583;
  assign T583 = {20'h0, T452};
  assign T452 = T46 ? reg_epc : 44'h0;
  assign T453 = T458 | T454;
  assign T454 = T457 ? reg_sup1 : 64'h0;
  assign T455 = T456 ? wdata : reg_sup1;
  assign T456 = wen & T457;
  assign T457 = T10[3'h5:3'h5];
  assign T458 = T463 | T459;
  assign T459 = T462 ? reg_sup0 : 64'h0;
  assign T460 = T461 ? wdata : reg_sup0;
  assign T461 = wen & T462;
  assign T462 = T10[3'h4:3'h4];
  assign T463 = T477 | T464;
  assign T464 = T476 ? T465 : 64'h0;
  assign T465 = {R471, R466};
  assign T584 = reset ? 6'h0 : T467;
  assign T467 = T470 ? T468 : R466;
  assign T468 = T469[3'h5:1'h0];
  assign T469 = T585 + 7'h1;
  assign T585 = {1'h0, R466};
  assign T470 = io_retire != 1'h0;
  assign T586 = reset ? 58'h0 : T472;
  assign T472 = T474 ? T473 : R471;
  assign T473 = R471 + 58'h1;
  assign T474 = T470 & T475;
  assign T475 = T469[3'h6:3'h6];
  assign T476 = T10[5'h1d:5'h1d];
  assign T477 = T480 | T478;
  assign T478 = T479 ? T19 : 64'h0;
  assign T479 = T10[5'h1c:5'h1c];
  assign T480 = T587 | T481;
  assign T481 = T482 ? T19 : 64'h0;
  assign T482 = T10[5'h1b:5'h1b];
  assign T587 = {56'h0, T483};
  assign T483 = T590 | T484;
  assign T484 = T18 ? T485 : 8'h0;
  assign T485 = {reg_frm, reg_fflags};
  assign T588 = T486[3'h4:1'h0];
  assign T486 = T17 ? wdata : T487;
  assign T487 = T490 ? wdata : T589;
  assign T589 = {59'h0, T488};
  assign T488 = io_fcsr_flags_valid ? T489 : reg_fflags;
  assign T489 = reg_fflags | io_fcsr_flags_bits;
  assign T490 = wen & T491;
  assign T491 = T10[1'h0:1'h0];
  assign T590 = {3'h0, T492};
  assign T492 = T494 | T591;
  assign T591 = {2'h0, T493};
  assign T493 = T9 ? reg_frm : 3'h0;
  assign T494 = T491 ? reg_fflags : 5'h0;
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T592;
  assign T592 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T495;
  assign T495 = cpu_req_valid & T401;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T496 = T498 ? 1'h0 : T497;
  assign T497 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T498 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T499;
  assign T499 = T501 & T500;
  assign T500 = host_pcr_rep_valid ^ 1'h1;
  assign T501 = host_pcr_req_valid ^ 1'h1;
  ManagementMachine temac_manage(.clk(clk), .reset(reset),
       //.io_stall_out(  )
       .io_write_to_cfga( T133 ),
       .io_cfgd_in( reg_cfgd ),
       .io_s_axi_awvalid( temac_manage_io_s_axi_awvalid ),
       .io_s_axi_awready( io_temac_s_axi_awready ),
       .io_s_axi_wvalid( temac_manage_io_s_axi_wvalid ),
       .io_s_axi_wready( io_temac_s_axi_wready ),
       .io_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_s_axi_bready( temac_manage_io_s_axi_bready ),
       .io_s_axi_arvalid( temac_manage_io_s_axi_arvalid ),
       .io_s_axi_arready( io_temac_s_axi_arready ),
       .io_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_s_axi_rready( temac_manage_io_s_axi_rready ),
       .io_sfp_tx_disable( temac_manage_io_sfp_tx_disable )
  );
  TransmitMachine temac_transmit(.clk(clk), .reset(reset),
       .io_tx_axis_fifo_tdata( temac_transmit_io_tx_axis_fifo_tdata ),
       .io_tx_axis_fifo_tvalid( temac_transmit_io_tx_axis_fifo_tvalid ),
       .io_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_tx_axis_fifo_tlast( temac_transmit_io_tx_axis_fifo_tlast ),
       .io_txd_in( reg_txd ),
       .io_write_to_txd( T371 )
  );
  ReceiveMachine temac_receive(.clk(clk), .reset(reset),
       .io_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_rx_axis_fifo_tready( temac_receive_io_rx_axis_fifo_tready ),
       .io_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_rxd_val( temac_receive_io_rxd_val ),
       .io_rxd_val_in( T594 ),
       .io_rxd_val_in_valid( T593 )
  );

  always @(posedge clk) begin
    if(T4) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T4) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T4) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T4) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(reset) begin
      reg_txd <= 64'h0;
    end else if(T371) begin
      reg_txd <= wdata;
    end
    if(reset) begin
      reg_cfgd <= 64'h0;
    end else if(T138) begin
      reg_cfgd <= wdata;
    end else if(io_temac_s_axi_rvalid) begin
      reg_cfgd <= T518;
    end
    reg_frm <= T502;
    if(reset) begin
      R20 <= 6'h0;
    end else if(T26) begin
      R20 <= T24;
    end else begin
      R20 <= T22;
    end
    if(reset) begin
      R28 <= 58'h0;
    end else if(T26) begin
      R28 <= T33;
    end else if(T32) begin
      R28 <= T31;
    end
    if(T45) begin
      reg_epc <= T43;
    end else if(io_exception) begin
      reg_epc <= T42;
    end
    if(T51) begin
      reg_evec <= T49;
    end
    if(T57) begin
      reg_ptbr <= T54;
    end
    if(reset) begin
      reg_status_s <= 1'h1;
    end else if(T68) begin
      reg_status_s <= T67;
    end else if(io_sret) begin
      reg_status_s <= reg_status_ps;
    end else if(io_exception) begin
      reg_status_s <= 1'h1;
    end
    if(reset) begin
      reg_status_ps <= 1'h0;
    end else if(T68) begin
      reg_status_ps <= T66;
    end else if(io_exception) begin
      reg_status_ps <= reg_status_s;
    end
    if(reset) begin
      reg_status_ei <= 1'h0;
    end else if(T68) begin
      reg_status_ei <= T78;
    end else if(io_sret) begin
      reg_status_ei <= reg_status_pei;
    end else if(io_exception) begin
      reg_status_ei <= 1'h0;
    end
    if(reset) begin
      reg_status_pei <= 1'h0;
    end else if(T68) begin
      reg_status_pei <= T77;
    end else if(io_exception) begin
      reg_status_pei <= reg_status_ei;
    end
    if(reset) begin
      reg_status_ef <= 1'h0;
    end else if(T68) begin
      reg_status_ef <= T81;
    end
    if(reset) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= T85;
    end
    if(reset) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= T89;
    end
    if(reset) begin
      reg_status_vm <= 1'h0;
    end else if(T68) begin
      reg_status_vm <= T92;
    end
    if(reset) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= T95;
    end
    if(reset) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= T99;
    end
    if(reset) begin
      reg_status_im <= 8'h0;
    end else if(T68) begin
      reg_status_im <= T102;
    end
    if(reset) begin
      r_rx_axis_fifo_tvalid <= 1'h0;
    end else begin
      r_rx_axis_fifo_tvalid <= io_temac_rx_axis_fifo_tvalid;
    end
    if(reset) begin
      r_irq_ipi <= 1'h1;
    end else if(io_host_ipi_rep_valid) begin
      r_irq_ipi <= 1'h1;
    end else if(T111) begin
      r_irq_ipi <= T110;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T116) begin
      reg_fromhost <= wdata;
    end
    if(reset) begin
      r_irq_timer <= 1'h0;
    end else if(T129) begin
      r_irq_timer <= 1'h0;
    end else if(T124) begin
      r_irq_timer <= 1'h1;
    end
    if(T129) begin
      reg_compare <= T126;
    end
    if(reset) begin
      reg_cfga <= 64'h0;
    end else if(T133) begin
      reg_cfga <= wdata;
    end
    if(reset) begin
      R144 <= 6'h0;
    end else if(T148) begin
      R144 <= T146;
    end
    if(reset) begin
      R149 <= 58'h0;
    end else if(T152) begin
      R149 <= T151;
    end
    if(reset) begin
      R158 <= 6'h0;
    end else if(T162) begin
      R158 <= T160;
    end
    if(reset) begin
      R163 <= 58'h0;
    end else if(T166) begin
      R163 <= T165;
    end
    if(reset) begin
      R172 <= 6'h0;
    end else if(T176) begin
      R172 <= T174;
    end
    if(reset) begin
      R177 <= 58'h0;
    end else if(T180) begin
      R177 <= T179;
    end
    if(reset) begin
      R186 <= 6'h0;
    end else if(T190) begin
      R186 <= T188;
    end
    if(reset) begin
      R191 <= 58'h0;
    end else if(T194) begin
      R191 <= T193;
    end
    if(reset) begin
      R200 <= 6'h0;
    end else if(T204) begin
      R200 <= T202;
    end
    if(reset) begin
      R205 <= 58'h0;
    end else if(T208) begin
      R205 <= T207;
    end
    if(reset) begin
      R214 <= 6'h0;
    end else if(T218) begin
      R214 <= T216;
    end
    if(reset) begin
      R219 <= 58'h0;
    end else if(T222) begin
      R219 <= T221;
    end
    if(reset) begin
      R228 <= 6'h0;
    end else if(T232) begin
      R228 <= T230;
    end
    if(reset) begin
      R233 <= 58'h0;
    end else if(T236) begin
      R233 <= T235;
    end
    if(reset) begin
      R242 <= 6'h0;
    end else if(T246) begin
      R242 <= T244;
    end
    if(reset) begin
      R247 <= 58'h0;
    end else if(T250) begin
      R247 <= T249;
    end
    if(reset) begin
      R256 <= 6'h0;
    end else if(T260) begin
      R256 <= T258;
    end
    if(reset) begin
      R261 <= 58'h0;
    end else if(T264) begin
      R261 <= T263;
    end
    if(reset) begin
      R270 <= 6'h0;
    end else if(T274) begin
      R270 <= T272;
    end
    if(reset) begin
      R275 <= 58'h0;
    end else if(T278) begin
      R275 <= T277;
    end
    if(reset) begin
      R284 <= 6'h0;
    end else if(T288) begin
      R284 <= T286;
    end
    if(reset) begin
      R289 <= 58'h0;
    end else if(T292) begin
      R289 <= T291;
    end
    if(reset) begin
      R298 <= 6'h0;
    end else if(T302) begin
      R298 <= T300;
    end
    if(reset) begin
      R303 <= 58'h0;
    end else if(T306) begin
      R303 <= T305;
    end
    if(reset) begin
      R312 <= 6'h0;
    end else if(T316) begin
      R312 <= T314;
    end
    if(reset) begin
      R317 <= 58'h0;
    end else if(T320) begin
      R317 <= T319;
    end
    if(reset) begin
      R326 <= 6'h0;
    end else if(T330) begin
      R326 <= T328;
    end
    if(reset) begin
      R331 <= 58'h0;
    end else if(T334) begin
      R331 <= T333;
    end
    if(reset) begin
      R340 <= 6'h0;
    end else if(T344) begin
      R340 <= T342;
    end
    if(reset) begin
      R345 <= 58'h0;
    end else if(T348) begin
      R345 <= T347;
    end
    if(reset) begin
      R354 <= 6'h0;
    end else if(T358) begin
      R354 <= T356;
    end
    if(reset) begin
      R359 <= 58'h0;
    end else if(T362) begin
      R359 <= T361;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T386) begin
      reg_tohost <= wdata;
    end else if(T383) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T395) begin
      reg_stats <= T394;
    end
    if(io_exception) begin
      reg_cause <= io_cause;
    end
    reg_badvaddr <= T581;
    if(T456) begin
      reg_sup1 <= wdata;
    end
    if(T461) begin
      reg_sup0 <= wdata;
    end
    if(reset) begin
      R466 <= 6'h0;
    end else if(T470) begin
      R466 <= T468;
    end
    if(reset) begin
      R471 <= 58'h0;
    end else if(T474) begin
      R471 <= T473;
    end
    reg_fflags <= T588;
    if(T498) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module Datapath(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [2:0] io_ctrl_sel_pc,
    input  io_ctrl_killd,
    input  io_ctrl_ren_1,
    input  io_ctrl_ren_0,
    input [2:0] io_ctrl_sel_alu2,
    input [1:0] io_ctrl_sel_alu1,
    input [2:0] io_ctrl_sel_imm,
    input  io_ctrl_fn_dw,
    input [3:0] io_ctrl_fn_alu,
    input  io_ctrl_div_mul_val,
    input  io_ctrl_div_mul_kill,
    //input  io_ctrl_div_val
    //input  io_ctrl_div_kill
    input [2:0] io_ctrl_csr,
    input  io_ctrl_sret,
    input  io_ctrl_mem_load,
    input  io_ctrl_wb_load,
    input  io_ctrl_ex_fp_val,
    input  io_ctrl_mem_fp_val,
    input  io_ctrl_ex_wen,
    input  io_ctrl_ex_valid,
    input  io_ctrl_mem_jalr,
    input  io_ctrl_mem_branch,
    input  io_ctrl_mem_wen,
    input  io_ctrl_wb_wen,
    input [2:0] io_ctrl_ex_mem_type,
    input  io_ctrl_ex_rs2_val,
    input  io_ctrl_ex_rocc_val,
    input  io_ctrl_mem_rocc_val,
    input  io_ctrl_bypass_1,
    input  io_ctrl_bypass_0,
    input [1:0] io_ctrl_bypass_src_1,
    input [1:0] io_ctrl_bypass_src_0,
    input  io_ctrl_ll_ready,
    input  io_ctrl_retire,
    input  io_ctrl_exception,
    input [63:0] io_ctrl_cause,
    input  io_ctrl_badvaddr_wen,
    output[31:0] io_ctrl_inst,
    //output io_ctrl_jalr_eq
    output io_ctrl_mem_br_taken,
    output io_ctrl_mem_misprediction,
    output io_ctrl_div_mul_rdy,
    output io_ctrl_ll_wen,
    output[4:0] io_ctrl_ll_waddr,
    output[4:0] io_ctrl_ex_waddr,
    output io_ctrl_mem_rs1_ra,
    output[4:0] io_ctrl_mem_waddr,
    output[4:0] io_ctrl_wb_waddr,
    output[7:0] io_ctrl_status_ip,
    output[7:0] io_ctrl_status_im,
    output[6:0] io_ctrl_status_zero,
    output io_ctrl_status_er,
    output io_ctrl_status_vm,
    output io_ctrl_status_s64,
    output io_ctrl_status_u64,
    output io_ctrl_status_ef,
    output io_ctrl_status_pei,
    output io_ctrl_status_ei,
    output io_ctrl_status_ps,
    output io_ctrl_status_s,
    output io_ctrl_fp_sboard_clr,
    output[4:0] io_ctrl_fp_sboard_clra,
    output io_ctrl_csr_replay,
    input  io_dmem_req_ready,
    //output io_dmem_req_valid
    //output io_dmem_req_bits_kill
    //output[2:0] io_dmem_req_bits_typ
    //output io_dmem_req_bits_phys
    output[43:0] io_dmem_req_bits_addr,
    output[8:0] io_dmem_req_bits_tag,
    //output[4:0] io_dmem_req_bits_cmd
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [8:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [8:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    //output io_imem_req_valid
    output[43:0] io_imem_req_bits_pc,
    //output io_imem_resp_ready
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    //output io_imem_btb_update_valid
    //output io_imem_btb_update_bits_prediction_valid
    //output io_imem_btb_update_bits_prediction_bits_taken
    //output[42:0] io_imem_btb_update_bits_prediction_bits_target
    //output[5:0] io_imem_btb_update_bits_prediction_bits_entry
    //output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history
    //output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    //output io_imem_btb_update_bits_taken
    //output io_imem_btb_update_bits_isJump
    //output io_imem_btb_update_bits_isCall
    //output io_imem_btb_update_bits_isReturn
    //output io_imem_btb_update_bits_mispredict
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    //output io_imem_invalidate
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    output io_rocc_resp_ready,
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [2:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [511:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[2:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready,
    output io_temac_sfp_tx_disable
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  reg  ex_reg_kill;
  wire T7;
  reg  mem_reg_kill;
  wire[31:0] T8;
  wire[63:0] T9;
  reg [63:0] R10;
  reg [63:0] R11;
  wire[63:0] ex_rs_1;
  wire[63:0] T12;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[63:0] id_rs_1;
  wire[63:0] T16;
  wire[63:0] T17;
  reg [63:0] T18 [30:0];
  wire[63:0] T19;
  wire T20;
  wire T21;
  wire[4:0] T22;
  wire T23;
  wire T24;
  wire[4:0] wb_waddr;
  wire wb_wen;
  wire[4:0] T25;
  wire[4:0] T26;
  wire[4:0] T27;
  wire[63:0] wb_wdata;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  reg [63:0] wb_reg_wdata;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] mem_int_wdata;
  reg [63:0] mem_reg_wdata;
  wire[63:0] T33;
  wire[63:0] T205;
  wire[44:0] mem_br_target;
  wire[44:0] T34;
  wire[44:0] T35;
  reg [43:0] mem_reg_pc;
  wire[43:0] T36;
  reg [43:0] ex_reg_pc;
  wire[43:0] T37;
  wire[44:0] T206;
  wire[21:0] T38;
  wire[21:0] T39;
  wire[21:0] T40;
  wire[21:0] T41;
  wire[11:0] T42;
  wire[4:0] T43;
  wire[3:0] T44;
  wire[6:0] T45;
  wire[5:0] T46;
  wire T47;
  wire T48;
  wire[9:0] T49;
  wire[8:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[21:0] T207;
  wire[14:0] T58;
  wire[14:0] T59;
  wire[11:0] T60;
  wire[4:0] T61;
  wire[3:0] T62;
  wire[6:0] T63;
  wire[5:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire[6:0] T208;
  wire T209;
  wire T71;
  wire[22:0] T210;
  wire T211;
  wire[18:0] T212;
  wire T213;
  wire T72;
  wire T73;
  wire[63:0] ll_wdata;
  wire[63:0] T74;
  wire T75;
  wire T76;
  wire dmem_resp_xpu;
  wire T77;
  wire T78;
  wire dmem_resp_valid;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T83;
  wire[61:0] T84;
  wire T85;
  wire T86;
  wire[63:0] T87;
  wire[63:0] T88;
  wire[63:0] T214;
  wire bypass_0;
  wire[63:0] bypass_1;
  wire T89;
  wire[1:0] T90;
  wire[63:0] T91;
  wire[63:0] bypass_2;
  wire[63:0] bypass_3;
  wire T92;
  wire T93;
  reg  ex_reg_rs_bypass_1;
  wire T94;
  wire[4:0] T95;
  wire[4:0] T96;
  wire[63:0] T97;
  reg [63:0] R98;
  reg [63:0] R99;
  wire[63:0] ex_rs_0;
  wire[63:0] T100;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T101;
  wire[1:0] T102;
  wire[1:0] T103;
  wire[63:0] id_rs_0;
  wire[63:0] T104;
  wire[63:0] T105;
  wire[4:0] T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T112;
  wire[61:0] T113;
  wire T114;
  wire T115;
  wire[63:0] T116;
  wire[63:0] T117;
  wire[63:0] T215;
  wire T118;
  wire[1:0] T119;
  wire[63:0] T120;
  wire T121;
  wire T122;
  reg  ex_reg_rs_bypass_0;
  wire T123;
  wire[4:0] T124;
  wire[4:0] T125;
  wire T126;
  wire[63:0] T127;
  wire[4:0] T128;
  wire[4:0] T129;
  wire[43:0] T130;
  reg [43:0] wb_reg_pc;
  wire[43:0] T131;
  wire T132;
  wire[32:0] T133;
  wire[32:0] T134;
  wire T135;
  wire[1135:0] T136;
  wire[63:0] T228;
  wire[63:0] T229;
  wire[63:0] T230;
  wire[63:0] T231;
  wire T232;
  wire[63:0] T233;
  wire T234;
  wire[1:0] T235;
  wire[11:0] T236;
  wire T237;
  wire T238;
  wire T138;
  wire dmem_resp_replay;
  reg  ex_reg_ctrl_fn_dw;
  wire T239;
  wire T240;
  reg [3:0] ex_reg_ctrl_fn_alu;
  wire[3:0] T241;
  wire[63:0] ex_op1;
  wire[63:0] T242;
  wire[43:0] T243;
  wire[43:0] T244;
  wire T245;
  reg [1:0] ex_reg_sel_alu1;
  wire[1:0] T246;
  wire[19:0] T247;
  wire T248;
  wire[63:0] T249;
  wire T250;
  wire[63:0] T251;
  wire[63:0] ex_op2;
  wire[63:0] T252;
  wire[31:0] T253;
  wire[31:0] T254;
  wire[3:0] T255;
  wire T256;
  reg [2:0] ex_reg_sel_alu2;
  wire[2:0] T257;
  wire[27:0] T258;
  wire T259;
  wire[31:0] ex_imm;
  wire[31:0] T260;
  wire[11:0] T261;
  wire[4:0] T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  reg [2:0] ex_reg_sel_imm;
  wire[2:0] T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[3:0] T273;
  wire[3:0] T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire T278;
  wire[3:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[6:0] T284;
  wire[5:0] T285;
  wire[5:0] T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire[19:0] T304;
  wire[18:0] T305;
  wire[7:0] T306;
  wire[7:0] T307;
  wire[7:0] T308;
  wire[7:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[10:0] T313;
  wire[10:0] T314;
  wire[10:0] T315;
  wire[10:0] T316;
  wire T317;
  wire T318;
  wire[31:0] T319;
  wire T320;
  wire[63:0] T321;
  wire T322;
  wire T137;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T139;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T140;
  wire[6:0] T141;
  wire[4:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire[4:0] T147;
  wire[6:0] T148;
  wire[4:0] T216;
  wire[7:0] dmem_resp_waddr;
  wire[8:0] T149;
  wire T150;
  wire dmem_resp_fpu;
  wire T151;
  wire[42:0] T217;
  wire[42:0] T218;
  wire[42:0] T219;
  wire[43:0] T220;
  wire[44:0] T152;
  wire[44:0] T153;
  wire[44:0] T221;
  wire[43:0] T154;
  wire T155;
  wire[44:0] mem_npc;
  wire[44:0] T222;
  wire[43:0] T156;
  wire[42:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[1:0] T161;
  wire T162;
  wire T163;
  wire T164;
  wire[21:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire[63:0] T172;
  wire[8:0] T223;
  wire[5:0] T173;
  wire[43:0] T174;
  wire[43:0] T175;
  wire[42:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire[21:0] T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire[4:0] T224;
  wire T190;
  wire[4:0] T191;
  wire[4:0] T192;
  wire T193;
  wire[4:0] T194;
  wire[4:0] T195;
  wire[4:0] T225;
  wire[7:0] T196;
  wire[7:0] T226;
  wire[4:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[44:0] T227;
  wire T204;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;
  wire pcr_io_host_pcr_req_ready;
  wire pcr_io_host_pcr_rep_valid;
  wire[63:0] pcr_io_host_pcr_rep_bits;
  wire pcr_io_host_ipi_req_valid;
  wire pcr_io_host_ipi_req_bits;
  wire pcr_io_host_ipi_rep_ready;
  wire pcr_io_host_debug_stats_pcr;
  wire[63:0] pcr_io_rw_rdata;
  wire pcr_io_temac_rx_axis_fifo_tready;
  wire[7:0] pcr_io_temac_tx_axis_fifo_tdata;
  wire pcr_io_temac_tx_axis_fifo_tvalid;
  wire pcr_io_temac_tx_axis_fifo_tlast;
  wire[11:0] pcr_io_temac_s_axi_awaddr;
  wire pcr_io_temac_s_axi_awvalid;
  wire[31:0] pcr_io_temac_s_axi_wdata;
  wire pcr_io_temac_s_axi_wvalid;
  wire pcr_io_temac_s_axi_bready;
  wire[11:0] pcr_io_temac_s_axi_araddr;
  wire pcr_io_temac_s_axi_arvalid;
  wire pcr_io_temac_s_axi_rready;
  wire pcr_io_temac_sfp_tx_disable;
  wire[7:0] pcr_io_status_ip;
  wire[7:0] pcr_io_status_im;
  wire[6:0] pcr_io_status_zero;
  wire pcr_io_status_er;
  wire pcr_io_status_vm;
  wire pcr_io_status_s64;
  wire pcr_io_status_u64;
  wire pcr_io_status_ef;
  wire pcr_io_status_pei;
  wire pcr_io_status_ei;
  wire pcr_io_status_ps;
  wire pcr_io_status_s;
  wire[31:0] pcr_io_ptbr;
  wire[43:0] pcr_io_evec;
  wire pcr_io_fatc;
  wire pcr_io_replay;
  wire[63:0] pcr_io_time;
  wire[2:0] pcr_io_fcsr_rm;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_kill = {1{$random}};
    mem_reg_kill = {1{$random}};
    R10 = {2{$random}};
    R11 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T18[initvar] = {2{$random}};
    wb_reg_wdata = {2{$random}};
    mem_reg_wdata = {2{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R98 = {2{$random}};
    R99 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    ex_reg_ctrl_fn_dw = {1{$random}};
    ex_reg_ctrl_fn_alu = {1{$random}};
    ex_reg_sel_alu1 = {1{$random}};
    ex_reg_sel_alu2 = {1{$random}};
    ex_reg_sel_imm = {1{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
  end
`endif

  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T7 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T6 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data : ex_reg_inst;
  assign T5 = io_ctrl_killd ^ 1'h1;
  assign T6 = ex_reg_kill ^ 1'h1;
  assign T7 = mem_reg_kill ^ 1'h1;
  assign T8 = wb_reg_inst;
  assign T9 = R10;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T87 : T12;
  assign T12 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T13 = T82 ? io_ctrl_bypass_src_1 : T14;
  assign T14 = T81 ? T15 : ex_reg_rs_lsb_1;
  assign T15 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T16;
  assign T16 = T79 ? wb_wdata : T17;
  assign T17 = T18[T26];
  assign T20 = T23 & T21;
  assign T21 = T22 < 5'h1f;
  assign T22 = T25[3'h4:1'h0];
  assign T23 = wb_wen & T24;
  assign T24 = wb_waddr != 5'h0;
  assign wb_waddr = io_ctrl_ll_wen ? io_ctrl_ll_waddr : io_ctrl_wb_waddr;
  assign wb_wen = io_ctrl_ll_wen | io_ctrl_wb_wen;
  assign T25 = ~ wb_waddr;
  assign T26 = ~ T27;
  assign T27 = io_imem_resp_bits_data[5'h18:5'h14];
  assign wb_wdata = T28;
  assign T28 = T76 ? io_dmem_resp_bits_data_subword : T29;
  assign T29 = io_ctrl_ll_wen ? ll_wdata : T30;
  assign T30 = T73 ? pcr_io_rw_rdata : wb_reg_wdata;
  assign T31 = T7 ? T32 : wb_reg_wdata;
  assign T32 = T72 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = io_ctrl_mem_jalr ? T205 : mem_reg_wdata;
  assign T33 = T6 ? alu_io_out : mem_reg_wdata;
  assign T205 = {T212, mem_br_target};
  assign mem_br_target = T206 + T34;
  assign T34 = T35;
  assign T35 = {1'h0, mem_reg_pc};
  assign T36 = T6 ? ex_reg_pc : mem_reg_pc;
  assign T37 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T206 = {T210, T38};
  assign T38 = T71 ? T207 : T39;
  assign T39 = T55 ? T40 : 22'h4;
  assign T40 = T41;
  assign T41 = {T49, T42};
  assign T42 = {T45, T43};
  assign T43 = {T44, 1'h0};
  assign T44 = mem_reg_inst[5'h18:5'h15];
  assign T45 = {T47, T46};
  assign T46 = mem_reg_inst[5'h1e:5'h19];
  assign T47 = T48;
  assign T48 = mem_reg_inst[5'h14:5'h14];
  assign T49 = {T53, T50};
  assign T50 = {T53, T51};
  assign T51 = T52;
  assign T52 = mem_reg_inst[5'h13:4'hc];
  assign T53 = T54;
  assign T54 = mem_reg_inst[5'h1f:5'h1f];
  assign T55 = T57 & T56;
  assign T56 = io_ctrl_mem_branch ^ 1'h1;
  assign T57 = io_ctrl_mem_jalr ^ 1'h1;
  assign T207 = {T208, T58};
  assign T58 = T59;
  assign T59 = {T67, T60};
  assign T60 = {T63, T61};
  assign T61 = {T62, 1'h0};
  assign T62 = mem_reg_inst[4'hb:4'h8];
  assign T63 = {T65, T64};
  assign T64 = mem_reg_inst[5'h1e:5'h19];
  assign T65 = T66;
  assign T66 = mem_reg_inst[3'h7:3'h7];
  assign T67 = {T69, T68};
  assign T68 = {T69, T69};
  assign T69 = T70;
  assign T70 = mem_reg_inst[5'h1f:5'h1f];
  assign T208 = T209 ? 7'h7f : 7'h0;
  assign T209 = T58[4'he:4'he];
  assign T71 = io_ctrl_mem_branch & io_ctrl_mem_br_taken;
  assign T210 = T211 ? 23'h7fffff : 23'h0;
  assign T211 = T38[5'h15:5'h15];
  assign T212 = T213 ? 19'h7ffff : 19'h0;
  assign T213 = mem_br_target[6'h2c:6'h2c];
  assign T72 = io_ctrl_mem_fp_val & io_ctrl_mem_wen;
  assign T73 = io_ctrl_csr != 3'h0;
  assign ll_wdata = T74;
  assign T74 = T75 ? io_rocc_resp_bits_data : div_io_resp_bits_data;
  assign T75 = io_rocc_resp_ready & io_rocc_resp_valid;
  assign T76 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_xpu = T77 ^ 1'h1;
  assign T77 = T78;
  assign T78 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T79 = T23 & T80;
  assign T80 = wb_waddr == T27;
  assign T81 = T5 & io_ctrl_ren_1;
  assign T82 = T5 & io_ctrl_bypass_1;
  assign T83 = T85 ? T84 : ex_reg_rs_msb_1;
  assign T84 = id_rs_1 >> 2'h2;
  assign T85 = T81 & T86;
  assign T86 = io_ctrl_bypass_1 ^ 1'h1;
  assign T87 = T93 ? T91 : T88;
  assign T88 = T89 ? bypass_1 : T214;
  assign T214 = {63'h0, bypass_0};
  assign bypass_0 = 1'h0;
  assign bypass_1 = mem_reg_wdata;
  assign T89 = T90[1'h0:1'h0];
  assign T90 = ex_reg_rs_lsb_1;
  assign T91 = T92 ? bypass_3 : bypass_2;
  assign bypass_2 = wb_reg_wdata;
  assign bypass_3 = io_dmem_resp_bits_data;
  assign T92 = T90[1'h0:1'h0];
  assign T93 = T90[1'h1:1'h1];
  assign T94 = T5 ? io_ctrl_bypass_1 : ex_reg_rs_bypass_1;
  assign T95 = T96;
  assign T96 = wb_reg_inst[5'h18:5'h14];
  assign T97 = R98;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T116 : T100;
  assign T100 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T101 = T111 ? io_ctrl_bypass_src_0 : T102;
  assign T102 = T110 ? T103 : ex_reg_rs_lsb_0;
  assign T103 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T104;
  assign T104 = T108 ? wb_wdata : T105;
  assign T105 = T18[T106];
  assign T106 = ~ T107;
  assign T107 = io_imem_resp_bits_data[5'h13:4'hf];
  assign T108 = T23 & T109;
  assign T109 = wb_waddr == T107;
  assign T110 = T5 & io_ctrl_ren_0;
  assign T111 = T5 & io_ctrl_bypass_0;
  assign T112 = T114 ? T113 : ex_reg_rs_msb_0;
  assign T113 = id_rs_0 >> 2'h2;
  assign T114 = T110 & T115;
  assign T115 = io_ctrl_bypass_0 ^ 1'h1;
  assign T116 = T122 ? T120 : T117;
  assign T117 = T118 ? bypass_1 : T215;
  assign T215 = {63'h0, bypass_0};
  assign T118 = T119[1'h0:1'h0];
  assign T119 = ex_reg_rs_lsb_0;
  assign T120 = T121 ? bypass_3 : bypass_2;
  assign T121 = T119[1'h0:1'h0];
  assign T122 = T119[1'h1:1'h1];
  assign T123 = T5 ? io_ctrl_bypass_0 : ex_reg_rs_bypass_0;
  assign T124 = T125;
  assign T125 = wb_reg_inst[5'h13:4'hf];
  assign T126 = wb_wen;
  assign T127 = wb_wdata;
  assign T128 = T129;
  assign T129 = wb_wen ? wb_waddr : 5'h0;
  assign T130 = wb_reg_pc;
  assign T131 = T7 ? mem_reg_pc : wb_reg_pc;
  assign T132 = io_ctrl_retire;
  assign T133 = T134;
  assign T134 = pcr_io_time[6'h20:1'h0];
  assign T135 = io_host_id;
  assign T228 = T234 ? T233 : T229;
  assign T229 = T232 ? T230 : wb_reg_wdata;
  assign T230 = pcr_io_rw_rdata & T231;
  assign T231 = ~ wb_reg_wdata;
  assign T232 = io_ctrl_csr == 3'h3;
  assign T233 = pcr_io_rw_rdata | wb_reg_wdata;
  assign T234 = io_ctrl_csr == 3'h2;
  assign T235 = io_ctrl_csr[1'h1:1'h0];
  assign T236 = wb_reg_inst[5'h1f:5'h14];
  assign T237 = T138 ? 1'h0 : T238;
  assign T238 = T75 ? 1'h0 : io_ctrl_ll_ready;
  assign T138 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T239 = T5 ? T240 : ex_reg_ctrl_fn_dw;
  assign T240 = io_ctrl_fn_dw;
  assign T241 = T5 ? io_ctrl_fn_alu : ex_reg_ctrl_fn_alu;
  assign ex_op1 = T250 ? T249 : T242;
  assign T242 = {T247, T243};
  assign T243 = T245 ? T244 : 44'h0;
  assign T244 = ex_reg_pc;
  assign T245 = ex_reg_sel_alu1 == 2'h2;
  assign T246 = T5 ? io_ctrl_sel_alu1 : ex_reg_sel_alu1;
  assign T247 = T248 ? 20'hfffff : 20'h0;
  assign T248 = T243[6'h2b:6'h2b];
  assign T249 = ex_rs_0;
  assign T250 = ex_reg_sel_alu1 == 2'h1;
  assign T251 = ex_op2;
  assign ex_op2 = T322 ? T321 : T252;
  assign T252 = {T319, T253};
  assign T253 = T318 ? ex_imm : T254;
  assign T254 = {T258, T255};
  assign T255 = T256 ? 4'h4 : 4'h0;
  assign T256 = ex_reg_sel_alu2 == 3'h1;
  assign T257 = T5 ? io_ctrl_sel_alu2 : ex_reg_sel_alu2;
  assign T258 = T259 ? 28'hfffffff : 28'h0;
  assign T259 = T255[2'h3:2'h3];
  assign ex_imm = T260;
  assign T260 = {T304, T261};
  assign T261 = {T284, T262};
  assign T262 = {T273, T263};
  assign T263 = T272 ? T271 : T264;
  assign T264 = T270 ? T269 : T265;
  assign T265 = T267 ? T266 : 1'h0;
  assign T266 = ex_reg_inst[4'hf:4'hf];
  assign T267 = ex_reg_sel_imm == 3'h5;
  assign T268 = T5 ? io_ctrl_sel_imm : ex_reg_sel_imm;
  assign T269 = ex_reg_inst[5'h14:5'h14];
  assign T270 = ex_reg_sel_imm == 3'h4;
  assign T271 = ex_reg_inst[3'h7:3'h7];
  assign T272 = ex_reg_sel_imm == 3'h0;
  assign T273 = T283 ? 4'h0 : T274;
  assign T274 = T280 ? T279 : T275;
  assign T275 = T278 ? T277 : T276;
  assign T276 = ex_reg_inst[5'h18:5'h15];
  assign T277 = ex_reg_inst[5'h13:5'h10];
  assign T278 = ex_reg_sel_imm == 3'h5;
  assign T279 = ex_reg_inst[4'hb:4'h8];
  assign T280 = T282 | T281;
  assign T281 = ex_reg_sel_imm == 3'h1;
  assign T282 = ex_reg_sel_imm == 3'h0;
  assign T283 = ex_reg_sel_imm == 3'h2;
  assign T284 = {T290, T285};
  assign T285 = T287 ? 6'h0 : T286;
  assign T286 = ex_reg_inst[5'h1e:5'h19];
  assign T287 = T289 | T288;
  assign T288 = ex_reg_sel_imm == 3'h5;
  assign T289 = ex_reg_sel_imm == 3'h2;
  assign T290 = T301 ? 1'h0 : T291;
  assign T291 = T300 ? T298 : T292;
  assign T292 = T297 ? T295 : T293;
  assign T293 = T294;
  assign T294 = ex_reg_inst[5'h1f:5'h1f];
  assign T295 = T296;
  assign T296 = ex_reg_inst[3'h7:3'h7];
  assign T297 = ex_reg_sel_imm == 3'h1;
  assign T298 = T299;
  assign T299 = ex_reg_inst[5'h14:5'h14];
  assign T300 = ex_reg_sel_imm == 3'h3;
  assign T301 = T303 | T302;
  assign T302 = ex_reg_sel_imm == 3'h5;
  assign T303 = ex_reg_sel_imm == 3'h2;
  assign T304 = {T293, T305};
  assign T305 = {T313, T306};
  assign T306 = T310 ? T309 : T307;
  assign T307 = T308;
  assign T308 = ex_reg_inst[5'h13:4'hc];
  assign T309 = T293 ? 8'hff : 8'h0;
  assign T310 = T312 & T311;
  assign T311 = ex_reg_sel_imm != 3'h3;
  assign T312 = ex_reg_sel_imm != 3'h2;
  assign T313 = T317 ? T315 : T314;
  assign T314 = T293 ? 11'h7ff : 11'h0;
  assign T315 = T316;
  assign T316 = ex_reg_inst[5'h1e:5'h14];
  assign T317 = ex_reg_sel_imm == 3'h2;
  assign T318 = ex_reg_sel_alu2 == 3'h3;
  assign T319 = T320 ? 32'hffffffff : 32'h0;
  assign T320 = T253[5'h1f:5'h1f];
  assign T321 = ex_rs_1;
  assign T322 = ex_reg_sel_alu2 == 3'h2;
  assign io_temac_sfp_tx_disable = pcr_io_temac_sfp_tx_disable;
  assign io_temac_s_axi_rready = pcr_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = pcr_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = pcr_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = pcr_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = pcr_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = pcr_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = pcr_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = pcr_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = pcr_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = pcr_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = pcr_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = pcr_io_temac_rx_axis_fifo_tready;
  assign io_rocc_resp_ready = T137;
  assign T137 = T138 ? 1'h0 : io_ctrl_ll_ready;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T139 = io_ctrl_mem_rocc_val ? mem_reg_rs2 : wb_reg_rs2;
  assign T140 = io_ctrl_ex_rs2_val ? ex_rs_1 : mem_reg_rs2;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_inst_opcode = T141;
  assign T141 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T142;
  assign T142 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T143;
  assign T143 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T144;
  assign T144 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T145;
  assign T145 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T146;
  assign T146 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T147;
  assign T147 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T148;
  assign T148 = wb_reg_inst[5'h1f:5'h19];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = T216;
  assign T216 = dmem_resp_waddr[3'h4:1'h0];
  assign dmem_resp_waddr = T149 >> 1'h1;
  assign T149 = io_dmem_resp_bits_tag;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T150;
  assign T150 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T151;
  assign T151 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = pcr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data;
  assign io_imem_btb_update_bits_returnAddr = T217;
  assign T217 = mem_int_wdata[6'h2a:1'h0];
  assign io_imem_btb_update_bits_target = T218;
  assign T218 = io_imem_req_bits_pc[6'h2a:1'h0];
  assign io_imem_btb_update_bits_pc = T219;
  assign T219 = mem_reg_pc[6'h2a:1'h0];
  assign io_imem_req_bits_pc = T220;
  assign T220 = T152[6'h2b:1'h0];
  assign T152 = T153;
  assign T153 = T171 ? mem_npc : T221;
  assign T221 = {1'h0, T154};
  assign T154 = T155 ? pcr_io_evec : wb_reg_pc;
  assign T155 = io_ctrl_sel_pc == 3'h3;
  assign mem_npc = io_ctrl_mem_jalr ? T222 : mem_br_target;
  assign T222 = {1'h0, T156};
  assign T156 = {T158, T157};
  assign T157 = mem_reg_wdata[6'h2a:1'h0];
  assign T158 = T168 ? T167 : T159;
  assign T159 = T163 ? T162 : T160;
  assign T160 = T161[1'h0:1'h0];
  assign T161 = mem_reg_wdata[6'h2b:6'h2a];
  assign T162 = T161 == 2'h3;
  assign T163 = T166 | T164;
  assign T164 = T165 == 22'h3ffffe;
  assign T165 = mem_reg_wdata >> 6'h2a;
  assign T166 = T165 == 22'h3fffff;
  assign T167 = T161 != 2'h0;
  assign T168 = T170 | T169;
  assign T169 = T165 == 22'h1;
  assign T170 = T165 == 22'h0;
  assign T171 = io_ctrl_sel_pc == 3'h1;
  assign io_ptw_status_s = pcr_io_status_s;
  assign io_ptw_status_ps = pcr_io_status_ps;
  assign io_ptw_status_ei = pcr_io_status_ei;
  assign io_ptw_status_pei = pcr_io_status_pei;
  assign io_ptw_status_ef = pcr_io_status_ef;
  assign io_ptw_status_u64 = pcr_io_status_u64;
  assign io_ptw_status_s64 = pcr_io_status_s64;
  assign io_ptw_status_vm = pcr_io_status_vm;
  assign io_ptw_status_er = pcr_io_status_er;
  assign io_ptw_status_zero = pcr_io_status_zero;
  assign io_ptw_status_im = pcr_io_status_im;
  assign io_ptw_status_ip = pcr_io_status_ip;
  assign io_ptw_sret = io_ctrl_sret;
  assign io_ptw_invalidate = pcr_io_fatc;
  assign io_ptw_ptbr = pcr_io_ptbr;
  assign io_dmem_req_bits_data = T172;
  assign T172 = io_ctrl_mem_fp_val ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_tag = T223;
  assign T223 = {3'h0, T173};
  assign T173 = {io_ctrl_ex_waddr, io_ctrl_ex_fp_val};
  assign io_dmem_req_bits_addr = T174;
  assign T174 = T175;
  assign T175 = {T177, T176};
  assign T176 = alu_io_adder_out[6'h2a:1'h0];
  assign T177 = T187 ? T186 : T178;
  assign T178 = T182 ? T181 : T179;
  assign T179 = T180[1'h0:1'h0];
  assign T180 = alu_io_adder_out[6'h2b:6'h2a];
  assign T181 = T180 == 2'h3;
  assign T182 = T185 | T183;
  assign T183 = T184 == 22'h3ffffe;
  assign T184 = ex_rs_0 >> 6'h2a;
  assign T185 = T184 == 22'h3fffff;
  assign T186 = T180 != 2'h0;
  assign T187 = T189 | T188;
  assign T188 = T184 == 22'h1;
  assign T189 = T184 == 22'h0;
  assign io_ctrl_csr_replay = pcr_io_replay;
  assign io_ctrl_fp_sboard_clra = T224;
  assign T224 = dmem_resp_waddr[3'h4:1'h0];
  assign io_ctrl_fp_sboard_clr = T190;
  assign T190 = dmem_resp_replay & dmem_resp_fpu;
  assign io_ctrl_status_s = pcr_io_status_s;
  assign io_ctrl_status_ps = pcr_io_status_ps;
  assign io_ctrl_status_ei = pcr_io_status_ei;
  assign io_ctrl_status_pei = pcr_io_status_pei;
  assign io_ctrl_status_ef = pcr_io_status_ef;
  assign io_ctrl_status_u64 = pcr_io_status_u64;
  assign io_ctrl_status_s64 = pcr_io_status_s64;
  assign io_ctrl_status_vm = pcr_io_status_vm;
  assign io_ctrl_status_er = pcr_io_status_er;
  assign io_ctrl_status_zero = pcr_io_status_zero;
  assign io_ctrl_status_im = pcr_io_status_im;
  assign io_ctrl_status_ip = pcr_io_status_ip;
  assign io_ctrl_wb_waddr = T191;
  assign T191 = wb_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_waddr = T192;
  assign T192 = mem_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_rs1_ra = T193;
  assign T193 = T194 == 5'h1;
  assign T194 = mem_reg_inst[5'h13:4'hf];
  assign io_ctrl_ex_waddr = T195;
  assign T195 = ex_reg_inst[4'hb:3'h7];
  assign io_ctrl_ll_waddr = T225;
  assign T225 = T196[3'h4:1'h0];
  assign T196 = T138 ? dmem_resp_waddr : T226;
  assign T226 = {3'h0, T197};
  assign T197 = T75 ? io_rocc_resp_bits_rd : div_io_resp_bits_tag;
  assign io_ctrl_ll_wen = T198;
  assign T198 = T138 ? 1'h1 : T199;
  assign T199 = T75 ? 1'h1 : T200;
  assign T200 = T237 & div_io_resp_valid;
  assign io_ctrl_div_mul_rdy = div_io_req_ready;
  assign io_ctrl_mem_misprediction = T201;
  assign T201 = T203 | T202;
  assign T202 = io_ctrl_ex_valid ^ 1'h1;
  assign T203 = mem_npc != T227;
  assign T227 = {1'h0, ex_reg_pc};
  assign io_ctrl_mem_br_taken = T204;
  assign T204 = mem_reg_wdata[1'h0:1'h0];
  assign io_ctrl_inst = io_imem_resp_bits_data;
  assign io_host_debug_stats_pcr = pcr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = pcr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = pcr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = pcr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = pcr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = pcr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = pcr_io_host_pcr_req_ready;
  ALU alu(
       .io_dw( ex_reg_ctrl_fn_dw ),
       .io_fn( ex_reg_ctrl_fn_alu ),
       .io_in2( T251 ),
       .io_in1( ex_op1 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( io_ctrl_div_mul_val ),
       .io_req_bits_fn( ex_reg_ctrl_fn_alu ),
       .io_req_bits_dw( ex_reg_ctrl_fn_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( io_ctrl_ex_waddr ),
       .io_kill( io_ctrl_div_mul_kill ),
       .io_resp_ready( T237 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );
  CSRFile pcr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( pcr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( pcr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( pcr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( pcr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( pcr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( pcr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( pcr_io_host_debug_stats_pcr ),
       .io_rw_addr( T236 ),
       .io_rw_cmd( T235 ),
       .io_rw_rdata( pcr_io_rw_rdata ),
       .io_rw_wdata( T228 ),
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( pcr_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( pcr_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( pcr_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( pcr_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( pcr_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( pcr_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( pcr_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( pcr_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( pcr_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( pcr_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( pcr_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( pcr_io_temac_s_axi_rready ),
       .io_temac_sfp_tx_disable( pcr_io_temac_sfp_tx_disable ),
       .io_status_ip( pcr_io_status_ip ),
       .io_status_im( pcr_io_status_im ),
       .io_status_zero( pcr_io_status_zero ),
       .io_status_er( pcr_io_status_er ),
       .io_status_vm( pcr_io_status_vm ),
       .io_status_s64( pcr_io_status_s64 ),
       .io_status_u64( pcr_io_status_u64 ),
       .io_status_ef( pcr_io_status_ef ),
       .io_status_pei( pcr_io_status_pei ),
       .io_status_ei( pcr_io_status_ei ),
       .io_status_ps( pcr_io_status_ps ),
       .io_status_s( pcr_io_status_s ),
       .io_ptbr( pcr_io_ptbr ),
       .io_evec( pcr_io_evec ),
       .io_exception( io_ctrl_exception ),
       .io_retire( io_ctrl_retire ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( io_ctrl_cause ),
       .io_badvaddr_wen( io_ctrl_badvaddr_wen ),
       .io_pc( wb_reg_pc ),
       .io_sret( io_ctrl_sret ),
       .io_fatc( pcr_io_fatc ),
       .io_replay( pcr_io_replay ),
       .io_time( pcr_io_time ),
       .io_fcsr_rm( pcr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );

  always @(posedge clk) begin
    if(T7) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T6) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data;
    end
    ex_reg_kill <= io_ctrl_killd;
    mem_reg_kill <= ex_reg_kill;
    R10 <= R11;
    if(ex_reg_rs_bypass_1) begin
      R11 <= T87;
    end else begin
      R11 <= T12;
    end
    if(T82) begin
      ex_reg_rs_lsb_1 <= io_ctrl_bypass_src_1;
    end else if(T81) begin
      ex_reg_rs_lsb_1 <= T15;
    end
    if (T20)
      T18[T25] <= wb_wdata;
    if(T7) begin
      wb_reg_wdata <= T32;
    end
    if(T6) begin
      mem_reg_wdata <= alu_io_out;
    end
    if(T6) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T85) begin
      ex_reg_rs_msb_1 <= T84;
    end
    if(T5) begin
      ex_reg_rs_bypass_1 <= io_ctrl_bypass_1;
    end
    R98 <= R99;
    if(ex_reg_rs_bypass_0) begin
      R99 <= T116;
    end else begin
      R99 <= T100;
    end
    if(T111) begin
      ex_reg_rs_lsb_0 <= io_ctrl_bypass_src_0;
    end else if(T110) begin
      ex_reg_rs_lsb_0 <= T103;
    end
    if(T114) begin
      ex_reg_rs_msb_0 <= T113;
    end
    if(T5) begin
      ex_reg_rs_bypass_0 <= io_ctrl_bypass_0;
    end
    if(T7) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if(T5) begin
      ex_reg_ctrl_fn_dw <= T240;
    end
    if(T5) begin
      ex_reg_ctrl_fn_alu <= io_ctrl_fn_alu;
    end
    if(T5) begin
      ex_reg_sel_alu1 <= io_ctrl_sel_alu1;
    end
    if(T5) begin
      ex_reg_sel_alu2 <= io_ctrl_sel_alu2;
    end
    if(T5) begin
      ex_reg_sel_imm <= io_ctrl_sel_imm;
    end
    if(io_ctrl_mem_rocc_val) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(io_ctrl_ex_rs2_val) begin
      mem_reg_rs2 <= ex_rs_1;
    end
`ifndef SYNTHESIS
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T135, T133, T132, T130, T128, T127, T126, T124, T97, T95, T9, T8, T1);
`endif
  end
endmodule

module FPUDecoder(
    input [31:0] io_inst,
    output[4:0] io_sigs_cmd,
    output io_sigs_ldst,
    output io_sigs_wen,
    output io_sigs_ren1,
    output io_sigs_ren2,
    output io_sigs_ren3,
    output io_sigs_swap23,
    output io_sigs_single,
    output io_sigs_fromint,
    output io_sigs_toint,
    output io_sigs_fastpipe,
    output io_sigs_fma,
    output io_sigs_round
);

  wire T0;
  wire T1;
  wire[31:0] T2;
  wire T3;
  wire T4;
  wire[31:0] T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  wire T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire T16;
  wire[31:0] T17;
  wire T18;
  wire T19;
  wire[31:0] T20;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire[31:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire T41;
  wire[31:0] T42;
  wire T43;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire[31:0] T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire[31:0] T55;
  wire T56;
  wire T57;
  wire[31:0] T58;
  wire T59;
  wire T60;
  wire[31:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[31:0] T65;
  wire T66;
  wire T67;
  wire[31:0] T68;
  wire T69;
  wire T70;
  wire[31:0] T71;
  wire T72;
  wire T73;
  wire[31:0] T74;
  wire T75;
  wire T76;
  wire[31:0] T77;
  wire T78;
  wire T79;
  wire[31:0] T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[31:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire[31:0] T114;
  wire[4:0] T115;
  wire[3:0] T116;
  wire[2:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire[31:0] T121;
  wire T122;
  wire[31:0] T123;
  wire T124;
  wire T125;
  wire[31:0] T126;
  wire T127;
  wire[31:0] T128;
  wire T129;
  wire T130;
  wire[31:0] T131;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire T135;
  wire[31:0] T136;
  wire T137;
  wire[31:0] T138;


  assign io_sigs_round = T0;
  assign T0 = T3 | T1;
  assign T1 = T2 == 32'he0000053;
  assign T2 = io_inst & 32'hedf0707f;
  assign T3 = T6 | T4;
  assign T4 = T5 == 32'he0000053;
  assign T5 = io_inst & 32'hfdf0607f;
  assign T6 = T9 | T7;
  assign T7 = T8 == 32'hc0000053;
  assign T8 = io_inst & 32'hedc0007f;
  assign T9 = T12 | T10;
  assign T10 = T11 == 32'h42000053;
  assign T11 = io_inst & 32'h7ff0007f;
  assign T12 = T15 | T13;
  assign T13 = T14 == 32'h40100053;
  assign T14 = io_inst & 32'h7ff0007f;
  assign T15 = T18 | T16;
  assign T16 = T17 == 32'h53;
  assign T17 = io_inst & 32'hec00007f;
  assign T18 = T21 | T19;
  assign T19 = T20 == 32'h53;
  assign T20 = io_inst & 32'hf400007f;
  assign T21 = T22 == 32'h43;
  assign T22 = io_inst & 32'h4000073;
  assign io_sigs_fma = T23;
  assign T23 = T24 | T16;
  assign T24 = T21 | T19;
  assign io_sigs_fastpipe = T25;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h42000053;
  assign T27 = io_inst & 32'hfff0007f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h40100053;
  assign T30 = io_inst & 32'hfff0007f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h20000053;
  assign T33 = io_inst & 32'hf400607f;
  assign T34 = T35 == 32'h20000053;
  assign T35 = io_inst & 32'hfc00507f;
  assign io_sigs_toint = T36;
  assign T36 = T37 | T4;
  assign T37 = T40 | T38;
  assign T38 = T39 == 32'hc0000053;
  assign T39 = io_inst & 32'hfdc0007f;
  assign T40 = T43 | T41;
  assign T41 = T42 == 32'ha0000053;
  assign T42 = io_inst & 32'hfc00507f;
  assign T43 = T46 | T44;
  assign T44 = T45 == 32'ha0000053;
  assign T45 = io_inst & 32'hfc00607f;
  assign T46 = T47 == 32'h2027;
  assign T47 = io_inst & 32'h607f;
  assign io_sigs_fromint = T48;
  assign T48 = T51 | T49;
  assign T49 = T50 == 32'hf0000053;
  assign T50 = io_inst & 32'hfdf0707f;
  assign T51 = T52 == 32'hd0000053;
  assign T52 = io_inst & 32'hfdc0007f;
  assign io_sigs_single = T53;
  assign T53 = T56 | T54;
  assign T54 = T55 == 32'he0000053;
  assign T55 = io_inst & 32'heff0707f;
  assign T56 = T59 | T57;
  assign T57 = T58 == 32'he0000053;
  assign T58 = io_inst & 32'hfff0607f;
  assign T59 = T62 | T60;
  assign T60 = T61 == 32'hc0000053;
  assign T61 = io_inst & 32'hefc0007f;
  assign T62 = T63 | T13;
  assign T63 = T66 | T64;
  assign T64 = T65 == 32'h20000053;
  assign T65 = io_inst & 32'h7e00507f;
  assign T66 = T69 | T67;
  assign T67 = T68 == 32'h20000053;
  assign T68 = io_inst & 32'h7e00607f;
  assign T69 = T72 | T70;
  assign T70 = T71 == 32'h20000053;
  assign T71 = io_inst & 32'hf600607f;
  assign T72 = T75 | T73;
  assign T73 = T74 == 32'h2007;
  assign T74 = io_inst & 32'h705f;
  assign T75 = T78 | T76;
  assign T76 = T77 == 32'h53;
  assign T77 = io_inst & 32'hee00007f;
  assign T78 = T81 | T79;
  assign T79 = T80 == 32'h53;
  assign T80 = io_inst & 32'hf600007f;
  assign T81 = T82 == 32'h43;
  assign T82 = io_inst & 32'h6000073;
  assign io_sigs_swap23 = T19;
  assign io_sigs_ren3 = T21;
  assign io_sigs_ren2 = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h20000053;
  assign T85 = io_inst & 32'h7c00507f;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h20000053;
  assign T88 = io_inst & 32'h7c00607f;
  assign T89 = T90 | T32;
  assign T90 = T91 | T46;
  assign T91 = T92 | T16;
  assign T92 = T21 | T19;
  assign io_sigs_ren1 = T93;
  assign T93 = T94 | T4;
  assign T94 = T95 | T38;
  assign T95 = T96 | T10;
  assign T96 = T97 | T13;
  assign T97 = T98 | T84;
  assign T98 = T99 | T87;
  assign T99 = T100 | T32;
  assign T100 = T101 | T16;
  assign T101 = T21 | T19;
  assign io_sigs_wen = T102;
  assign T102 = T103 | T49;
  assign T103 = T104 | T51;
  assign T104 = T105 | T26;
  assign T105 = T106 | T29;
  assign T106 = T107 | T32;
  assign T107 = T108 | T34;
  assign T108 = T111 | T109;
  assign T109 = T110 == 32'h2007;
  assign T110 = io_inst & 32'h607f;
  assign T111 = T112 | T16;
  assign T112 = T21 | T19;
  assign io_sigs_ldst = T113;
  assign T113 = T114 == 32'h2007;
  assign T114 = io_inst & 32'h605f;
  assign io_sigs_cmd = T115;
  assign T115 = {T137, T116};
  assign T116 = {T134, T117};
  assign T117 = {T129, T118};
  assign T118 = {T124, T119};
  assign T119 = T122 | T120;
  assign T120 = T121 == 32'h8000010;
  assign T121 = io_inst & 32'h8000010;
  assign T122 = T123 == 32'h4;
  assign T123 = io_inst & 32'h4;
  assign T124 = T127 | T125;
  assign T125 = T126 == 32'h10000010;
  assign T126 = io_inst & 32'h10000010;
  assign T127 = T128 == 32'h8;
  assign T128 = io_inst & 32'h8;
  assign T129 = T132 | T130;
  assign T130 = T131 == 32'h20000000;
  assign T131 = io_inst & 32'h20000000;
  assign T132 = T133 == 32'h0;
  assign T133 = io_inst & 32'h40;
  assign T134 = T132 | T135;
  assign T135 = T136 == 32'h40000000;
  assign T136 = io_inst & 32'h40000000;
  assign T137 = T138 == 32'h0;
  assign T138 = io_inst & 32'h10;
endmodule

module mulAddSubRecodedFloatN_0(
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[27:0] T4;
  wire[27:0] T529;
  wire[25:0] T5;
  wire[26:0] roundMask;
  wire[26:0] T6;
  wire[24:0] T7;
  wire[24:0] T530;
  wire T8;
  wire[24:0] T9;
  wire[8:0] T10;
  wire T11;
  wire[8:0] T12;
  wire[24:0] T13;
  wire[1024:0] T14;
  wire[9:0] T15;
  wire[9:0] sExpX3_13;
  wire[10:0] sExpX3;
  wire[10:0] T531;
  wire[6:0] estNormDist;
  wire[6:0] T16;
  wire[6:0] estNormNeg_dist;
  wire[6:0] T17;
  wire[6:0] T18;
  wire[6:0] T19;
  wire[6:0] T20;
  wire[6:0] T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[6:0] T24;
  wire[6:0] T25;
  wire[6:0] T26;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[6:0] T29;
  wire[6:0] T30;
  wire[6:0] T31;
  wire[6:0] T32;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[6:0] T40;
  wire[6:0] T41;
  wire[6:0] T42;
  wire[6:0] T43;
  wire[6:0] T44;
  wire[6:0] T45;
  wire[6:0] T46;
  wire[6:0] T47;
  wire[6:0] T48;
  wire[6:0] T49;
  wire[6:0] T50;
  wire[6:0] T51;
  wire[6:0] T52;
  wire[6:0] T53;
  wire[6:0] T54;
  wire[6:0] T55;
  wire[6:0] T56;
  wire[6:0] T57;
  wire[6:0] T58;
  wire[6:0] T59;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire T65;
  wire[50:0] T66;
  wire[50:0] T67;
  wire[49:0] T68;
  wire[49:0] T69;
  wire[74:0] sigSum;
  wire[74:0] alignedNegSigC;
  wire[75:0] T70;
  wire T71;
  wire doSubMags;
  wire opSignC;
  wire T72;
  wire T73;
  wire signProd;
  wire T74;
  wire T75;
  wire signB;
  wire signA;
  wire T76;
  wire[23:0] T77;
  wire[23:0] CExtraMask;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[6:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[5:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[3:0] T89;
  wire[7:0] T90;
  wire[23:0] T91;
  wire[128:0] T92;
  wire[6:0] CAlignDist;
  wire[10:0] T93;
  wire[10:0] T94;
  wire[10:0] sNatCAlignDist;
  wire[10:0] T532;
  wire[8:0] expC;
  wire[10:0] sExpAlignedProd;
  wire[10:0] T95;
  wire[10:0] T533;
  wire[8:0] expA;
  wire[10:0] T96;
  wire[7:0] T97;
  wire[8:0] expB;
  wire[2:0] T98;
  wire[2:0] T534;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire CAlignDist_floor;
  wire T103;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T104;
  wire isZeroA;
  wire[2:0] T105;
  wire[7:0] T106;
  wire[7:0] T535;
  wire[3:0] T107;
  wire[7:0] T108;
  wire[7:0] T536;
  wire[5:0] T109;
  wire[7:0] T110;
  wire[7:0] T537;
  wire[6:0] T111;
  wire[15:0] T112;
  wire[15:0] T113;
  wire[15:0] T114;
  wire[14:0] T115;
  wire[15:0] T116;
  wire[15:0] T117;
  wire[15:0] T118;
  wire[13:0] T119;
  wire[15:0] T120;
  wire[15:0] T121;
  wire[15:0] T122;
  wire[11:0] T123;
  wire[15:0] T124;
  wire[15:0] T125;
  wire[15:0] T126;
  wire[7:0] T127;
  wire[15:0] T128;
  wire[15:0] T129;
  wire[15:0] T538;
  wire[7:0] T130;
  wire[15:0] T131;
  wire[15:0] T539;
  wire[11:0] T132;
  wire[15:0] T133;
  wire[15:0] T540;
  wire[13:0] T134;
  wire[15:0] T135;
  wire[15:0] T541;
  wire[14:0] T136;
  wire[23:0] sigC;
  wire[22:0] fractC;
  wire T137;
  wire isZeroC;
  wire[2:0] T138;
  wire[74:0] T139;
  wire[74:0] T140;
  wire[74:0] T141;
  wire[73:0] T142;
  wire[49:0] T143;
  wire[49:0] T542;
  wire[23:0] negSigC;
  wire[23:0] T144;
  wire[74:0] T543;
  wire[48:0] T145;
  wire[47:0] T146;
  wire[23:0] sigB;
  wire[22:0] fractB;
  wire T147;
  wire[23:0] sigA;
  wire[22:0] fractA;
  wire T148;
  wire[50:0] T544;
  wire[49:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire notCDom_signSigSum;
  wire[6:0] CDom_estNormDist;
  wire[6:0] T545;
  wire[4:0] T198;
  wire[6:0] T199;
  wire T200;
  wire CAlignDist_0;
  wire T201;
  wire[9:0] T202;
  wire isCDominant;
  wire T203;
  wire T204;
  wire[9:0] T205;
  wire T206;
  wire[10:0] sExpSum;
  wire[10:0] T546;
  wire[7:0] T207;
  wire[7:0] T208;
  wire[7:0] T209;
  wire[6:0] T210;
  wire[7:0] T211;
  wire[7:0] T212;
  wire[7:0] T213;
  wire[5:0] T214;
  wire[7:0] T215;
  wire[7:0] T216;
  wire[7:0] T217;
  wire[3:0] T218;
  wire[7:0] T219;
  wire[7:0] T220;
  wire[7:0] T547;
  wire[3:0] T221;
  wire[7:0] T222;
  wire[7:0] T548;
  wire[5:0] T223;
  wire[7:0] T224;
  wire[7:0] T549;
  wire[6:0] T225;
  wire[15:0] T226;
  wire[15:0] T227;
  wire[15:0] T228;
  wire[14:0] T229;
  wire[15:0] T230;
  wire[15:0] T231;
  wire[15:0] T232;
  wire[13:0] T233;
  wire[15:0] T234;
  wire[15:0] T235;
  wire[15:0] T236;
  wire[11:0] T237;
  wire[15:0] T238;
  wire[15:0] T239;
  wire[15:0] T240;
  wire[7:0] T241;
  wire[15:0] T242;
  wire[15:0] T243;
  wire[15:0] T550;
  wire[7:0] T244;
  wire[15:0] T245;
  wire[15:0] T551;
  wire[11:0] T246;
  wire[15:0] T247;
  wire[15:0] T552;
  wire[13:0] T248;
  wire[15:0] T249;
  wire[15:0] T553;
  wire[14:0] T250;
  wire[26:0] T251;
  wire[26:0] T554;
  wire T252;
  wire[27:0] sigX3;
  wire[42:0] T253;
  wire T254;
  wire T255;
  wire[15:0] T256;
  wire[15:0] absSigSumExtraMask;
  wire[14:0] T257;
  wire[6:0] T258;
  wire[2:0] T259;
  wire T260;
  wire[2:0] T261;
  wire[6:0] T262;
  wire[14:0] T263;
  wire[16:0] T264;
  wire[3:0] normTo2ShiftDist;
  wire[3:0] estNormDist_5;
  wire[3:0] T265;
  wire[1:0] T266;
  wire T267;
  wire[1:0] T268;
  wire T269;
  wire[3:0] T270;
  wire[1:0] T271;
  wire T272;
  wire[1:0] T273;
  wire[3:0] T274;
  wire T275;
  wire[1:0] T276;
  wire T277;
  wire[1:0] T278;
  wire T279;
  wire[7:0] T280;
  wire[7:0] T281;
  wire[7:0] T282;
  wire[6:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[7:0] T286;
  wire[5:0] T287;
  wire[7:0] T288;
  wire[7:0] T289;
  wire[7:0] T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T293;
  wire[7:0] T555;
  wire[3:0] T294;
  wire[7:0] T295;
  wire[7:0] T556;
  wire[5:0] T296;
  wire[7:0] T297;
  wire[7:0] T557;
  wire[6:0] T298;
  wire[15:0] T299;
  wire[42:0] cFirstNormAbsSigSum;
  wire[42:0] T558;
  wire[41:0] T300;
  wire[41:0] notCDom_pos_firstNormAbsSigSum;
  wire[41:0] T301;
  wire[41:0] T302;
  wire[31:0] T303;
  wire[31:0] T559;
  wire[9:0] T304;
  wire[41:0] T560;
  wire[33:0] T305;
  wire T306;
  wire T307;
  wire[1:0] firstReduceSigSum;
  wire T308;
  wire[17:0] T309;
  wire T310;
  wire[15:0] T311;
  wire T312;
  wire T313;
  wire[1:0] firstReduceNotSigSum;
  wire T314;
  wire[17:0] T315;
  wire[74:0] notSigSum;
  wire T316;
  wire[15:0] T317;
  wire[32:0] T318;
  wire T319;
  wire[41:0] T320;
  wire[41:0] T321;
  wire[41:0] T322;
  wire[15:0] T323;
  wire[15:0] T561;
  wire[25:0] T324;
  wire T325;
  wire T326;
  wire[41:0] CDom_firstNormAbsSigSum;
  wire[41:0] T327;
  wire[41:0] T328;
  wire[41:0] T329;
  wire T330;
  wire[40:0] T331;
  wire[41:0] T562;
  wire T332;
  wire T333;
  wire T334;
  wire[41:0] T335;
  wire[41:0] T336;
  wire[41:0] T337;
  wire T338;
  wire[40:0] T339;
  wire[41:0] T563;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[41:0] T344;
  wire[41:0] T345;
  wire[41:0] T346;
  wire T347;
  wire[40:0] T348;
  wire[41:0] T564;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire[41:0] T353;
  wire[41:0] T354;
  wire T355;
  wire[40:0] T356;
  wire[41:0] T565;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire[42:0] T362;
  wire[42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[42:0] T363;
  wire[42:0] T364;
  wire[10:0] T365;
  wire[42:0] T566;
  wire[32:0] T366;
  wire T367;
  wire[31:0] T368;
  wire T369;
  wire[42:0] T370;
  wire[42:0] T567;
  wire[41:0] T371;
  wire[42:0] T372;
  wire[26:0] T373;
  wire T374;
  wire T375;
  wire[42:0] T568;
  wire T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[41:0] T380;
  wire[41:0] T381;
  wire roundPosBit;
  wire[27:0] T382;
  wire[27:0] T569;
  wire[26:0] roundPosMask;
  wire[26:0] T570;
  wire[25:0] T383;
  wire[25:0] T384;
  wire T385;
  wire allRound;
  wire allRoundExtra;
  wire[27:0] T386;
  wire[27:0] T571;
  wire[25:0] T387;
  wire[27:0] T388;
  wire doIncrSig;
  wire T389;
  wire T390;
  wire T391;
  wire commonCase;
  wire T392;
  wire notSpecial_addZeros;
  wire T393;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T394;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T395;
  wire isSpecialA;
  wire[1:0] T396;
  wire underflow;
  wire underflowY;
  wire T397;
  wire T398;
  wire[9:0] T572;
  wire[7:0] T399;
  wire sigX3Shift1;
  wire[1:0] T400;
  wire T401;
  wire overflow;
  wire overflowY;
  wire[2:0] T402;
  wire[10:0] sExpY;
  wire[10:0] T403;
  wire[10:0] T404;
  wire T405;
  wire[1:0] T406;
  wire[25:0] sigY3;
  wire[25:0] T407;
  wire[25:0] T408;
  wire[25:0] T409;
  wire[25:0] T410;
  wire[25:0] roundUp_sigY3;
  wire[25:0] T411;
  wire[25:0] T412;
  wire[27:0] T413;
  wire[27:0] T573;
  wire roundEven;
  wire T414;
  wire T415;
  wire T416;
  wire roundingMode_nearest_even;
  wire T417;
  wire T418;
  wire T419;
  wire[25:0] T420;
  wire[25:0] T421;
  wire roundUp;
  wire T422;
  wire T423;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T424;
  wire doNegSignSum;
  wire T425;
  wire T426;
  wire T427;
  wire isZeroY;
  wire[2:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire[25:0] T442;
  wire[25:0] T443;
  wire[27:0] T444;
  wire[27:0] T574;
  wire[26:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[10:0] T449;
  wire[10:0] T450;
  wire T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire[1:0] T455;
  wire invalid;
  wire notSigNaN_invalid;
  wire T456;
  wire T457;
  wire isInfC;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire isInfB;
  wire T462;
  wire T463;
  wire isInfA;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire isNaNB;
  wire T468;
  wire T469;
  wire isNaNA;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire isSigNaNC;
  wire T475;
  wire T476;
  wire isNaNC;
  wire T477;
  wire T478;
  wire isSigNaNB;
  wire T479;
  wire T480;
  wire isSigNaNA;
  wire T481;
  wire T482;
  wire[32:0] T483;
  wire[31:0] T484;
  wire[22:0] fractOut;
  wire[22:0] T485;
  wire[22:0] T575;
  wire T486;
  wire isSatOut;
  wire T487;
  wire overflowY_roundMagUp;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire isNaNOut;
  wire T492;
  wire T493;
  wire[22:0] fractY;
  wire[22:0] T494;
  wire[22:0] T495;
  wire[8:0] expOut;
  wire[8:0] T496;
  wire[8:0] T497;
  wire[8:0] T498;
  wire notNaN_isInfOut;
  wire T499;
  wire T500;
  wire T501;
  wire[8:0] T502;
  wire[8:0] T503;
  wire[8:0] T504;
  wire[8:0] T505;
  wire[8:0] T506;
  wire[8:0] T507;
  wire[8:0] T508;
  wire[8:0] T509;
  wire[8:0] T510;
  wire[8:0] T511;
  wire[8:0] T512;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T513;
  wire[8:0] T514;
  wire T515;
  wire T516;
  wire[8:0] expY;
  wire signOut;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;


  assign io_exceptionFlags = T0;
  assign T0 = {T455, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T385 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 28'h0;
  assign T4 = sigX3 & T529;
  assign T529 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T251 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T530;
  assign T530 = {24'h0, T8};
  assign T8 = sigX3[5'h1a:5'h1a];
  assign T9 = {T226, T10};
  assign T10 = {T207, T11};
  assign T11 = T12[4'h8:4'h8];
  assign T12 = T13[5'h18:5'h10];
  assign T13 = T14[8'h83:7'h6b];
  assign T14 = $signed(1025'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T15;
  assign T15 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'h9:1'h0];
  assign sExpX3 = sExpSum - T531;
  assign T531 = {4'h0, estNormDist};
  assign estNormDist = isCDominant ? CDom_estNormDist : T16;
  assign T16 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = T197 ? 7'h18 : T17;
  assign T17 = T196 ? 7'h19 : T18;
  assign T18 = T195 ? 7'h1a : T19;
  assign T19 = T194 ? 7'h1b : T20;
  assign T20 = T193 ? 7'h1c : T21;
  assign T21 = T192 ? 7'h1d : T22;
  assign T22 = T191 ? 7'h1e : T23;
  assign T23 = T190 ? 7'h1f : T24;
  assign T24 = T189 ? 7'h20 : T25;
  assign T25 = T188 ? 7'h21 : T26;
  assign T26 = T187 ? 7'h22 : T27;
  assign T27 = T186 ? 7'h23 : T28;
  assign T28 = T185 ? 7'h24 : T29;
  assign T29 = T184 ? 7'h25 : T30;
  assign T30 = T183 ? 7'h26 : T31;
  assign T31 = T182 ? 7'h27 : T32;
  assign T32 = T181 ? 7'h28 : T33;
  assign T33 = T180 ? 7'h29 : T34;
  assign T34 = T179 ? 7'h2a : T35;
  assign T35 = T178 ? 7'h2b : T36;
  assign T36 = T177 ? 7'h2c : T37;
  assign T37 = T176 ? 7'h2d : T38;
  assign T38 = T175 ? 7'h2e : T39;
  assign T39 = T174 ? 7'h2f : T40;
  assign T40 = T173 ? 7'h30 : T41;
  assign T41 = T172 ? 7'h31 : T42;
  assign T42 = T171 ? 7'h32 : T43;
  assign T43 = T170 ? 7'h33 : T44;
  assign T44 = T169 ? 7'h34 : T45;
  assign T45 = T168 ? 7'h35 : T46;
  assign T46 = T167 ? 7'h36 : T47;
  assign T47 = T166 ? 7'h37 : T48;
  assign T48 = T165 ? 7'h38 : T49;
  assign T49 = T164 ? 7'h39 : T50;
  assign T50 = T163 ? 7'h3a : T51;
  assign T51 = T162 ? 7'h3b : T52;
  assign T52 = T161 ? 7'h3c : T53;
  assign T53 = T160 ? 7'h3d : T54;
  assign T54 = T159 ? 7'h3e : T55;
  assign T55 = T158 ? 7'h3f : T56;
  assign T56 = T157 ? 7'h40 : T57;
  assign T57 = T156 ? 7'h41 : T58;
  assign T58 = T155 ? 7'h42 : T59;
  assign T59 = T154 ? 7'h43 : T60;
  assign T60 = T153 ? 7'h44 : T61;
  assign T61 = T152 ? 7'h45 : T62;
  assign T62 = T151 ? 7'h46 : T63;
  assign T63 = T150 ? 7'h47 : T64;
  assign T64 = T65 ? 7'h48 : 7'h49;
  assign T65 = T66[1'h1:1'h1];
  assign T66 = T544 ^ T67;
  assign T67 = T68 << 1'h1;
  assign T68 = 50'h0 | T69;
  assign T69 = sigSum[6'h32:1'h1];
  assign sigSum = T543 + alignedNegSigC;
  assign alignedNegSigC = T70[7'h4a:1'h0];
  assign T70 = {T139, T71};
  assign T71 = T76 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T73 ^ T72;
  assign T72 = io_op[1'h0:1'h0];
  assign T73 = io_c[6'h20:6'h20];
  assign signProd = T75 ^ T74;
  assign T74 = io_op[1'h1:1'h1];
  assign T75 = signA ^ signB;
  assign signB = io_b[6'h20:6'h20];
  assign signA = io_a[6'h20:6'h20];
  assign T76 = T77 != 24'h0;
  assign T77 = sigC & CExtraMask;
  assign CExtraMask = {T112, T78};
  assign T78 = T110 | T79;
  assign T79 = T80 & 8'haa;
  assign T80 = T81 << 1'h1;
  assign T81 = T82[3'h6:1'h0];
  assign T82 = T108 | T83;
  assign T83 = T84 & 8'hcc;
  assign T84 = T85 << 2'h2;
  assign T85 = T86[3'h5:1'h0];
  assign T86 = T106 | T87;
  assign T87 = T88 & 8'hf0;
  assign T88 = T89 << 3'h4;
  assign T89 = T90[2'h3:1'h0];
  assign T90 = T91[5'h17:5'h10];
  assign T91 = T92[7'h4d:6'h36];
  assign T92 = $signed(129'h100000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = T93[3'h6:1'h0];
  assign T93 = CAlignDist_floor ? 11'h0 : T94;
  assign T94 = T101 ? sNatCAlignDist : 11'h4a;
  assign sNatCAlignDist = sExpAlignedProd - T532;
  assign T532 = {2'h0, expC};
  assign expC = io_c[5'h1f:5'h17];
  assign sExpAlignedProd = T95 + 11'h1b;
  assign T95 = T96 + T533;
  assign T533 = {2'h0, expA};
  assign expA = io_a[5'h1f:5'h17];
  assign T96 = {T98, T97};
  assign T97 = expB[3'h7:1'h0];
  assign expB = io_b[5'h1f:5'h17];
  assign T98 = 3'h0 - T534;
  assign T534 = {2'h0, T99};
  assign T99 = T100 ^ 1'h1;
  assign T100 = expB[4'h8:4'h8];
  assign T101 = T102 < 10'h4a;
  assign T102 = sNatCAlignDist[4'h9:1'h0];
  assign CAlignDist_floor = isZeroProd | T103;
  assign T103 = sNatCAlignDist[4'ha:4'ha];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T104 == 3'h0;
  assign T104 = expB[4'h8:3'h6];
  assign isZeroA = T105 == 3'h0;
  assign T105 = expA[4'h8:3'h6];
  assign T106 = T535 & 8'hf;
  assign T535 = {4'h0, T107};
  assign T107 = T90 >> 3'h4;
  assign T108 = T536 & 8'h33;
  assign T536 = {2'h0, T109};
  assign T109 = T86 >> 2'h2;
  assign T110 = T537 & 8'h55;
  assign T537 = {1'h0, T111};
  assign T111 = T82 >> 1'h1;
  assign T112 = T135 | T113;
  assign T113 = T114 & 16'haaaa;
  assign T114 = T115 << 1'h1;
  assign T115 = T116[4'he:1'h0];
  assign T116 = T133 | T117;
  assign T117 = T118 & 16'hcccc;
  assign T118 = T119 << 2'h2;
  assign T119 = T120[4'hd:1'h0];
  assign T120 = T131 | T121;
  assign T121 = T122 & 16'hf0f0;
  assign T122 = T123 << 3'h4;
  assign T123 = T124[4'hb:1'h0];
  assign T124 = T129 | T125;
  assign T125 = T126 & 16'hff00;
  assign T126 = T127 << 4'h8;
  assign T127 = T128[3'h7:1'h0];
  assign T128 = T91[4'hf:1'h0];
  assign T129 = T538 & 16'hff;
  assign T538 = {8'h0, T130};
  assign T130 = T128 >> 4'h8;
  assign T131 = T539 & 16'hf0f;
  assign T539 = {4'h0, T132};
  assign T132 = T124 >> 3'h4;
  assign T133 = T540 & 16'h3333;
  assign T540 = {2'h0, T134};
  assign T134 = T120 >> 2'h2;
  assign T135 = T541 & 16'h5555;
  assign T541 = {1'h0, T136};
  assign T136 = T116 >> 1'h1;
  assign sigC = {T137, fractC};
  assign fractC = io_c[5'h16:1'h0];
  assign T137 = isZeroC ^ 1'h1;
  assign isZeroC = T138 == 3'h0;
  assign T138 = expC[4'h8:3'h6];
  assign T139 = $signed(T140) >>> CAlignDist;
  assign T140 = T141;
  assign T141 = {doSubMags, T142};
  assign T142 = {negSigC, T143};
  assign T143 = 50'h0 - T542;
  assign T542 = {49'h0, doSubMags};
  assign negSigC = doSubMags ? T144 : sigC;
  assign T144 = ~ sigC;
  assign T543 = {26'h0, T145};
  assign T145 = T146 << 1'h1;
  assign T146 = sigA * sigB;
  assign sigB = {T147, fractB};
  assign fractB = io_b[5'h16:1'h0];
  assign T147 = isZeroB ^ 1'h1;
  assign sigA = {T148, fractA};
  assign fractA = io_a[5'h16:1'h0];
  assign T148 = isZeroA ^ 1'h1;
  assign T544 = {1'h0, T149};
  assign T149 = 50'h0 ^ T69;
  assign T150 = T66[2'h2:2'h2];
  assign T151 = T66[2'h3:2'h3];
  assign T152 = T66[3'h4:3'h4];
  assign T153 = T66[3'h5:3'h5];
  assign T154 = T66[3'h6:3'h6];
  assign T155 = T66[3'h7:3'h7];
  assign T156 = T66[4'h8:4'h8];
  assign T157 = T66[4'h9:4'h9];
  assign T158 = T66[4'ha:4'ha];
  assign T159 = T66[4'hb:4'hb];
  assign T160 = T66[4'hc:4'hc];
  assign T161 = T66[4'hd:4'hd];
  assign T162 = T66[4'he:4'he];
  assign T163 = T66[4'hf:4'hf];
  assign T164 = T66[5'h10:5'h10];
  assign T165 = T66[5'h11:5'h11];
  assign T166 = T66[5'h12:5'h12];
  assign T167 = T66[5'h13:5'h13];
  assign T168 = T66[5'h14:5'h14];
  assign T169 = T66[5'h15:5'h15];
  assign T170 = T66[5'h16:5'h16];
  assign T171 = T66[5'h17:5'h17];
  assign T172 = T66[5'h18:5'h18];
  assign T173 = T66[5'h19:5'h19];
  assign T174 = T66[5'h1a:5'h1a];
  assign T175 = T66[5'h1b:5'h1b];
  assign T176 = T66[5'h1c:5'h1c];
  assign T177 = T66[5'h1d:5'h1d];
  assign T178 = T66[5'h1e:5'h1e];
  assign T179 = T66[5'h1f:5'h1f];
  assign T180 = T66[6'h20:6'h20];
  assign T181 = T66[6'h21:6'h21];
  assign T182 = T66[6'h22:6'h22];
  assign T183 = T66[6'h23:6'h23];
  assign T184 = T66[6'h24:6'h24];
  assign T185 = T66[6'h25:6'h25];
  assign T186 = T66[6'h26:6'h26];
  assign T187 = T66[6'h27:6'h27];
  assign T188 = T66[6'h28:6'h28];
  assign T189 = T66[6'h29:6'h29];
  assign T190 = T66[6'h2a:6'h2a];
  assign T191 = T66[6'h2b:6'h2b];
  assign T192 = T66[6'h2c:6'h2c];
  assign T193 = T66[6'h2d:6'h2d];
  assign T194 = T66[6'h2e:6'h2e];
  assign T195 = T66[6'h2f:6'h2f];
  assign T196 = T66[6'h30:6'h30];
  assign T197 = T66[6'h31:6'h31];
  assign notCDom_signSigSum = sigSum[6'h33:6'h33];
  assign CDom_estNormDist = T200 ? CAlignDist : T545;
  assign T545 = {2'h0, T198};
  assign T198 = T199[3'h4:1'h0];
  assign T199 = CAlignDist - 7'h1;
  assign T200 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T201;
  assign T201 = T202 == 10'h0;
  assign T202 = sNatCAlignDist[4'h9:1'h0];
  assign isCDominant = T206 & T203;
  assign T203 = CAlignDist_floor | T204;
  assign T204 = T205 < 10'h19;
  assign T205 = sNatCAlignDist[4'h9:1'h0];
  assign T206 = isZeroC ^ 1'h1;
  assign sExpSum = CAlignDist_floor ? T546 : sExpAlignedProd;
  assign T546 = {2'h0, expC};
  assign T207 = T224 | T208;
  assign T208 = T209 & 8'haa;
  assign T209 = T210 << 1'h1;
  assign T210 = T211[3'h6:1'h0];
  assign T211 = T222 | T212;
  assign T212 = T213 & 8'hcc;
  assign T213 = T214 << 2'h2;
  assign T214 = T215[3'h5:1'h0];
  assign T215 = T220 | T216;
  assign T216 = T217 & 8'hf0;
  assign T217 = T218 << 3'h4;
  assign T218 = T219[2'h3:1'h0];
  assign T219 = T12[3'h7:1'h0];
  assign T220 = T547 & 8'hf;
  assign T547 = {4'h0, T221};
  assign T221 = T219 >> 3'h4;
  assign T222 = T548 & 8'h33;
  assign T548 = {2'h0, T223};
  assign T223 = T215 >> 2'h2;
  assign T224 = T549 & 8'h55;
  assign T549 = {1'h0, T225};
  assign T225 = T211 >> 1'h1;
  assign T226 = T249 | T227;
  assign T227 = T228 & 16'haaaa;
  assign T228 = T229 << 1'h1;
  assign T229 = T230[4'he:1'h0];
  assign T230 = T247 | T231;
  assign T231 = T232 & 16'hcccc;
  assign T232 = T233 << 2'h2;
  assign T233 = T234[4'hd:1'h0];
  assign T234 = T245 | T235;
  assign T235 = T236 & 16'hf0f0;
  assign T236 = T237 << 3'h4;
  assign T237 = T238[4'hb:1'h0];
  assign T238 = T243 | T239;
  assign T239 = T240 & 16'hff00;
  assign T240 = T241 << 4'h8;
  assign T241 = T242[3'h7:1'h0];
  assign T242 = T13[4'hf:1'h0];
  assign T243 = T550 & 16'hff;
  assign T550 = {8'h0, T244};
  assign T244 = T242 >> 4'h8;
  assign T245 = T551 & 16'hf0f;
  assign T551 = {4'h0, T246};
  assign T246 = T238 >> 3'h4;
  assign T247 = T552 & 16'h3333;
  assign T552 = {2'h0, T248};
  assign T248 = T234 >> 2'h2;
  assign T249 = T553 & 16'h5555;
  assign T553 = {1'h0, T250};
  assign T250 = T230 >> 1'h1;
  assign T251 = 27'h0 - T554;
  assign T554 = {26'h0, T252};
  assign T252 = sExpX3[4'ha:4'ha];
  assign sigX3 = T253[5'h1b:1'h0];
  assign T253 = {T380, T254};
  assign T254 = doIncrSig ? T376 : T255;
  assign T255 = T256 != 16'h0;
  assign T256 = T299 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T257, 1'h1};
  assign T257 = {T280, T258};
  assign T258 = {T270, T259};
  assign T259 = {T266, T260};
  assign T260 = T261[2'h2:2'h2];
  assign T261 = T262[3'h6:3'h4];
  assign T262 = T263[4'he:4'h8];
  assign T263 = T264[4'hf:1'h1];
  assign T264 = $signed(17'h10000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T265;
  assign T265 = estNormDist[2'h3:1'h0];
  assign T266 = {T269, T267};
  assign T267 = T268[1'h1:1'h1];
  assign T268 = T261[1'h1:1'h0];
  assign T269 = T268[1'h0:1'h0];
  assign T270 = {T276, T271};
  assign T271 = {T275, T272};
  assign T272 = T273[1'h1:1'h1];
  assign T273 = T274[2'h3:2'h2];
  assign T274 = T262[2'h3:1'h0];
  assign T275 = T273[1'h0:1'h0];
  assign T276 = {T279, T277};
  assign T277 = T278[1'h1:1'h1];
  assign T278 = T274[1'h1:1'h0];
  assign T279 = T278[1'h0:1'h0];
  assign T280 = T297 | T281;
  assign T281 = T282 & 8'haa;
  assign T282 = T283 << 1'h1;
  assign T283 = T284[3'h6:1'h0];
  assign T284 = T295 | T285;
  assign T285 = T286 & 8'hcc;
  assign T286 = T287 << 2'h2;
  assign T287 = T288[3'h5:1'h0];
  assign T288 = T293 | T289;
  assign T289 = T290 & 8'hf0;
  assign T290 = T291 << 3'h4;
  assign T291 = T292[2'h3:1'h0];
  assign T292 = T263[3'h7:1'h0];
  assign T293 = T555 & 8'hf;
  assign T555 = {4'h0, T294};
  assign T294 = T292 >> 3'h4;
  assign T295 = T556 & 8'h33;
  assign T556 = {2'h0, T296};
  assign T296 = T288 >> 2'h2;
  assign T297 = T557 & 8'h55;
  assign T557 = {1'h0, T298};
  assign T298 = T284 >> 1'h1;
  assign T299 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T362 : T558;
  assign T558 = {1'h0, T300};
  assign T300 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T326 ? T320 : T301;
  assign T301 = T319 ? T560 : T302;
  assign T302 = {T304, T303};
  assign T303 = 32'h0 - T559;
  assign T559 = {31'h0, doSubMags};
  assign T304 = sigSum[4'ha:1'h1];
  assign T560 = {8'h0, T305};
  assign T305 = {T318, T306};
  assign T306 = doSubMags ? T312 : T307;
  assign T307 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T310, T308};
  assign T308 = T309 != 18'h0;
  assign T309 = sigSum[5'h11:1'h0];
  assign T310 = T311 != 16'h0;
  assign T311 = sigSum[6'h21:5'h12];
  assign T312 = ~ T313;
  assign T313 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T316, T314};
  assign T314 = T315 != 18'h0;
  assign T315 = notSigSum[5'h11:1'h0];
  assign notSigSum = ~ sigSum;
  assign T316 = T317 != 16'h0;
  assign T317 = notSigSum[6'h21:5'h12];
  assign T318 = sigSum[6'h32:5'h12];
  assign T319 = estNormNeg_dist[3'h4:3'h4];
  assign T320 = T325 ? T322 : T321;
  assign T321 = sigSum[6'h2a:1'h1];
  assign T322 = {T324, T323};
  assign T323 = 16'h0 - T561;
  assign T561 = {15'h0, doSubMags};
  assign T324 = sigSum[5'h1a:1'h1];
  assign T325 = estNormNeg_dist[3'h4:3'h4];
  assign T326 = estNormNeg_dist[3'h5:3'h5];
  assign CDom_firstNormAbsSigSum = T327;
  assign T327 = T335 | T328;
  assign T328 = T562 & T329;
  assign T329 = {T331, T330};
  assign T330 = firstReduceNotSigSum[1'h0:1'h0];
  assign T331 = notSigSum[6'h3a:5'h12];
  assign T562 = T332 ? 42'h3ffffffffff : 42'h0;
  assign T332 = T333;
  assign T333 = doSubMags & T334;
  assign T334 = CDom_estNormDist[3'h4:3'h4];
  assign T335 = T344 | T336;
  assign T336 = T563 & T337;
  assign T337 = {T339, T338};
  assign T338 = firstReduceNotSigSum != 2'h0;
  assign T339 = notSigSum[7'h4a:6'h22];
  assign T563 = T340 ? 42'h3ffffffffff : 42'h0;
  assign T340 = T341;
  assign T341 = doSubMags & T342;
  assign T342 = ~ T343;
  assign T343 = CDom_estNormDist[3'h4:3'h4];
  assign T344 = T353 | T345;
  assign T345 = T564 & T346;
  assign T346 = {T348, T347};
  assign T347 = firstReduceSigSum[1'h0:1'h0];
  assign T348 = sigSum[6'h3a:5'h12];
  assign T564 = T349 ? 42'h3ffffffffff : 42'h0;
  assign T349 = T350;
  assign T350 = T352 & T351;
  assign T351 = CDom_estNormDist[3'h4:3'h4];
  assign T352 = ~ doSubMags;
  assign T353 = T565 & T354;
  assign T354 = {T356, T355};
  assign T355 = firstReduceSigSum != 2'h0;
  assign T356 = sigSum[7'h4a:6'h22];
  assign T565 = T357 ? 42'h3ffffffffff : 42'h0;
  assign T357 = T358;
  assign T358 = T361 & T359;
  assign T359 = ~ T360;
  assign T360 = CDom_estNormDist[3'h4:3'h4];
  assign T361 = ~ doSubMags;
  assign T362 = isCDominant ? T568 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T375 ? T370 : T363;
  assign T363 = T369 ? T566 : T364;
  assign T364 = T365 << 6'h20;
  assign T365 = notSigSum[4'hb:1'h1];
  assign T566 = {10'h0, T366};
  assign T366 = {T368, T367};
  assign T367 = firstReduceNotSigSum[1'h0:1'h0];
  assign T368 = notSigSum[6'h31:5'h12];
  assign T369 = estNormNeg_dist[3'h4:3'h4];
  assign T370 = T374 ? T372 : T567;
  assign T567 = {1'h0, T371};
  assign T371 = notSigSum[6'h2a:1'h1];
  assign T372 = T373 << 5'h10;
  assign T373 = notSigSum[5'h1b:1'h1];
  assign T374 = estNormNeg_dist[3'h4:3'h4];
  assign T375 = estNormNeg_dist[3'h5:3'h5];
  assign T568 = {1'h0, CDom_firstNormAbsSigSum};
  assign T376 = T377 == 16'h0;
  assign T377 = T378 & absSigSumExtraMask;
  assign T378 = ~ T379;
  assign T379 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign T380 = T381 >> normTo2ShiftDist;
  assign T381 = cFirstNormAbsSigSum[6'h2a:1'h1];
  assign roundPosBit = T382 != 28'h0;
  assign T382 = sigX3 & T569;
  assign T569 = {1'h0, roundPosMask};
  assign roundPosMask = T570 & roundMask;
  assign T570 = {1'h0, T383};
  assign T383 = ~ T384;
  assign T384 = roundMask >> 1'h1;
  assign T385 = ~ allRound;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T386 == 28'h0;
  assign T386 = T388 & T571;
  assign T571 = {2'h0, T387};
  assign T387 = roundMask >> 1'h1;
  assign T388 = ~ sigX3;
  assign doIncrSig = T389 & doSubMags;
  assign T389 = T391 & T390;
  assign T390 = ~ notCDom_signSigSum;
  assign T391 = ~ isCDominant;
  assign commonCase = T393 & T392;
  assign T392 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T393 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T394 == 2'h3;
  assign T394 = expC[4'h8:3'h7];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T395 == 2'h3;
  assign T395 = expB[4'h8:3'h7];
  assign isSpecialA = T396 == 2'h3;
  assign T396 = expA[4'h8:3'h7];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T397;
  assign T397 = T401 | T398;
  assign T398 = sExpX3_13 <= T572;
  assign T572 = {2'h0, T399};
  assign T399 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign sigX3Shift1 = T400 == 2'h0;
  assign T400 = sigX3[5'h1b:5'h1a];
  assign T401 = sExpX3[4'ha:4'ha];
  assign overflow = commonCase & overflowY;
  assign overflowY = T402 == 3'h3;
  assign T402 = sExpY[4'h9:3'h7];
  assign sExpY = T449 | T403;
  assign T403 = T405 ? T404 : 11'h0;
  assign T404 = sExpX3 - 11'h1;
  assign T405 = T406 == 2'h0;
  assign T406 = sigY3[5'h19:5'h18];
  assign sigY3 = T420 | T407;
  assign T407 = roundEven ? T408 : 26'h0;
  assign T408 = roundUp_sigY3 & T409;
  assign T409 = ~ T410;
  assign T410 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T411[5'h19:1'h0];
  assign T411 = T412 + 26'h1;
  assign T412 = T413 >> 2'h2;
  assign T413 = sigX3 | T573;
  assign T573 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T417 : T414;
  assign T414 = T416 & T415;
  assign T415 = ~ anyRoundExtra;
  assign T416 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T417 = T418 & allRoundExtra;
  assign T418 = roundingMode_nearest_even & T419;
  assign T419 = ~ roundPosBit;
  assign T420 = T442 | T421;
  assign T421 = roundUp ? roundUp_sigY3 : 26'h0;
  assign roundUp = T429 | T422;
  assign T422 = T423 & 1'h1;
  assign T423 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T427 & T424;
  assign T424 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T425 : notCDom_signSigSum;
  assign T425 = doSubMags & T426;
  assign T426 = ~ isZeroC;
  assign T427 = ~ isZeroY;
  assign isZeroY = T428 == 3'h0;
  assign T428 = sigX3[5'h1b:5'h19];
  assign T429 = T432 | T430;
  assign T430 = T431 & roundPosBit;
  assign T431 = doIncrSig & roundingMode_nearest_even;
  assign T432 = T434 | T433;
  assign T433 = doIncrSig & allRound;
  assign T434 = T438 | T435;
  assign T435 = T436 & anyRound;
  assign T436 = T437 & roundDirectUp;
  assign T437 = ~ doIncrSig;
  assign T438 = T439 & anyRoundExtra;
  assign T439 = T440 & roundPosBit;
  assign T440 = T441 & roundingMode_nearest_even;
  assign T441 = ~ doIncrSig;
  assign T442 = T446 ? T443 : 26'h0;
  assign T443 = T444 >> 2'h2;
  assign T444 = sigX3 & T574;
  assign T574 = {1'h0, T445};
  assign T445 = ~ roundMask;
  assign T446 = T448 & T447;
  assign T447 = ~ roundEven;
  assign T448 = ~ roundUp;
  assign T449 = T452 | T450;
  assign T450 = T451 ? sExpX3 : 11'h0;
  assign T451 = sigY3[5'h18:5'h18];
  assign T452 = T454 ? T453 : 11'h0;
  assign T453 = sExpX3 + 11'h1;
  assign T454 = sigY3[5'h19:5'h19];
  assign T455 = {invalid, 1'h0};
  assign invalid = T474 | notSigNaN_invalid;
  assign notSigNaN_invalid = T471 | T456;
  assign T456 = T457 & doSubMags;
  assign T457 = T460 & isInfC;
  assign isInfC = isSpecialC & T458;
  assign T458 = T459 ^ 1'h1;
  assign T459 = expC[3'h6:3'h6];
  assign T460 = T466 & T461;
  assign T461 = isInfA | isInfB;
  assign isInfB = isSpecialB & T462;
  assign T462 = T463 ^ 1'h1;
  assign T463 = expB[3'h6:3'h6];
  assign isInfA = isSpecialA & T464;
  assign T464 = T465 ^ 1'h1;
  assign T465 = expA[3'h6:3'h6];
  assign T466 = T469 & T467;
  assign T467 = ~ isNaNB;
  assign isNaNB = isSpecialB & T468;
  assign T468 = expB[3'h6:3'h6];
  assign T469 = ~ isNaNA;
  assign isNaNA = isSpecialA & T470;
  assign T470 = expA[3'h6:3'h6];
  assign T471 = T473 | T472;
  assign T472 = isZeroA & isInfB;
  assign T473 = isInfA & isZeroB;
  assign T474 = T478 | isSigNaNC;
  assign isSigNaNC = isNaNC & T475;
  assign T475 = T476 ^ 1'h1;
  assign T476 = fractC[5'h16:5'h16];
  assign isNaNC = isSpecialC & T477;
  assign T477 = expC[3'h6:3'h6];
  assign T478 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T479;
  assign T479 = T480 ^ 1'h1;
  assign T480 = fractB[5'h16:5'h16];
  assign isSigNaNA = isNaNA & T481;
  assign T481 = T482 ^ 1'h1;
  assign T482 = fractA[5'h16:5'h16];
  assign io_out = T483;
  assign T483 = {signOut, T484};
  assign T484 = {expOut, fractOut};
  assign fractOut = fractY | T485;
  assign T485 = 23'h0 - T575;
  assign T575 = {22'h0, T486};
  assign T486 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T487;
  assign T487 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T490 | T488;
  assign T488 = roundingMode_max & T489;
  assign T489 = ~ signY;
  assign T490 = roundingMode_nearest_even | T491;
  assign T491 = roundingMode_min & signY;
  assign isNaNOut = T492 | notSigNaN_invalid;
  assign T492 = T493 | isNaNC;
  assign T493 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T495 : T494;
  assign T494 = sigY3[5'h17:1'h1];
  assign T495 = sigY3[5'h16:1'h0];
  assign expOut = T497 | T496;
  assign T496 = isNaNOut ? 9'h1c0 : 9'h0;
  assign T497 = T502 | T498;
  assign T498 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign notNaN_isInfOut = T500 | T499;
  assign T499 = overflow & overflowY_roundMagUp;
  assign T500 = T501 | isInfC;
  assign T501 = isInfA | isInfB;
  assign T502 = T504 | T503;
  assign T503 = isSatOut ? 9'h17f : 9'h0;
  assign T504 = T507 & T505;
  assign T505 = ~ T506;
  assign T506 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T507 = T510 & T508;
  assign T508 = ~ T509;
  assign T509 = isSatOut ? 9'h80 : 9'h0;
  assign T510 = expY & T511;
  assign T511 = ~ T512;
  assign T512 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign notSpecial_isZeroOut = T516 | totalUnderflowY;
  assign totalUnderflowY = T515 | T513;
  assign T513 = T514 < 9'h6b;
  assign T514 = sExpY[4'h8:1'h0];
  assign T515 = sExpY[4'h9:4'h9];
  assign T516 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'h8:1'h0];
  assign signOut = T518 | T517;
  assign T517 = commonCase & signY;
  assign T518 = T522 | T519;
  assign T519 = T520 & opSignC;
  assign T520 = T521 & isSpecialC;
  assign T521 = mulSpecial ^ 1'h1;
  assign T522 = T526 | T523;
  assign T523 = T524 & signProd;
  assign T524 = mulSpecial & T525;
  assign T525 = isSpecialC ^ 1'h1;
  assign T526 = T527 | isNaNOut;
  assign T527 = T528 & opSignC;
  assign T528 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_0(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T7;
  reg [2:0] in_rm;
  wire[2:0] T8;
  wire[32:0] T9;
  reg [64:0] in_in3;
  wire[64:0] T10;
  wire[64:0] T11;
  wire[64:0] T12;
  wire[32:0] zero;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[32:0] T19;
  reg [64:0] in_in2;
  wire[64:0] T20;
  wire[64:0] T21;
  wire T22;
  wire[32:0] T23;
  reg [64:0] in_in1;
  wire[64:0] T24;
  wire[1:0] T25;
  reg [4:0] in_cmd;
  wire[4:0] T26;
  wire[4:0] T27;
  wire[4:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg [4:0] R0;
  wire[4:0] T1;
  wire[4:0] res_exc;
  reg  valid;
  reg [64:0] R2;
  wire[64:0] T3;
  wire[64:0] res_data;
  wire[64:0] T5;
  reg  R4;
  wire T6;
  wire[32:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R0 = {1{$random}};
    valid = {1{$random}};
    R2 = {3{$random}};
    R4 = {1{$random}};
  end
`endif

  assign T7 = in_rm[1'h1:1'h0];
  assign T8 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T9 = in_in3[6'h20:1'h0];
  assign T10 = T16 ? T12 : T11;
  assign T11 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T12 = {32'h0, zero};
  assign zero = T13 << 6'h20;
  assign T13 = T15 ^ T14;
  assign T14 = io_in_bits_in2[6'h20:6'h20];
  assign T15 = io_in_bits_in1[6'h20:6'h20];
  assign T16 = io_in_valid & T17;
  assign T17 = T18 ^ 1'h1;
  assign T18 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T19 = in_in2[6'h20:1'h0];
  assign T20 = T22 ? 65'h80000000 : T21;
  assign T21 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T22 = io_in_valid & io_in_bits_swap23;
  assign T23 = in_in1[6'h20:1'h0];
  assign T24 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T25 = in_cmd[1'h1:1'h0];
  assign T26 = io_in_valid ? T28 : T27;
  assign T27 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T28 = {3'h0, T29};
  assign T29 = {T31, T30};
  assign T30 = io_in_bits_cmd[1'h0:1'h0];
  assign T31 = T33 & T32;
  assign T32 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T33 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R0;
  assign T1 = valid ? res_exc : R0;
  assign res_exc = fma_io_exceptionFlags;
  assign io_out_bits_data = R2;
  assign T3 = valid ? res_data : R2;
  assign res_data = T5;
  assign T5 = {32'h0, fma_io_out};
  assign io_out_valid = R4;
  assign T6 = reset ? 1'h0 : valid;
  mulAddSubRecodedFloatN_0 fma(
       .io_op( T25 ),
       .io_a( T23 ),
       .io_b( T19 ),
       .io_c( T9 ),
       .io_roundingMode( T7 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T16) begin
      in_in3 <= T12;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T22) begin
      in_in2 <= 65'h80000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T28;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(valid) begin
      R0 <= res_exc;
    end
    valid <= io_in_valid;
    if(valid) begin
      R2 <= res_data;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else begin
      R4 <= valid;
    end
  end
endmodule

module mulAddSubRecodedFloatN_1(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[56:0] T4;
  wire[56:0] T744;
  wire[54:0] T5;
  wire[55:0] roundMask;
  wire[55:0] T6;
  wire[53:0] T7;
  wire[53:0] T745;
  wire T8;
  wire[53:0] T9;
  wire[21:0] T10;
  wire[5:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[5:0] T15;
  wire[21:0] T16;
  wire[53:0] T17;
  wire[8192:0] T18;
  wire[12:0] T19;
  wire[12:0] sExpX3_13;
  wire[13:0] sExpX3;
  wire[13:0] T746;
  wire[7:0] estNormDist;
  wire[7:0] T20;
  wire[7:0] estNormNeg_dist;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[7:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[7:0] T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[7:0] T58;
  wire[7:0] T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire[7:0] T75;
  wire[7:0] T76;
  wire[7:0] T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire[7:0] T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T119;
  wire[7:0] T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire T127;
  wire[108:0] T128;
  wire[108:0] T129;
  wire[107:0] T130;
  wire[107:0] T131;
  wire[161:0] sigSum;
  wire[161:0] alignedNegSigC;
  wire[162:0] T132;
  wire T133;
  wire doSubMags;
  wire opSignC;
  wire T134;
  wire T135;
  wire signProd;
  wire T136;
  wire T137;
  wire signB;
  wire signA;
  wire T138;
  wire[52:0] T139;
  wire[52:0] CExtraMask;
  wire[20:0] T140;
  wire[4:0] T141;
  wire T142;
  wire[4:0] T143;
  wire[20:0] T144;
  wire[52:0] T145;
  wire[256:0] T146;
  wire[7:0] CAlignDist;
  wire[13:0] T147;
  wire[13:0] T148;
  wire[13:0] sNatCAlignDist;
  wire[13:0] T747;
  wire[11:0] expC;
  wire[13:0] sExpAlignedProd;
  wire[13:0] T149;
  wire[13:0] T748;
  wire[11:0] expA;
  wire[13:0] T150;
  wire[10:0] T151;
  wire[11:0] expB;
  wire[2:0] T152;
  wire[2:0] T749;
  wire T153;
  wire T154;
  wire T155;
  wire[12:0] T156;
  wire CAlignDist_floor;
  wire T157;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T158;
  wire isZeroA;
  wire[2:0] T159;
  wire[3:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[1:0] T163;
  wire[3:0] T164;
  wire T165;
  wire[1:0] T166;
  wire T167;
  wire[1:0] T168;
  wire T169;
  wire[15:0] T170;
  wire[15:0] T171;
  wire[15:0] T172;
  wire[14:0] T173;
  wire[15:0] T174;
  wire[15:0] T175;
  wire[15:0] T176;
  wire[13:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[15:0] T180;
  wire[11:0] T181;
  wire[15:0] T182;
  wire[15:0] T183;
  wire[15:0] T184;
  wire[7:0] T185;
  wire[15:0] T186;
  wire[15:0] T187;
  wire[15:0] T750;
  wire[7:0] T188;
  wire[15:0] T189;
  wire[15:0] T751;
  wire[11:0] T190;
  wire[15:0] T191;
  wire[15:0] T752;
  wire[13:0] T192;
  wire[15:0] T193;
  wire[15:0] T753;
  wire[14:0] T194;
  wire[31:0] T195;
  wire[31:0] T196;
  wire[31:0] T197;
  wire[30:0] T198;
  wire[31:0] T199;
  wire[31:0] T200;
  wire[31:0] T201;
  wire[29:0] T202;
  wire[31:0] T203;
  wire[31:0] T204;
  wire[31:0] T205;
  wire[27:0] T206;
  wire[31:0] T207;
  wire[31:0] T208;
  wire[31:0] T209;
  wire[23:0] T210;
  wire[31:0] T211;
  wire[31:0] T212;
  wire[31:0] T213;
  wire[15:0] T214;
  wire[31:0] T215;
  wire[31:0] T216;
  wire[31:0] T754;
  wire[15:0] T217;
  wire[31:0] T218;
  wire[31:0] T755;
  wire[23:0] T219;
  wire[31:0] T220;
  wire[31:0] T756;
  wire[27:0] T221;
  wire[31:0] T222;
  wire[31:0] T757;
  wire[29:0] T223;
  wire[31:0] T224;
  wire[31:0] T758;
  wire[30:0] T225;
  wire[52:0] sigC;
  wire[51:0] fractC;
  wire T226;
  wire isZeroC;
  wire[2:0] T227;
  wire[161:0] T228;
  wire[161:0] T229;
  wire[161:0] T230;
  wire[160:0] T231;
  wire[107:0] T232;
  wire[107:0] T759;
  wire[52:0] negSigC;
  wire[52:0] T233;
  wire[161:0] T760;
  wire[106:0] T234;
  wire[105:0] T235;
  wire[52:0] sigB;
  wire[51:0] fractB;
  wire T236;
  wire[52:0] sigA;
  wire[51:0] fractA;
  wire T237;
  wire[108:0] T761;
  wire[107:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire notCDom_signSigSum;
  wire[7:0] CDom_estNormDist;
  wire[7:0] T762;
  wire[5:0] T345;
  wire[7:0] T346;
  wire T347;
  wire CAlignDist_0;
  wire T348;
  wire[12:0] T349;
  wire isCDominant;
  wire T350;
  wire T351;
  wire[12:0] T352;
  wire T353;
  wire[13:0] sExpSum;
  wire[13:0] T763;
  wire T354;
  wire[3:0] T355;
  wire[1:0] T356;
  wire T357;
  wire[1:0] T358;
  wire[3:0] T359;
  wire T360;
  wire[1:0] T361;
  wire T362;
  wire[1:0] T363;
  wire T364;
  wire[15:0] T365;
  wire[15:0] T366;
  wire[15:0] T367;
  wire[14:0] T368;
  wire[15:0] T369;
  wire[15:0] T370;
  wire[15:0] T371;
  wire[13:0] T372;
  wire[15:0] T373;
  wire[15:0] T374;
  wire[15:0] T375;
  wire[11:0] T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[7:0] T380;
  wire[15:0] T381;
  wire[15:0] T382;
  wire[15:0] T764;
  wire[7:0] T383;
  wire[15:0] T384;
  wire[15:0] T765;
  wire[11:0] T385;
  wire[15:0] T386;
  wire[15:0] T766;
  wire[13:0] T387;
  wire[15:0] T388;
  wire[15:0] T767;
  wire[14:0] T389;
  wire[31:0] T390;
  wire[31:0] T391;
  wire[31:0] T392;
  wire[30:0] T393;
  wire[31:0] T394;
  wire[31:0] T395;
  wire[31:0] T396;
  wire[29:0] T397;
  wire[31:0] T398;
  wire[31:0] T399;
  wire[31:0] T400;
  wire[27:0] T401;
  wire[31:0] T402;
  wire[31:0] T403;
  wire[31:0] T404;
  wire[23:0] T405;
  wire[31:0] T406;
  wire[31:0] T407;
  wire[31:0] T408;
  wire[15:0] T409;
  wire[31:0] T410;
  wire[31:0] T411;
  wire[31:0] T768;
  wire[15:0] T412;
  wire[31:0] T413;
  wire[31:0] T769;
  wire[23:0] T414;
  wire[31:0] T415;
  wire[31:0] T770;
  wire[27:0] T416;
  wire[31:0] T417;
  wire[31:0] T771;
  wire[29:0] T418;
  wire[31:0] T419;
  wire[31:0] T772;
  wire[30:0] T420;
  wire[55:0] T421;
  wire[55:0] T773;
  wire T422;
  wire[56:0] sigX3;
  wire[87:0] T423;
  wire T424;
  wire T425;
  wire[31:0] T426;
  wire[31:0] absSigSumExtraMask;
  wire[30:0] T427;
  wire[14:0] T428;
  wire[6:0] T429;
  wire[2:0] T430;
  wire T431;
  wire[2:0] T432;
  wire[6:0] T433;
  wire[14:0] T434;
  wire[30:0] T435;
  wire[32:0] T436;
  wire[4:0] normTo2ShiftDist;
  wire[4:0] estNormDist_5;
  wire[4:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[1:0] T440;
  wire T441;
  wire[3:0] T442;
  wire[1:0] T443;
  wire T444;
  wire[1:0] T445;
  wire[3:0] T446;
  wire T447;
  wire[1:0] T448;
  wire T449;
  wire[1:0] T450;
  wire T451;
  wire[7:0] T452;
  wire[7:0] T453;
  wire[7:0] T454;
  wire[6:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[5:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[3:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T774;
  wire[3:0] T466;
  wire[7:0] T467;
  wire[7:0] T775;
  wire[5:0] T468;
  wire[7:0] T469;
  wire[7:0] T776;
  wire[6:0] T470;
  wire[15:0] T471;
  wire[15:0] T472;
  wire[15:0] T473;
  wire[14:0] T474;
  wire[15:0] T475;
  wire[15:0] T476;
  wire[15:0] T477;
  wire[13:0] T478;
  wire[15:0] T479;
  wire[15:0] T480;
  wire[15:0] T481;
  wire[11:0] T482;
  wire[15:0] T483;
  wire[15:0] T484;
  wire[15:0] T485;
  wire[7:0] T486;
  wire[15:0] T487;
  wire[15:0] T488;
  wire[15:0] T777;
  wire[7:0] T489;
  wire[15:0] T490;
  wire[15:0] T778;
  wire[11:0] T491;
  wire[15:0] T492;
  wire[15:0] T779;
  wire[13:0] T493;
  wire[15:0] T494;
  wire[15:0] T780;
  wire[14:0] T495;
  wire[31:0] T496;
  wire[87:0] cFirstNormAbsSigSum;
  wire[87:0] T781;
  wire[86:0] T497;
  wire[86:0] notCDom_pos_firstNormAbsSigSum;
  wire[86:0] T498;
  wire[86:0] T499;
  wire[53:0] T500;
  wire[53:0] T782;
  wire[32:0] T501;
  wire[86:0] T502;
  wire[86:0] T503;
  wire[85:0] T504;
  wire[85:0] T783;
  wire T505;
  wire[86:0] T784;
  wire[65:0] T506;
  wire T507;
  wire T508;
  wire[1:0] firstReduceSigSum;
  wire T509;
  wire[43:0] T510;
  wire T511;
  wire[31:0] T512;
  wire T513;
  wire T514;
  wire[1:0] firstReduceNotSigSum;
  wire T515;
  wire[43:0] T516;
  wire[161:0] notSigSum;
  wire T517;
  wire[31:0] T518;
  wire[64:0] T519;
  wire T520;
  wire T521;
  wire[86:0] T522;
  wire[86:0] T523;
  wire T524;
  wire T525;
  wire[10:0] T526;
  wire T527;
  wire[10:0] T528;
  wire[85:0] T529;
  wire[86:0] T530;
  wire[21:0] T531;
  wire[21:0] T785;
  wire[64:0] T532;
  wire T533;
  wire T534;
  wire[86:0] CDom_firstNormAbsSigSum;
  wire[86:0] T535;
  wire[86:0] T536;
  wire[86:0] T537;
  wire T538;
  wire[85:0] T539;
  wire[86:0] T786;
  wire T540;
  wire T541;
  wire T542;
  wire[86:0] T543;
  wire[86:0] T544;
  wire[86:0] T545;
  wire T546;
  wire[85:0] T547;
  wire[86:0] T787;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire[86:0] T552;
  wire[86:0] T553;
  wire[86:0] T554;
  wire T555;
  wire[85:0] T556;
  wire[86:0] T788;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire[86:0] T561;
  wire[86:0] T562;
  wire T563;
  wire[85:0] T564;
  wire[86:0] T789;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire[87:0] T570;
  wire[87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[87:0] T571;
  wire[87:0] T572;
  wire[33:0] T573;
  wire[87:0] T574;
  wire[87:0] T575;
  wire[1:0] T576;
  wire[87:0] T790;
  wire[64:0] T577;
  wire T578;
  wire[63:0] T579;
  wire T580;
  wire T581;
  wire[87:0] T582;
  wire[87:0] T583;
  wire T584;
  wire[10:0] T585;
  wire[86:0] T586;
  wire[87:0] T587;
  wire[65:0] T588;
  wire T589;
  wire T590;
  wire[87:0] T791;
  wire T591;
  wire[31:0] T592;
  wire[31:0] T593;
  wire[31:0] T594;
  wire[86:0] T595;
  wire[86:0] T596;
  wire roundPosBit;
  wire[56:0] T597;
  wire[56:0] T792;
  wire[55:0] roundPosMask;
  wire[55:0] T793;
  wire[54:0] T598;
  wire[54:0] T599;
  wire T600;
  wire allRound;
  wire allRoundExtra;
  wire[56:0] T601;
  wire[56:0] T794;
  wire[54:0] T602;
  wire[56:0] T603;
  wire doIncrSig;
  wire T604;
  wire T605;
  wire T606;
  wire commonCase;
  wire T607;
  wire notSpecial_addZeros;
  wire T608;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T609;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T610;
  wire isSpecialA;
  wire[1:0] T611;
  wire underflow;
  wire underflowY;
  wire T612;
  wire T613;
  wire[12:0] T795;
  wire[10:0] T614;
  wire sigX3Shift1;
  wire[1:0] T615;
  wire T616;
  wire overflow;
  wire overflowY;
  wire[2:0] T617;
  wire[13:0] sExpY;
  wire[13:0] T618;
  wire[13:0] T619;
  wire T620;
  wire[1:0] T621;
  wire[54:0] sigY3;
  wire[54:0] T622;
  wire[54:0] T623;
  wire[54:0] T624;
  wire[54:0] T625;
  wire[54:0] roundUp_sigY3;
  wire[54:0] T626;
  wire[54:0] T627;
  wire[56:0] T628;
  wire[56:0] T796;
  wire roundEven;
  wire T629;
  wire T630;
  wire T631;
  wire roundingMode_nearest_even;
  wire T632;
  wire T633;
  wire T634;
  wire[54:0] T635;
  wire[54:0] T636;
  wire roundUp;
  wire T637;
  wire T638;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T639;
  wire doNegSignSum;
  wire T640;
  wire T641;
  wire T642;
  wire isZeroY;
  wire[2:0] T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire[54:0] T657;
  wire[54:0] T658;
  wire[56:0] T659;
  wire[56:0] T797;
  wire[55:0] T660;
  wire T661;
  wire T662;
  wire T663;
  wire[13:0] T664;
  wire[13:0] T665;
  wire T666;
  wire[13:0] T667;
  wire[13:0] T668;
  wire T669;
  wire[1:0] T670;
  wire invalid;
  wire notSigNaN_invalid;
  wire T671;
  wire T672;
  wire isInfC;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire isInfB;
  wire T677;
  wire T678;
  wire isInfA;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire isNaNB;
  wire T683;
  wire T684;
  wire isNaNA;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire isSigNaNC;
  wire T690;
  wire T691;
  wire isNaNC;
  wire T692;
  wire T693;
  wire isSigNaNB;
  wire T694;
  wire T695;
  wire isSigNaNA;
  wire T696;
  wire T697;
  wire[64:0] T698;
  wire[63:0] T699;
  wire[51:0] fractOut;
  wire[51:0] T700;
  wire[51:0] T798;
  wire T701;
  wire isSatOut;
  wire T702;
  wire overflowY_roundMagUp;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire isNaNOut;
  wire T707;
  wire T708;
  wire[51:0] fractY;
  wire[51:0] T709;
  wire[51:0] T710;
  wire[11:0] expOut;
  wire[11:0] T711;
  wire[11:0] T712;
  wire[11:0] T713;
  wire notNaN_isInfOut;
  wire T714;
  wire T715;
  wire T716;
  wire[11:0] T717;
  wire[11:0] T718;
  wire[11:0] T719;
  wire[11:0] T720;
  wire[11:0] T721;
  wire[11:0] T722;
  wire[11:0] T723;
  wire[11:0] T724;
  wire[11:0] T725;
  wire[11:0] T726;
  wire[11:0] T727;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T728;
  wire[11:0] T729;
  wire T730;
  wire T731;
  wire[11:0] expY;
  wire signOut;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;


  assign io_exceptionFlags = T0;
  assign T0 = {T670, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T600 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 57'h0;
  assign T4 = sigX3 & T744;
  assign T744 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T421 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T745;
  assign T745 = {53'h0, T8};
  assign T8 = sigX3[6'h37:6'h37];
  assign T9 = {T390, T10};
  assign T10 = {T365, T11};
  assign T11 = {T355, T12};
  assign T12 = {T354, T13};
  assign T13 = T14[1'h1:1'h1];
  assign T14 = T15[3'h5:3'h4];
  assign T15 = T16[5'h15:5'h10];
  assign T16 = T17[6'h35:6'h20];
  assign T17 = T18[11'h403:10'h3ce];
  assign T18 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T19;
  assign T19 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'hc:1'h0];
  assign sExpX3 = sExpSum - T746;
  assign T746 = {6'h0, estNormDist};
  assign estNormDist = isCDominant ? CDom_estNormDist : T20;
  assign T20 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = T344 ? 8'h35 : T21;
  assign T21 = T343 ? 8'h36 : T22;
  assign T22 = T342 ? 8'h37 : T23;
  assign T23 = T341 ? 8'h38 : T24;
  assign T24 = T340 ? 8'h39 : T25;
  assign T25 = T339 ? 8'h3a : T26;
  assign T26 = T338 ? 8'h3b : T27;
  assign T27 = T337 ? 8'h3c : T28;
  assign T28 = T336 ? 8'h3d : T29;
  assign T29 = T335 ? 8'h3e : T30;
  assign T30 = T334 ? 8'h3f : T31;
  assign T31 = T333 ? 8'h40 : T32;
  assign T32 = T332 ? 8'h41 : T33;
  assign T33 = T331 ? 8'h42 : T34;
  assign T34 = T330 ? 8'h43 : T35;
  assign T35 = T329 ? 8'h44 : T36;
  assign T36 = T328 ? 8'h45 : T37;
  assign T37 = T327 ? 8'h46 : T38;
  assign T38 = T326 ? 8'h47 : T39;
  assign T39 = T325 ? 8'h48 : T40;
  assign T40 = T324 ? 8'h49 : T41;
  assign T41 = T323 ? 8'h4a : T42;
  assign T42 = T322 ? 8'h4b : T43;
  assign T43 = T321 ? 8'h4c : T44;
  assign T44 = T320 ? 8'h4d : T45;
  assign T45 = T319 ? 8'h4e : T46;
  assign T46 = T318 ? 8'h4f : T47;
  assign T47 = T317 ? 8'h50 : T48;
  assign T48 = T316 ? 8'h51 : T49;
  assign T49 = T315 ? 8'h52 : T50;
  assign T50 = T314 ? 8'h53 : T51;
  assign T51 = T313 ? 8'h54 : T52;
  assign T52 = T312 ? 8'h55 : T53;
  assign T53 = T311 ? 8'h56 : T54;
  assign T54 = T310 ? 8'h57 : T55;
  assign T55 = T309 ? 8'h58 : T56;
  assign T56 = T308 ? 8'h59 : T57;
  assign T57 = T307 ? 8'h5a : T58;
  assign T58 = T306 ? 8'h5b : T59;
  assign T59 = T305 ? 8'h5c : T60;
  assign T60 = T304 ? 8'h5d : T61;
  assign T61 = T303 ? 8'h5e : T62;
  assign T62 = T302 ? 8'h5f : T63;
  assign T63 = T301 ? 8'h60 : T64;
  assign T64 = T300 ? 8'h61 : T65;
  assign T65 = T299 ? 8'h62 : T66;
  assign T66 = T298 ? 8'h63 : T67;
  assign T67 = T297 ? 8'h64 : T68;
  assign T68 = T296 ? 8'h65 : T69;
  assign T69 = T295 ? 8'h66 : T70;
  assign T70 = T294 ? 8'h67 : T71;
  assign T71 = T293 ? 8'h68 : T72;
  assign T72 = T292 ? 8'h69 : T73;
  assign T73 = T291 ? 8'h6a : T74;
  assign T74 = T290 ? 8'h6b : T75;
  assign T75 = T289 ? 8'h6c : T76;
  assign T76 = T288 ? 8'h6d : T77;
  assign T77 = T287 ? 8'h6e : T78;
  assign T78 = T286 ? 8'h6f : T79;
  assign T79 = T285 ? 8'h70 : T80;
  assign T80 = T284 ? 8'h71 : T81;
  assign T81 = T283 ? 8'h72 : T82;
  assign T82 = T282 ? 8'h73 : T83;
  assign T83 = T281 ? 8'h74 : T84;
  assign T84 = T280 ? 8'h75 : T85;
  assign T85 = T279 ? 8'h76 : T86;
  assign T86 = T278 ? 8'h77 : T87;
  assign T87 = T277 ? 8'h78 : T88;
  assign T88 = T276 ? 8'h79 : T89;
  assign T89 = T275 ? 8'h7a : T90;
  assign T90 = T274 ? 8'h7b : T91;
  assign T91 = T273 ? 8'h7c : T92;
  assign T92 = T272 ? 8'h7d : T93;
  assign T93 = T271 ? 8'h7e : T94;
  assign T94 = T270 ? 8'h7f : T95;
  assign T95 = T269 ? 8'h80 : T96;
  assign T96 = T268 ? 8'h81 : T97;
  assign T97 = T267 ? 8'h82 : T98;
  assign T98 = T266 ? 8'h83 : T99;
  assign T99 = T265 ? 8'h84 : T100;
  assign T100 = T264 ? 8'h85 : T101;
  assign T101 = T263 ? 8'h86 : T102;
  assign T102 = T262 ? 8'h87 : T103;
  assign T103 = T261 ? 8'h88 : T104;
  assign T104 = T260 ? 8'h89 : T105;
  assign T105 = T259 ? 8'h8a : T106;
  assign T106 = T258 ? 8'h8b : T107;
  assign T107 = T257 ? 8'h8c : T108;
  assign T108 = T256 ? 8'h8d : T109;
  assign T109 = T255 ? 8'h8e : T110;
  assign T110 = T254 ? 8'h8f : T111;
  assign T111 = T253 ? 8'h90 : T112;
  assign T112 = T252 ? 8'h91 : T113;
  assign T113 = T251 ? 8'h92 : T114;
  assign T114 = T250 ? 8'h93 : T115;
  assign T115 = T249 ? 8'h94 : T116;
  assign T116 = T248 ? 8'h95 : T117;
  assign T117 = T247 ? 8'h96 : T118;
  assign T118 = T246 ? 8'h97 : T119;
  assign T119 = T245 ? 8'h98 : T120;
  assign T120 = T244 ? 8'h99 : T121;
  assign T121 = T243 ? 8'h9a : T122;
  assign T122 = T242 ? 8'h9b : T123;
  assign T123 = T241 ? 8'h9c : T124;
  assign T124 = T240 ? 8'h9d : T125;
  assign T125 = T239 ? 8'h9e : T126;
  assign T126 = T127 ? 8'h9f : 8'ha0;
  assign T127 = T128[1'h1:1'h1];
  assign T128 = T761 ^ T129;
  assign T129 = T130 << 1'h1;
  assign T130 = 108'h0 | T131;
  assign T131 = sigSum[7'h6c:1'h1];
  assign sigSum = T760 + alignedNegSigC;
  assign alignedNegSigC = T132[8'ha1:1'h0];
  assign T132 = {T228, T133};
  assign T133 = T138 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T135 ^ T134;
  assign T134 = io_op[1'h0:1'h0];
  assign T135 = io_c[7'h40:7'h40];
  assign signProd = T137 ^ T136;
  assign T136 = io_op[1'h1:1'h1];
  assign T137 = signA ^ signB;
  assign signB = io_b[7'h40:7'h40];
  assign signA = io_a[7'h40:7'h40];
  assign T138 = T139 != 53'h0;
  assign T139 = sigC & CExtraMask;
  assign CExtraMask = {T195, T140};
  assign T140 = {T170, T141};
  assign T141 = {T160, T142};
  assign T142 = T143[3'h4:3'h4];
  assign T143 = T144[5'h14:5'h10];
  assign T144 = T145[6'h34:6'h20];
  assign T145 = T146[8'h93:7'h5f];
  assign T146 = $signed(257'h10000000000000000000000000000000000000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = T147[3'h7:1'h0];
  assign T147 = CAlignDist_floor ? 14'h0 : T148;
  assign T148 = T155 ? sNatCAlignDist : 14'ha1;
  assign sNatCAlignDist = sExpAlignedProd - T747;
  assign T747 = {2'h0, expC};
  assign expC = io_c[6'h3f:6'h34];
  assign sExpAlignedProd = T149 + 14'h38;
  assign T149 = T150 + T748;
  assign T748 = {2'h0, expA};
  assign expA = io_a[6'h3f:6'h34];
  assign T150 = {T152, T151};
  assign T151 = expB[4'ha:1'h0];
  assign expB = io_b[6'h3f:6'h34];
  assign T152 = 3'h0 - T749;
  assign T749 = {2'h0, T153};
  assign T153 = T154 ^ 1'h1;
  assign T154 = expB[4'hb:4'hb];
  assign T155 = T156 < 13'ha1;
  assign T156 = sNatCAlignDist[4'hc:1'h0];
  assign CAlignDist_floor = isZeroProd | T157;
  assign T157 = sNatCAlignDist[4'hd:4'hd];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T158 == 3'h0;
  assign T158 = expB[4'hb:4'h9];
  assign isZeroA = T159 == 3'h0;
  assign T159 = expA[4'hb:4'h9];
  assign T160 = {T166, T161};
  assign T161 = {T165, T162};
  assign T162 = T163[1'h1:1'h1];
  assign T163 = T164[2'h3:2'h2];
  assign T164 = T143[2'h3:1'h0];
  assign T165 = T163[1'h0:1'h0];
  assign T166 = {T169, T167};
  assign T167 = T168[1'h1:1'h1];
  assign T168 = T164[1'h1:1'h0];
  assign T169 = T168[1'h0:1'h0];
  assign T170 = T193 | T171;
  assign T171 = T172 & 16'haaaa;
  assign T172 = T173 << 1'h1;
  assign T173 = T174[4'he:1'h0];
  assign T174 = T191 | T175;
  assign T175 = T176 & 16'hcccc;
  assign T176 = T177 << 2'h2;
  assign T177 = T178[4'hd:1'h0];
  assign T178 = T189 | T179;
  assign T179 = T180 & 16'hf0f0;
  assign T180 = T181 << 3'h4;
  assign T181 = T182[4'hb:1'h0];
  assign T182 = T187 | T183;
  assign T183 = T184 & 16'hff00;
  assign T184 = T185 << 4'h8;
  assign T185 = T186[3'h7:1'h0];
  assign T186 = T144[4'hf:1'h0];
  assign T187 = T750 & 16'hff;
  assign T750 = {8'h0, T188};
  assign T188 = T186 >> 4'h8;
  assign T189 = T751 & 16'hf0f;
  assign T751 = {4'h0, T190};
  assign T190 = T182 >> 3'h4;
  assign T191 = T752 & 16'h3333;
  assign T752 = {2'h0, T192};
  assign T192 = T178 >> 2'h2;
  assign T193 = T753 & 16'h5555;
  assign T753 = {1'h0, T194};
  assign T194 = T174 >> 1'h1;
  assign T195 = T224 | T196;
  assign T196 = T197 & 32'haaaaaaaa;
  assign T197 = T198 << 1'h1;
  assign T198 = T199[5'h1e:1'h0];
  assign T199 = T222 | T200;
  assign T200 = T201 & 32'hcccccccc;
  assign T201 = T202 << 2'h2;
  assign T202 = T203[5'h1d:1'h0];
  assign T203 = T220 | T204;
  assign T204 = T205 & 32'hf0f0f0f0;
  assign T205 = T206 << 3'h4;
  assign T206 = T207[5'h1b:1'h0];
  assign T207 = T218 | T208;
  assign T208 = T209 & 32'hff00ff00;
  assign T209 = T210 << 4'h8;
  assign T210 = T211[5'h17:1'h0];
  assign T211 = T216 | T212;
  assign T212 = T213 & 32'hffff0000;
  assign T213 = T214 << 5'h10;
  assign T214 = T215[4'hf:1'h0];
  assign T215 = T145[5'h1f:1'h0];
  assign T216 = T754 & 32'hffff;
  assign T754 = {16'h0, T217};
  assign T217 = T215 >> 5'h10;
  assign T218 = T755 & 32'hff00ff;
  assign T755 = {8'h0, T219};
  assign T219 = T211 >> 4'h8;
  assign T220 = T756 & 32'hf0f0f0f;
  assign T756 = {4'h0, T221};
  assign T221 = T207 >> 3'h4;
  assign T222 = T757 & 32'h33333333;
  assign T757 = {2'h0, T223};
  assign T223 = T203 >> 2'h2;
  assign T224 = T758 & 32'h55555555;
  assign T758 = {1'h0, T225};
  assign T225 = T199 >> 1'h1;
  assign sigC = {T226, fractC};
  assign fractC = io_c[6'h33:1'h0];
  assign T226 = isZeroC ^ 1'h1;
  assign isZeroC = T227 == 3'h0;
  assign T227 = expC[4'hb:4'h9];
  assign T228 = $signed(T229) >>> CAlignDist;
  assign T229 = T230;
  assign T230 = {doSubMags, T231};
  assign T231 = {negSigC, T232};
  assign T232 = 108'h0 - T759;
  assign T759 = {107'h0, doSubMags};
  assign negSigC = doSubMags ? T233 : sigC;
  assign T233 = ~ sigC;
  assign T760 = {55'h0, T234};
  assign T234 = T235 << 1'h1;
  assign T235 = sigA * sigB;
  assign sigB = {T236, fractB};
  assign fractB = io_b[6'h33:1'h0];
  assign T236 = isZeroB ^ 1'h1;
  assign sigA = {T237, fractA};
  assign fractA = io_a[6'h33:1'h0];
  assign T237 = isZeroA ^ 1'h1;
  assign T761 = {1'h0, T238};
  assign T238 = 108'h0 ^ T131;
  assign T239 = T128[2'h2:2'h2];
  assign T240 = T128[2'h3:2'h3];
  assign T241 = T128[3'h4:3'h4];
  assign T242 = T128[3'h5:3'h5];
  assign T243 = T128[3'h6:3'h6];
  assign T244 = T128[3'h7:3'h7];
  assign T245 = T128[4'h8:4'h8];
  assign T246 = T128[4'h9:4'h9];
  assign T247 = T128[4'ha:4'ha];
  assign T248 = T128[4'hb:4'hb];
  assign T249 = T128[4'hc:4'hc];
  assign T250 = T128[4'hd:4'hd];
  assign T251 = T128[4'he:4'he];
  assign T252 = T128[4'hf:4'hf];
  assign T253 = T128[5'h10:5'h10];
  assign T254 = T128[5'h11:5'h11];
  assign T255 = T128[5'h12:5'h12];
  assign T256 = T128[5'h13:5'h13];
  assign T257 = T128[5'h14:5'h14];
  assign T258 = T128[5'h15:5'h15];
  assign T259 = T128[5'h16:5'h16];
  assign T260 = T128[5'h17:5'h17];
  assign T261 = T128[5'h18:5'h18];
  assign T262 = T128[5'h19:5'h19];
  assign T263 = T128[5'h1a:5'h1a];
  assign T264 = T128[5'h1b:5'h1b];
  assign T265 = T128[5'h1c:5'h1c];
  assign T266 = T128[5'h1d:5'h1d];
  assign T267 = T128[5'h1e:5'h1e];
  assign T268 = T128[5'h1f:5'h1f];
  assign T269 = T128[6'h20:6'h20];
  assign T270 = T128[6'h21:6'h21];
  assign T271 = T128[6'h22:6'h22];
  assign T272 = T128[6'h23:6'h23];
  assign T273 = T128[6'h24:6'h24];
  assign T274 = T128[6'h25:6'h25];
  assign T275 = T128[6'h26:6'h26];
  assign T276 = T128[6'h27:6'h27];
  assign T277 = T128[6'h28:6'h28];
  assign T278 = T128[6'h29:6'h29];
  assign T279 = T128[6'h2a:6'h2a];
  assign T280 = T128[6'h2b:6'h2b];
  assign T281 = T128[6'h2c:6'h2c];
  assign T282 = T128[6'h2d:6'h2d];
  assign T283 = T128[6'h2e:6'h2e];
  assign T284 = T128[6'h2f:6'h2f];
  assign T285 = T128[6'h30:6'h30];
  assign T286 = T128[6'h31:6'h31];
  assign T287 = T128[6'h32:6'h32];
  assign T288 = T128[6'h33:6'h33];
  assign T289 = T128[6'h34:6'h34];
  assign T290 = T128[6'h35:6'h35];
  assign T291 = T128[6'h36:6'h36];
  assign T292 = T128[6'h37:6'h37];
  assign T293 = T128[6'h38:6'h38];
  assign T294 = T128[6'h39:6'h39];
  assign T295 = T128[6'h3a:6'h3a];
  assign T296 = T128[6'h3b:6'h3b];
  assign T297 = T128[6'h3c:6'h3c];
  assign T298 = T128[6'h3d:6'h3d];
  assign T299 = T128[6'h3e:6'h3e];
  assign T300 = T128[6'h3f:6'h3f];
  assign T301 = T128[7'h40:7'h40];
  assign T302 = T128[7'h41:7'h41];
  assign T303 = T128[7'h42:7'h42];
  assign T304 = T128[7'h43:7'h43];
  assign T305 = T128[7'h44:7'h44];
  assign T306 = T128[7'h45:7'h45];
  assign T307 = T128[7'h46:7'h46];
  assign T308 = T128[7'h47:7'h47];
  assign T309 = T128[7'h48:7'h48];
  assign T310 = T128[7'h49:7'h49];
  assign T311 = T128[7'h4a:7'h4a];
  assign T312 = T128[7'h4b:7'h4b];
  assign T313 = T128[7'h4c:7'h4c];
  assign T314 = T128[7'h4d:7'h4d];
  assign T315 = T128[7'h4e:7'h4e];
  assign T316 = T128[7'h4f:7'h4f];
  assign T317 = T128[7'h50:7'h50];
  assign T318 = T128[7'h51:7'h51];
  assign T319 = T128[7'h52:7'h52];
  assign T320 = T128[7'h53:7'h53];
  assign T321 = T128[7'h54:7'h54];
  assign T322 = T128[7'h55:7'h55];
  assign T323 = T128[7'h56:7'h56];
  assign T324 = T128[7'h57:7'h57];
  assign T325 = T128[7'h58:7'h58];
  assign T326 = T128[7'h59:7'h59];
  assign T327 = T128[7'h5a:7'h5a];
  assign T328 = T128[7'h5b:7'h5b];
  assign T329 = T128[7'h5c:7'h5c];
  assign T330 = T128[7'h5d:7'h5d];
  assign T331 = T128[7'h5e:7'h5e];
  assign T332 = T128[7'h5f:7'h5f];
  assign T333 = T128[7'h60:7'h60];
  assign T334 = T128[7'h61:7'h61];
  assign T335 = T128[7'h62:7'h62];
  assign T336 = T128[7'h63:7'h63];
  assign T337 = T128[7'h64:7'h64];
  assign T338 = T128[7'h65:7'h65];
  assign T339 = T128[7'h66:7'h66];
  assign T340 = T128[7'h67:7'h67];
  assign T341 = T128[7'h68:7'h68];
  assign T342 = T128[7'h69:7'h69];
  assign T343 = T128[7'h6a:7'h6a];
  assign T344 = T128[7'h6b:7'h6b];
  assign notCDom_signSigSum = sigSum[7'h6d:7'h6d];
  assign CDom_estNormDist = T347 ? CAlignDist : T762;
  assign T762 = {2'h0, T345};
  assign T345 = T346[3'h5:1'h0];
  assign T346 = CAlignDist - 8'h1;
  assign T347 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T348;
  assign T348 = T349 == 13'h0;
  assign T349 = sNatCAlignDist[4'hc:1'h0];
  assign isCDominant = T353 & T350;
  assign T350 = CAlignDist_floor | T351;
  assign T351 = T352 < 13'h36;
  assign T352 = sNatCAlignDist[4'hc:1'h0];
  assign T353 = isZeroC ^ 1'h1;
  assign sExpSum = CAlignDist_floor ? T763 : sExpAlignedProd;
  assign T763 = {2'h0, expC};
  assign T354 = T14[1'h0:1'h0];
  assign T355 = {T361, T356};
  assign T356 = {T360, T357};
  assign T357 = T358[1'h1:1'h1];
  assign T358 = T359[2'h3:2'h2];
  assign T359 = T15[2'h3:1'h0];
  assign T360 = T358[1'h0:1'h0];
  assign T361 = {T364, T362};
  assign T362 = T363[1'h1:1'h1];
  assign T363 = T359[1'h1:1'h0];
  assign T364 = T363[1'h0:1'h0];
  assign T365 = T388 | T366;
  assign T366 = T367 & 16'haaaa;
  assign T367 = T368 << 1'h1;
  assign T368 = T369[4'he:1'h0];
  assign T369 = T386 | T370;
  assign T370 = T371 & 16'hcccc;
  assign T371 = T372 << 2'h2;
  assign T372 = T373[4'hd:1'h0];
  assign T373 = T384 | T374;
  assign T374 = T375 & 16'hf0f0;
  assign T375 = T376 << 3'h4;
  assign T376 = T377[4'hb:1'h0];
  assign T377 = T382 | T378;
  assign T378 = T379 & 16'hff00;
  assign T379 = T380 << 4'h8;
  assign T380 = T381[3'h7:1'h0];
  assign T381 = T16[4'hf:1'h0];
  assign T382 = T764 & 16'hff;
  assign T764 = {8'h0, T383};
  assign T383 = T381 >> 4'h8;
  assign T384 = T765 & 16'hf0f;
  assign T765 = {4'h0, T385};
  assign T385 = T377 >> 3'h4;
  assign T386 = T766 & 16'h3333;
  assign T766 = {2'h0, T387};
  assign T387 = T373 >> 2'h2;
  assign T388 = T767 & 16'h5555;
  assign T767 = {1'h0, T389};
  assign T389 = T369 >> 1'h1;
  assign T390 = T419 | T391;
  assign T391 = T392 & 32'haaaaaaaa;
  assign T392 = T393 << 1'h1;
  assign T393 = T394[5'h1e:1'h0];
  assign T394 = T417 | T395;
  assign T395 = T396 & 32'hcccccccc;
  assign T396 = T397 << 2'h2;
  assign T397 = T398[5'h1d:1'h0];
  assign T398 = T415 | T399;
  assign T399 = T400 & 32'hf0f0f0f0;
  assign T400 = T401 << 3'h4;
  assign T401 = T402[5'h1b:1'h0];
  assign T402 = T413 | T403;
  assign T403 = T404 & 32'hff00ff00;
  assign T404 = T405 << 4'h8;
  assign T405 = T406[5'h17:1'h0];
  assign T406 = T411 | T407;
  assign T407 = T408 & 32'hffff0000;
  assign T408 = T409 << 5'h10;
  assign T409 = T410[4'hf:1'h0];
  assign T410 = T17[5'h1f:1'h0];
  assign T411 = T768 & 32'hffff;
  assign T768 = {16'h0, T412};
  assign T412 = T410 >> 5'h10;
  assign T413 = T769 & 32'hff00ff;
  assign T769 = {8'h0, T414};
  assign T414 = T406 >> 4'h8;
  assign T415 = T770 & 32'hf0f0f0f;
  assign T770 = {4'h0, T416};
  assign T416 = T402 >> 3'h4;
  assign T417 = T771 & 32'h33333333;
  assign T771 = {2'h0, T418};
  assign T418 = T398 >> 2'h2;
  assign T419 = T772 & 32'h55555555;
  assign T772 = {1'h0, T420};
  assign T420 = T394 >> 1'h1;
  assign T421 = 56'h0 - T773;
  assign T773 = {55'h0, T422};
  assign T422 = sExpX3[4'hd:4'hd];
  assign sigX3 = T423[6'h38:1'h0];
  assign T423 = {T595, T424};
  assign T424 = doIncrSig ? T591 : T425;
  assign T425 = T426 != 32'h0;
  assign T426 = T496 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T427, 1'h1};
  assign T427 = {T471, T428};
  assign T428 = {T452, T429};
  assign T429 = {T442, T430};
  assign T430 = {T438, T431};
  assign T431 = T432[2'h2:2'h2];
  assign T432 = T433[3'h6:3'h4];
  assign T433 = T434[4'he:4'h8];
  assign T434 = T435[5'h1e:5'h10];
  assign T435 = T436[5'h1f:1'h1];
  assign T436 = $signed(33'h100000000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T437;
  assign T437 = estNormDist[3'h4:1'h0];
  assign T438 = {T441, T439};
  assign T439 = T440[1'h1:1'h1];
  assign T440 = T432[1'h1:1'h0];
  assign T441 = T440[1'h0:1'h0];
  assign T442 = {T448, T443};
  assign T443 = {T447, T444};
  assign T444 = T445[1'h1:1'h1];
  assign T445 = T446[2'h3:2'h2];
  assign T446 = T433[2'h3:1'h0];
  assign T447 = T445[1'h0:1'h0];
  assign T448 = {T451, T449};
  assign T449 = T450[1'h1:1'h1];
  assign T450 = T446[1'h1:1'h0];
  assign T451 = T450[1'h0:1'h0];
  assign T452 = T469 | T453;
  assign T453 = T454 & 8'haa;
  assign T454 = T455 << 1'h1;
  assign T455 = T456[3'h6:1'h0];
  assign T456 = T467 | T457;
  assign T457 = T458 & 8'hcc;
  assign T458 = T459 << 2'h2;
  assign T459 = T460[3'h5:1'h0];
  assign T460 = T465 | T461;
  assign T461 = T462 & 8'hf0;
  assign T462 = T463 << 3'h4;
  assign T463 = T464[2'h3:1'h0];
  assign T464 = T434[3'h7:1'h0];
  assign T465 = T774 & 8'hf;
  assign T774 = {4'h0, T466};
  assign T466 = T464 >> 3'h4;
  assign T467 = T775 & 8'h33;
  assign T775 = {2'h0, T468};
  assign T468 = T460 >> 2'h2;
  assign T469 = T776 & 8'h55;
  assign T776 = {1'h0, T470};
  assign T470 = T456 >> 1'h1;
  assign T471 = T494 | T472;
  assign T472 = T473 & 16'haaaa;
  assign T473 = T474 << 1'h1;
  assign T474 = T475[4'he:1'h0];
  assign T475 = T492 | T476;
  assign T476 = T477 & 16'hcccc;
  assign T477 = T478 << 2'h2;
  assign T478 = T479[4'hd:1'h0];
  assign T479 = T490 | T480;
  assign T480 = T481 & 16'hf0f0;
  assign T481 = T482 << 3'h4;
  assign T482 = T483[4'hb:1'h0];
  assign T483 = T488 | T484;
  assign T484 = T485 & 16'hff00;
  assign T485 = T486 << 4'h8;
  assign T486 = T487[3'h7:1'h0];
  assign T487 = T435[4'hf:1'h0];
  assign T488 = T777 & 16'hff;
  assign T777 = {8'h0, T489};
  assign T489 = T487 >> 4'h8;
  assign T490 = T778 & 16'hf0f;
  assign T778 = {4'h0, T491};
  assign T491 = T483 >> 3'h4;
  assign T492 = T779 & 16'h3333;
  assign T779 = {2'h0, T493};
  assign T493 = T479 >> 2'h2;
  assign T494 = T780 & 16'h5555;
  assign T780 = {1'h0, T495};
  assign T495 = T475 >> 1'h1;
  assign T496 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T570 : T781;
  assign T781 = {1'h0, T497};
  assign T497 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T534 ? T522 : T498;
  assign T498 = T521 ? T502 : T499;
  assign T499 = {T501, T500};
  assign T500 = 54'h0 - T782;
  assign T782 = {53'h0, doSubMags};
  assign T501 = sigSum[6'h21:1'h1];
  assign T502 = T520 ? T784 : T503;
  assign T503 = {T505, T504};
  assign T504 = 86'h0 - T783;
  assign T783 = {85'h0, doSubMags};
  assign T505 = sigSum[1'h1:1'h1];
  assign T784 = {21'h0, T506};
  assign T506 = {T519, T507};
  assign T507 = doSubMags ? T513 : T508;
  assign T508 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T511, T509};
  assign T509 = T510 != 44'h0;
  assign T510 = sigSum[6'h2b:1'h0];
  assign T511 = T512 != 32'h0;
  assign T512 = sigSum[7'h4b:6'h2c];
  assign T513 = ~ T514;
  assign T514 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T517, T515};
  assign T515 = T516 != 44'h0;
  assign T516 = notSigSum[6'h2b:1'h0];
  assign notSigSum = ~ sigSum;
  assign T517 = T518 != 32'h0;
  assign T518 = notSigSum[7'h4b:6'h2c];
  assign T519 = sigSum[7'h6c:6'h2c];
  assign T520 = estNormNeg_dist[3'h4:3'h4];
  assign T521 = estNormNeg_dist[3'h5:3'h5];
  assign T522 = T533 ? T530 : T523;
  assign T523 = {T529, T524};
  assign T524 = doSubMags ? T527 : T525;
  assign T525 = T526 != 11'h0;
  assign T526 = sigSum[4'hb:1'h1];
  assign T527 = T528 == 11'h0;
  assign T528 = notSigSum[4'hb:1'h1];
  assign T529 = sigSum[7'h61:4'hc];
  assign T530 = {T532, T531};
  assign T531 = 22'h0 - T785;
  assign T785 = {21'h0, doSubMags};
  assign T532 = sigSum[7'h41:1'h1];
  assign T533 = estNormNeg_dist[3'h5:3'h5];
  assign T534 = estNormNeg_dist[3'h6:3'h6];
  assign CDom_firstNormAbsSigSum = T535;
  assign T535 = T543 | T536;
  assign T536 = T786 & T537;
  assign T537 = {T539, T538};
  assign T538 = firstReduceNotSigSum[1'h0:1'h0];
  assign T539 = notSigSum[8'h81:6'h2c];
  assign T786 = T540 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T540 = T541;
  assign T541 = doSubMags & T542;
  assign T542 = CDom_estNormDist[3'h5:3'h5];
  assign T543 = T552 | T544;
  assign T544 = T787 & T545;
  assign T545 = {T547, T546};
  assign T546 = firstReduceNotSigSum != 2'h0;
  assign T547 = notSigSum[8'ha1:7'h4c];
  assign T787 = T548 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T548 = T549;
  assign T549 = doSubMags & T550;
  assign T550 = ~ T551;
  assign T551 = CDom_estNormDist[3'h5:3'h5];
  assign T552 = T561 | T553;
  assign T553 = T788 & T554;
  assign T554 = {T556, T555};
  assign T555 = firstReduceSigSum[1'h0:1'h0];
  assign T556 = sigSum[8'h81:6'h2c];
  assign T788 = T557 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T557 = T558;
  assign T558 = T560 & T559;
  assign T559 = CDom_estNormDist[3'h5:3'h5];
  assign T560 = ~ doSubMags;
  assign T561 = T789 & T562;
  assign T562 = {T564, T563};
  assign T563 = firstReduceSigSum != 2'h0;
  assign T564 = sigSum[8'ha1:7'h4c];
  assign T789 = T565 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T565 = T566;
  assign T566 = T569 & T567;
  assign T567 = ~ T568;
  assign T568 = CDom_estNormDist[3'h5:3'h5];
  assign T569 = ~ doSubMags;
  assign T570 = isCDominant ? T791 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T590 ? T582 : T571;
  assign T571 = T581 ? T574 : T572;
  assign T572 = T573 << 6'h36;
  assign T573 = notSigSum[6'h22:1'h1];
  assign T574 = T580 ? T790 : T575;
  assign T575 = T576 << 7'h56;
  assign T576 = notSigSum[2'h2:1'h1];
  assign T790 = {23'h0, T577};
  assign T577 = {T579, T578};
  assign T578 = firstReduceNotSigSum[1'h0:1'h0];
  assign T579 = notSigSum[7'h6b:6'h2c];
  assign T580 = estNormNeg_dist[3'h4:3'h4];
  assign T581 = estNormNeg_dist[3'h5:3'h5];
  assign T582 = T589 ? T587 : T583;
  assign T583 = {T586, T584};
  assign T584 = T585 != 11'h0;
  assign T585 = notSigSum[4'hb:1'h1];
  assign T586 = notSigSum[7'h62:4'hc];
  assign T587 = T588 << 5'h16;
  assign T588 = notSigSum[7'h42:1'h1];
  assign T589 = estNormNeg_dist[3'h5:3'h5];
  assign T590 = estNormNeg_dist[3'h6:3'h6];
  assign T791 = {1'h0, CDom_firstNormAbsSigSum};
  assign T591 = T592 == 32'h0;
  assign T592 = T593 & absSigSumExtraMask;
  assign T593 = ~ T594;
  assign T594 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign T595 = T596 >> normTo2ShiftDist;
  assign T596 = cFirstNormAbsSigSum[7'h57:1'h1];
  assign roundPosBit = T597 != 57'h0;
  assign T597 = sigX3 & T792;
  assign T792 = {1'h0, roundPosMask};
  assign roundPosMask = T793 & roundMask;
  assign T793 = {1'h0, T598};
  assign T598 = ~ T599;
  assign T599 = roundMask >> 1'h1;
  assign T600 = ~ allRound;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T601 == 57'h0;
  assign T601 = T603 & T794;
  assign T794 = {2'h0, T602};
  assign T602 = roundMask >> 1'h1;
  assign T603 = ~ sigX3;
  assign doIncrSig = T604 & doSubMags;
  assign T604 = T606 & T605;
  assign T605 = ~ notCDom_signSigSum;
  assign T606 = ~ isCDominant;
  assign commonCase = T608 & T607;
  assign T607 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T608 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T609 == 2'h3;
  assign T609 = expC[4'hb:4'ha];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T610 == 2'h3;
  assign T610 = expB[4'hb:4'ha];
  assign isSpecialA = T611 == 2'h3;
  assign T611 = expA[4'hb:4'ha];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T612;
  assign T612 = T616 | T613;
  assign T613 = sExpX3_13 <= T795;
  assign T795 = {2'h0, T614};
  assign T614 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign sigX3Shift1 = T615 == 2'h0;
  assign T615 = sigX3[6'h38:6'h37];
  assign T616 = sExpX3[4'hd:4'hd];
  assign overflow = commonCase & overflowY;
  assign overflowY = T617 == 3'h3;
  assign T617 = sExpY[4'hc:4'ha];
  assign sExpY = T664 | T618;
  assign T618 = T620 ? T619 : 14'h0;
  assign T619 = sExpX3 - 14'h1;
  assign T620 = T621 == 2'h0;
  assign T621 = sigY3[6'h36:6'h35];
  assign sigY3 = T635 | T622;
  assign T622 = roundEven ? T623 : 55'h0;
  assign T623 = roundUp_sigY3 & T624;
  assign T624 = ~ T625;
  assign T625 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T626[6'h36:1'h0];
  assign T626 = T627 + 55'h1;
  assign T627 = T628 >> 2'h2;
  assign T628 = sigX3 | T796;
  assign T796 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T632 : T629;
  assign T629 = T631 & T630;
  assign T630 = ~ anyRoundExtra;
  assign T631 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T632 = T633 & allRoundExtra;
  assign T633 = roundingMode_nearest_even & T634;
  assign T634 = ~ roundPosBit;
  assign T635 = T657 | T636;
  assign T636 = roundUp ? roundUp_sigY3 : 55'h0;
  assign roundUp = T644 | T637;
  assign T637 = T638 & 1'h1;
  assign T638 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T642 & T639;
  assign T639 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T640 : notCDom_signSigSum;
  assign T640 = doSubMags & T641;
  assign T641 = ~ isZeroC;
  assign T642 = ~ isZeroY;
  assign isZeroY = T643 == 3'h0;
  assign T643 = sigX3[6'h38:6'h36];
  assign T644 = T647 | T645;
  assign T645 = T646 & roundPosBit;
  assign T646 = doIncrSig & roundingMode_nearest_even;
  assign T647 = T649 | T648;
  assign T648 = doIncrSig & allRound;
  assign T649 = T653 | T650;
  assign T650 = T651 & anyRound;
  assign T651 = T652 & roundDirectUp;
  assign T652 = ~ doIncrSig;
  assign T653 = T654 & anyRoundExtra;
  assign T654 = T655 & roundPosBit;
  assign T655 = T656 & roundingMode_nearest_even;
  assign T656 = ~ doIncrSig;
  assign T657 = T661 ? T658 : 55'h0;
  assign T658 = T659 >> 2'h2;
  assign T659 = sigX3 & T797;
  assign T797 = {1'h0, T660};
  assign T660 = ~ roundMask;
  assign T661 = T663 & T662;
  assign T662 = ~ roundEven;
  assign T663 = ~ roundUp;
  assign T664 = T667 | T665;
  assign T665 = T666 ? sExpX3 : 14'h0;
  assign T666 = sigY3[6'h35:6'h35];
  assign T667 = T669 ? T668 : 14'h0;
  assign T668 = sExpX3 + 14'h1;
  assign T669 = sigY3[6'h36:6'h36];
  assign T670 = {invalid, 1'h0};
  assign invalid = T689 | notSigNaN_invalid;
  assign notSigNaN_invalid = T686 | T671;
  assign T671 = T672 & doSubMags;
  assign T672 = T675 & isInfC;
  assign isInfC = isSpecialC & T673;
  assign T673 = T674 ^ 1'h1;
  assign T674 = expC[4'h9:4'h9];
  assign T675 = T681 & T676;
  assign T676 = isInfA | isInfB;
  assign isInfB = isSpecialB & T677;
  assign T677 = T678 ^ 1'h1;
  assign T678 = expB[4'h9:4'h9];
  assign isInfA = isSpecialA & T679;
  assign T679 = T680 ^ 1'h1;
  assign T680 = expA[4'h9:4'h9];
  assign T681 = T684 & T682;
  assign T682 = ~ isNaNB;
  assign isNaNB = isSpecialB & T683;
  assign T683 = expB[4'h9:4'h9];
  assign T684 = ~ isNaNA;
  assign isNaNA = isSpecialA & T685;
  assign T685 = expA[4'h9:4'h9];
  assign T686 = T688 | T687;
  assign T687 = isZeroA & isInfB;
  assign T688 = isInfA & isZeroB;
  assign T689 = T693 | isSigNaNC;
  assign isSigNaNC = isNaNC & T690;
  assign T690 = T691 ^ 1'h1;
  assign T691 = fractC[6'h33:6'h33];
  assign isNaNC = isSpecialC & T692;
  assign T692 = expC[4'h9:4'h9];
  assign T693 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T694;
  assign T694 = T695 ^ 1'h1;
  assign T695 = fractB[6'h33:6'h33];
  assign isSigNaNA = isNaNA & T696;
  assign T696 = T697 ^ 1'h1;
  assign T697 = fractA[6'h33:6'h33];
  assign io_out = T698;
  assign T698 = {signOut, T699};
  assign T699 = {expOut, fractOut};
  assign fractOut = fractY | T700;
  assign T700 = 52'h0 - T798;
  assign T798 = {51'h0, T701};
  assign T701 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T702;
  assign T702 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T705 | T703;
  assign T703 = roundingMode_max & T704;
  assign T704 = ~ signY;
  assign T705 = roundingMode_nearest_even | T706;
  assign T706 = roundingMode_min & signY;
  assign isNaNOut = T707 | notSigNaN_invalid;
  assign T707 = T708 | isNaNC;
  assign T708 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T710 : T709;
  assign T709 = sigY3[6'h34:1'h1];
  assign T710 = sigY3[6'h33:1'h0];
  assign expOut = T712 | T711;
  assign T711 = isNaNOut ? 12'he00 : 12'h0;
  assign T712 = T717 | T713;
  assign T713 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = T715 | T714;
  assign T714 = overflow & overflowY_roundMagUp;
  assign T715 = T716 | isInfC;
  assign T716 = isInfA | isInfB;
  assign T717 = T719 | T718;
  assign T718 = isSatOut ? 12'hbff : 12'h0;
  assign T719 = T722 & T720;
  assign T720 = ~ T721;
  assign T721 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T722 = T725 & T723;
  assign T723 = ~ T724;
  assign T724 = isSatOut ? 12'h400 : 12'h0;
  assign T725 = expY & T726;
  assign T726 = ~ T727;
  assign T727 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign notSpecial_isZeroOut = T731 | totalUnderflowY;
  assign totalUnderflowY = T730 | T728;
  assign T728 = T729 < 12'h3ce;
  assign T729 = sExpY[4'hb:1'h0];
  assign T730 = sExpY[4'hc:4'hc];
  assign T731 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'hb:1'h0];
  assign signOut = T733 | T732;
  assign T732 = commonCase & signY;
  assign T733 = T737 | T734;
  assign T734 = T735 & opSignC;
  assign T735 = T736 & isSpecialC;
  assign T736 = mulSpecial ^ 1'h1;
  assign T737 = T741 | T738;
  assign T738 = T739 & signProd;
  assign T739 = mulSpecial & T740;
  assign T740 = isSpecialC ^ 1'h1;
  assign T741 = T742 | isNaNOut;
  assign T742 = T743 & opSignC;
  assign T743 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_1(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T12;
  reg [2:0] in_rm;
  wire[2:0] T13;
  reg [64:0] in_in3;
  wire[64:0] T14;
  wire[64:0] T15;
  wire[64:0] zero;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg [64:0] in_in2;
  wire[64:0] T22;
  wire[64:0] T23;
  wire T24;
  reg [64:0] in_in1;
  wire[64:0] T25;
  wire[1:0] T26;
  reg [4:0] in_cmd;
  wire[4:0] T27;
  wire[4:0] T28;
  wire[4:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg [4:0] R0;
  wire[4:0] T1;
  reg [4:0] R2;
  wire[4:0] T3;
  wire[4:0] res_exc;
  reg  valid;
  reg  R4;
  wire T10;
  reg [64:0] R5;
  wire[64:0] T6;
  reg [64:0] R7;
  wire[64:0] T8;
  wire[64:0] res_data;
  reg  R9;
  wire T11;
  wire[64:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R0 = {1{$random}};
    R2 = {1{$random}};
    valid = {1{$random}};
    R4 = {1{$random}};
    R5 = {3{$random}};
    R7 = {3{$random}};
    R9 = {1{$random}};
  end
`endif

  assign T12 = in_rm[1'h1:1'h0];
  assign T13 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T14 = T19 ? zero : T15;
  assign T15 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign zero = T16 << 7'h40;
  assign T16 = T18 ^ T17;
  assign T17 = io_in_bits_in2[7'h40:7'h40];
  assign T18 = io_in_bits_in1[7'h40:7'h40];
  assign T19 = io_in_valid & T20;
  assign T20 = T21 ^ 1'h1;
  assign T21 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T22 = T24 ? 65'h8000000000000000 : T23;
  assign T23 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T24 = io_in_valid & io_in_bits_swap23;
  assign T25 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T26 = in_cmd[1'h1:1'h0];
  assign T27 = io_in_valid ? T29 : T28;
  assign T28 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T29 = {3'h0, T30};
  assign T30 = {T32, T31};
  assign T31 = io_in_bits_cmd[1'h0:1'h0];
  assign T32 = T34 & T33;
  assign T33 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T34 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R0;
  assign T1 = R4 ? R2 : R0;
  assign T3 = valid ? res_exc : R2;
  assign res_exc = fma_io_exceptionFlags;
  assign T10 = reset ? 1'h0 : valid;
  assign io_out_bits_data = R5;
  assign T6 = R4 ? R7 : R5;
  assign T8 = valid ? res_data : R7;
  assign res_data = fma_io_out;
  assign io_out_valid = R9;
  assign T11 = reset ? 1'h0 : R4;
  mulAddSubRecodedFloatN_1 fma(
       .io_op( T26 ),
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_c( in_in3 ),
       .io_roundingMode( T12 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T19) begin
      in_in3 <= zero;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T24) begin
      in_in2 <= 65'h8000000000000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T29;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(R4) begin
      R0 <= R2;
    end
    if(valid) begin
      R2 <= res_exc;
    end
    valid <= io_in_valid;
    if(reset) begin
      R4 <= 1'h0;
    end else begin
      R4 <= valid;
    end
    if(R4) begin
      R5 <= R7;
    end
    if(valid) begin
      R7 <= res_data;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else begin
      R9 <= R4;
    end
  end
endmodule

module recodedFloatNCompare(
    input [64:0] io_a,
    input [64:0] io_b,
    output io_a_eq_b,
    output io_a_lt_b,
    output io_a_eq_b_invalid,
    output io_a_lt_b_invalid
);

  wire T0;
  wire isNaNB;
  wire[2:0] codeB;
  wire[11:0] expB;
  wire isNaNA;
  wire[2:0] codeA;
  wire[11:0] expA;
  wire T1;
  wire isSignalingNaNB;
  wire T2;
  wire T3;
  wire[51:0] sigB;
  wire isSignalingNaNA;
  wire T4;
  wire T5;
  wire[51:0] sigA;
  wire T6;
  wire T7;
  wire T8;
  wire magLess;
  wire T9;
  wire T10;
  wire expEqual;
  wire T11;
  wire T12;
  wire T13;
  wire isZeroB;
  wire T14;
  wire isZeroA;
  wire T15;
  wire signA;
  wire T16;
  wire T17;
  wire magEqual;
  wire T18;
  wire T19;
  wire T20;
  wire signB;
  wire T21;
  wire T22;
  wire T23;
  wire signEqual;
  wire T24;
  wire T25;


  assign io_a_lt_b_invalid = T0;
  assign T0 = isNaNA | isNaNB;
  assign isNaNB = codeB == 3'h7;
  assign codeB = expB[4'hb:4'h9];
  assign expB = io_b[6'h3f:6'h34];
  assign isNaNA = codeA == 3'h7;
  assign codeA = expA[4'hb:4'h9];
  assign expA = io_a[6'h3f:6'h34];
  assign io_a_eq_b_invalid = T1;
  assign T1 = isSignalingNaNA | isSignalingNaNB;
  assign isSignalingNaNB = isNaNB & T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = sigB[6'h33:6'h33];
  assign sigB = io_b[6'h33:1'h0];
  assign isSignalingNaNA = isNaNA & T4;
  assign T4 = T5 ^ 1'h1;
  assign T5 = sigA[6'h33:6'h33];
  assign sigA = io_a[6'h33:1'h0];
  assign io_a_lt_b = T6;
  assign T6 = T21 & T7;
  assign T7 = signB ? T16 : T8;
  assign T8 = signA ? T12 : magLess;
  assign magLess = T11 | T9;
  assign T9 = expEqual & T10;
  assign T10 = sigA < sigB;
  assign expEqual = expA == expB;
  assign T11 = expA < expB;
  assign T12 = T13 ^ 1'h1;
  assign T13 = isZeroA & isZeroB;
  assign isZeroB = T14 ^ 1'h1;
  assign T14 = codeB != 3'h0;
  assign isZeroA = T15 ^ 1'h1;
  assign T15 = codeA != 3'h0;
  assign signA = io_a[7'h40:7'h40];
  assign T16 = T19 & T17;
  assign T17 = magEqual ^ 1'h1;
  assign magEqual = expEqual & T18;
  assign T18 = sigA == sigB;
  assign T19 = signA & T20;
  assign T20 = magLess ^ 1'h1;
  assign signB = io_b[7'h40:7'h40];
  assign T21 = io_a_lt_b_invalid ^ 1'h1;
  assign io_a_eq_b = T22;
  assign T22 = T24 & T23;
  assign T23 = isZeroA | signEqual;
  assign signEqual = signA == signB;
  assign T24 = T25 & magEqual;
  assign T25 = isNaNA ^ 1'h1;
endmodule

module FPToInt(input clk,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output io_out_bits_lt,
    output[63:0] io_out_bits_store,
    output[63:0] io_out_bits_toint,
    output[4:0] io_out_bits_exc
);

  reg [64:0] in_in2;
  wire[64:0] T346;
  wire[64:0] T347;
  wire[64:0] T348;
  wire[63:0] T349;
  wire[51:0] T350;
  wire[51:0] T351;
  wire[22:0] T352;
  wire[51:0] T353;
  wire[51:0] T354;
  wire T355;
  wire[2:0] T356;
  wire[11:0] T357;
  wire[11:0] T358;
  wire[11:0] T359;
  wire[11:0] T360;
  wire T361;
  wire[11:0] T362;
  wire[7:0] T363;
  wire T364;
  wire[11:0] T365;
  wire[10:0] T366;
  wire T367;
  wire[11:0] T368;
  wire T369;
  wire T370;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[4:0] T49;
  wire T50;
  wire T51;
  reg [64:0] in_in1;
  wire[64:0] T23;
  wire[64:0] T24;
  wire[64:0] T25;
  wire[63:0] T26;
  wire[51:0] T27;
  wire[51:0] T28;
  wire[22:0] T29;
  wire[51:0] T30;
  wire[51:0] T331;
  wire T31;
  wire[2:0] T32;
  wire[11:0] T33;
  wire[11:0] T34;
  wire[11:0] T35;
  wire[11:0] T36;
  wire T37;
  wire[11:0] T38;
  wire[7:0] T42;
  wire T39;
  wire[11:0] T332;
  wire[10:0] T40;
  wire T41;
  wire[11:0] T333;
  wire T43;
  wire T44;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] dcmp_exc;
  wire T2;
  wire[2:0] T3;
  wire[2:0] T330;
  wire[1:0] T4;
  wire[2:0] T5;
  reg [2:0] in_rm;
  wire[2:0] T6;
  wire T7;
  wire[4:0] T8;
  reg [4:0] in_cmd;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[3:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] T15;
  wire[2:0] T16;
  wire T17;
  wire[50:0] T18;
  wire[115:0] T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire[11:0] T22;
  wire T52;
  wire T53;
  wire[52:0] T54;
  wire[51:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[10:0] T66;
  wire T67;
  wire T68;
  wire[63:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[1:0] T87;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[10:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[1:0] T110;
  reg [1:0] in_typ;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[1:0] T127;
  wire T128;
  wire[4:0] T129;
  wire[63:0] T130;
  wire[63:0] T131;
  wire[63:0] T132;
  wire[63:0] unrec_out;
  wire[63:0] unrec_d;
  wire[62:0] T133;
  wire[51:0] T134;
  wire[51:0] T135;
  wire[51:0] T136;
  wire[52:0] T137;
  wire[5:0] T138;
  wire[5:0] T139;
  wire[11:0] T140;
  wire[52:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[9:0] T145;
  wire T146;
  wire[1:0] T147;
  wire T148;
  wire[2:0] T149;
  wire[51:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire[1:0] T162;
  wire[10:0] T163;
  wire[10:0] T164;
  wire[10:0] T334;
  wire[10:0] T165;
  wire[10:0] T166;
  wire T167;
  wire[63:0] T168;
  wire[31:0] unrec_s;
  wire[30:0] T169;
  wire[22:0] T170;
  wire[22:0] T171;
  wire[22:0] T172;
  wire[23:0] T173;
  wire[4:0] T174;
  wire[4:0] T175;
  wire[8:0] T176;
  wire[23:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire[6:0] T181;
  wire T182;
  wire[1:0] T183;
  wire T184;
  wire[2:0] T185;
  wire[22:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[1:0] T191;
  wire T192;
  wire T193;
  wire[1:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire[1:0] T198;
  wire[7:0] T199;
  wire[7:0] T200;
  wire[7:0] T335;
  wire[7:0] T201;
  wire[7:0] T202;
  wire T203;
  wire[31:0] T204;
  wire[31:0] T336;
  wire T205;
  reg  in_single;
  wire T206;
  wire[63:0] T337;
  wire[9:0] classify_out;
  wire[9:0] classify_d;
  wire[4:0] T207;
  wire[2:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[11:0] T215;
  wire T216;
  wire[1:0] T217;
  wire[2:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[9:0] T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[4:0] T237;
  wire[2:0] T238;
  wire[1:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire[1:0] T246;
  wire T247;
  wire T248;
  wire T249;
  wire[51:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire[9:0] classify_s;
  wire[4:0] T254;
  wire[2:0] T255;
  wire[1:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire[8:0] T262;
  wire T263;
  wire[1:0] T264;
  wire[2:0] T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire[6:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[1:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[4:0] T284;
  wire[2:0] T285;
  wire[1:0] T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[22:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire[63:0] T338;
  wire dcmp_out;
  wire[2:0] T302;
  wire[2:0] T339;
  wire[1:0] T303;
  wire[2:0] T304;
  wire[63:0] T305;
  wire[63:0] T340;
  wire[31:0] T306;
  wire[31:0] T307;
  wire[31:0] T341;
  wire T342;
  wire[63:0] T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] T312;
  wire[63:0] T313;
  wire T314;
  wire[63:0] T315;
  wire[63:0] T316;
  wire[63:0] T317;
  wire[63:0] T343;
  wire[31:0] T318;
  wire T319;
  wire T320;
  wire T321;
  wire[31:0] T344;
  wire T345;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg  valid;
  wire dcmp_io_a_eq_b;
  wire dcmp_io_a_lt_b;
  wire dcmp_io_a_eq_b_invalid;
  wire dcmp_io_a_lt_b_invalid;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_rm = {1{$random}};
    in_cmd = {1{$random}};
    in_typ = {1{$random}};
    in_single = {1{$random}};
    valid = {1{$random}};
  end
`endif

  assign T346 = T45 ? T348 : T347;
  assign T347 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T348 = {T370, T349};
  assign T349 = {T357, T350};
  assign T350 = T353 | T351;
  assign T351 = T352 << 5'h1d;
  assign T352 = io_in_bits_in2[5'h16:1'h0];
  assign T353 = 52'h0 - T354;
  assign T354 = {51'h0, T355};
  assign T355 = T356 == 3'h7;
  assign T356 = io_in_bits_in2[5'h1f:5'h1d];
  assign T357 = T369 ? T368 : T358;
  assign T358 = T367 ? T365 : T359;
  assign T359 = T364 ? T362 : T360;
  assign T360 = T361 ? 12'hc00 : 12'he00;
  assign T361 = T356 < 3'h7;
  assign T362 = {4'h8, T363};
  assign T363 = io_in_bits_in2[5'h1e:5'h17];
  assign T364 = T356 < 3'h6;
  assign T365 = {1'h0, T366};
  assign T366 = {3'h7, T363};
  assign T367 = T356 < 3'h4;
  assign T368 = {4'h0, T363};
  assign T369 = T356 < 3'h1;
  assign T370 = io_in_bits_in2[6'h20:6'h20];
  assign T45 = io_in_valid & T46;
  assign T46 = T50 & T47;
  assign T47 = T48 == 1'h0;
  assign T48 = T49 == 5'hc;
  assign T49 = io_in_bits_cmd & 5'hc;
  assign T50 = io_in_bits_single & T51;
  assign T51 = io_in_bits_ldst ^ 1'h1;
  assign T23 = T45 ? T25 : T24;
  assign T24 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T25 = {T44, T26};
  assign T26 = {T33, T27};
  assign T27 = T30 | T28;
  assign T28 = T29 << 5'h1d;
  assign T29 = io_in_bits_in1[5'h16:1'h0];
  assign T30 = 52'h0 - T331;
  assign T331 = {51'h0, T31};
  assign T31 = T32 == 3'h7;
  assign T32 = io_in_bits_in1[5'h1f:5'h1d];
  assign T33 = T43 ? T333 : T34;
  assign T34 = T41 ? T332 : T35;
  assign T35 = T39 ? T38 : T36;
  assign T36 = T37 ? 12'hc00 : 12'he00;
  assign T37 = T32 < 3'h7;
  assign T38 = {4'h8, T42};
  assign T42 = io_in_bits_in1[5'h1e:5'h17];
  assign T39 = T32 < 3'h6;
  assign T332 = {1'h0, T40};
  assign T40 = {3'h7, T42};
  assign T41 = T32 < 3'h4;
  assign T333 = {4'h0, T42};
  assign T43 = T32 < 3'h1;
  assign T44 = io_in_bits_in1[6'h20:6'h20];
  assign io_out_bits_exc = T0;
  assign T0 = T128 ? T10 : T1;
  assign T1 = T7 ? dcmp_exc : 5'h0;
  assign dcmp_exc = T2 << 3'h4;
  assign T2 = T3 != 3'h0;
  assign T3 = T5 & T330;
  assign T330 = {1'h0, T4};
  assign T4 = {dcmp_io_a_lt_b_invalid, dcmp_io_a_eq_b_invalid};
  assign T5 = ~ in_rm;
  assign T6 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T7 = T8 == 5'h4;
  assign T8 = in_cmd & 5'hc;
  assign T9 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T10 = {T58, T11};
  assign T11 = {3'h0, T12};
  assign T12 = T14 & T13;
  assign T13 = T58 ^ 1'h1;
  assign T14 = T15 != 2'h0;
  assign T15 = T16[1'h1:1'h0];
  assign T16 = {T57, T17};
  assign T17 = T18 != 51'h0;
  assign T18 = T19[6'h32:1'h0];
  assign T19 = T54 << T20;
  assign T20 = T52 ? 6'h0 : T21;
  assign T21 = T22[3'h5:1'h0];
  assign T22 = in_in1[6'h3f:6'h34];
  assign T52 = T53 ^ 1'h1;
  assign T53 = T22[4'hb:4'hb];
  assign T54 = {T56, T55};
  assign T55 = in_in1[6'h33:1'h0];
  assign T56 = T52 ^ 1'h1;
  assign T57 = T19[6'h34:6'h33];
  assign T58 = T126 | T59;
  assign T59 = T125 ? T119 : T60;
  assign T60 = T118 ? T112 : T61;
  assign T61 = T109 ? T103 : T62;
  assign T62 = T52 ? 1'h0 : T63;
  assign T63 = T102 ? T98 : T64;
  assign T64 = T97 ? T67 : T65;
  assign T65 = 11'h40 <= T66;
  assign T66 = T22[4'ha:1'h0];
  assign T67 = T70 | T68;
  assign T68 = T69 != 64'h0;
  assign T69 = T19[7'h73:6'h34];
  assign T70 = T96 | T71;
  assign T71 = T95 ? T84 : T72;
  assign T72 = T83 ? T82 : T73;
  assign T73 = T81 ? T74 : 1'h0;
  assign T74 = T79 & T75;
  assign T75 = T52 ? T76 : T14;
  assign T76 = T77 ^ 1'h1;
  assign T77 = T78 == 3'h0;
  assign T78 = T22[4'hb:4'h9];
  assign T79 = T80 ^ 1'h1;
  assign T80 = in_in1[7'h40:7'h40];
  assign T81 = in_rm == 3'h3;
  assign T82 = T80 & T75;
  assign T83 = in_rm == 3'h2;
  assign T84 = T52 ? T90 : T85;
  assign T85 = T88 | T86;
  assign T86 = T87 == 2'h3;
  assign T87 = T16[1'h1:1'h0];
  assign T88 = T89 == 2'h3;
  assign T89 = T16[2'h2:1'h1];
  assign T90 = T91 & T14;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T94 == 11'h7ff;
  assign T94 = T22[4'ha:1'h0];
  assign T95 = in_rm == 3'h0;
  assign T96 = T80 ^ 1'h1;
  assign T97 = T66 == 11'h3f;
  assign T98 = T101 & T99;
  assign T99 = T71 & T100;
  assign T100 = T69 == 64'hffffffffffffffff;
  assign T101 = T80 ^ 1'h1;
  assign T102 = T66 == 11'h3e;
  assign T103 = T52 ? T108 : T104;
  assign T104 = T80 | T105;
  assign T105 = T107 ? T99 : T106;
  assign T106 = 11'h40 <= T66;
  assign T107 = T66 == 11'h3f;
  assign T108 = T80 & T71;
  assign T109 = T110 == 2'h2;
  assign T110 = in_typ ^ 2'h1;
  assign T111 = io_in_valid ? io_in_bits_typ : in_typ;
  assign T112 = T52 ? 1'h0 : T113;
  assign T113 = T117 ? T98 : T114;
  assign T114 = T116 ? T67 : T115;
  assign T115 = 11'h20 <= T66;
  assign T116 = T66 == 11'h1f;
  assign T117 = T66 == 11'h1e;
  assign T118 = T110 == 2'h1;
  assign T119 = T52 ? T124 : T120;
  assign T120 = T80 | T121;
  assign T121 = T123 ? T99 : T122;
  assign T122 = 11'h20 <= T66;
  assign T123 = T66 == 11'h1f;
  assign T124 = T80 & T71;
  assign T125 = T110 == 2'h0;
  assign T126 = T127 == 2'h3;
  assign T127 = T22[4'hb:4'ha];
  assign T128 = T129 == 5'h8;
  assign T129 = in_cmd & 5'hc;
  assign io_out_bits_toint = T130;
  assign T130 = T128 ? T305 : T131;
  assign T131 = T7 ? T338 : T132;
  assign T132 = T301 ? T337 : unrec_out;
  assign unrec_out = in_single ? T168 : unrec_d;
  assign unrec_d = {T167, T133};
  assign T133 = {T163, T134};
  assign T134 = T151 ? T150 : T135;
  assign T135 = T142 ? T136 : 52'h0;
  assign T136 = T137[6'h33:1'h0];
  assign T137 = T141 >> T138;
  assign T138 = 6'h2 - T139;
  assign T139 = T140[3'h5:1'h0];
  assign T140 = in_in1[6'h3f:6'h34];
  assign T141 = {1'h1, T150};
  assign T142 = T148 | T143;
  assign T143 = T146 & T144;
  assign T144 = T145 < 10'h2;
  assign T145 = T140[4'h9:1'h0];
  assign T146 = T147 == 2'h1;
  assign T147 = T140[4'hb:4'ha];
  assign T148 = T149 == 3'h1;
  assign T149 = T140[4'hb:4'h9];
  assign T150 = in_in1[6'h33:1'h0];
  assign T151 = T156 | T152;
  assign T152 = T154 & T153;
  assign T153 = T140[4'h9:4'h9];
  assign T154 = T155 == 2'h3;
  assign T155 = T140[4'hb:4'ha];
  assign T156 = T159 | T157;
  assign T157 = T158 == 2'h2;
  assign T158 = T140[4'hb:4'ha];
  assign T159 = T161 & T160;
  assign T160 = T144 ^ 1'h1;
  assign T161 = T162 == 2'h1;
  assign T162 = T140[4'hb:4'ha];
  assign T163 = T156 ? T165 : T164;
  assign T164 = 11'h0 - T334;
  assign T334 = {10'h0, T154};
  assign T165 = T166 - 11'h401;
  assign T166 = T140[4'ha:1'h0];
  assign T167 = in_in1[7'h40:7'h40];
  assign T168 = {T204, unrec_s};
  assign unrec_s = {T203, T169};
  assign T169 = {T199, T170};
  assign T170 = T187 ? T186 : T171;
  assign T171 = T178 ? T172 : 23'h0;
  assign T172 = T173[5'h16:1'h0];
  assign T173 = T177 >> T174;
  assign T174 = 5'h2 - T175;
  assign T175 = T176[3'h4:1'h0];
  assign T176 = in_in1[5'h1f:5'h17];
  assign T177 = {1'h1, T186};
  assign T178 = T184 | T179;
  assign T179 = T182 & T180;
  assign T180 = T181 < 7'h2;
  assign T181 = T176[3'h6:1'h0];
  assign T182 = T183 == 2'h1;
  assign T183 = T176[4'h8:3'h7];
  assign T184 = T185 == 3'h1;
  assign T185 = T176[4'h8:3'h6];
  assign T186 = in_in1[5'h16:1'h0];
  assign T187 = T192 | T188;
  assign T188 = T190 & T189;
  assign T189 = T176[3'h6:3'h6];
  assign T190 = T191 == 2'h3;
  assign T191 = T176[4'h8:3'h7];
  assign T192 = T195 | T193;
  assign T193 = T194 == 2'h2;
  assign T194 = T176[4'h8:3'h7];
  assign T195 = T197 & T196;
  assign T196 = T180 ^ 1'h1;
  assign T197 = T198 == 2'h1;
  assign T198 = T176[4'h8:3'h7];
  assign T199 = T192 ? T201 : T200;
  assign T200 = 8'h0 - T335;
  assign T335 = {7'h0, T190};
  assign T201 = T202 - 8'h81;
  assign T202 = T176[3'h7:1'h0];
  assign T203 = in_in1[6'h20:6'h20];
  assign T204 = 32'h0 - T336;
  assign T336 = {31'h0, T205};
  assign T205 = unrec_s[5'h1f:5'h1f];
  assign T206 = io_in_valid ? io_in_bits_single : in_single;
  assign T337 = {54'h0, classify_out};
  assign classify_out = in_single ? classify_s : classify_d;
  assign classify_d = {T237, T207};
  assign T207 = {T232, T208};
  assign T208 = {T227, T209};
  assign T209 = {T219, T210};
  assign T210 = T212 & T211;
  assign T211 = in_in1[7'h40:7'h40];
  assign T212 = T216 & T213;
  assign T213 = T214 ^ 1'h1;
  assign T214 = T215[4'h9:4'h9];
  assign T215 = in_in1[6'h3f:6'h34];
  assign T216 = T217 == 2'h3;
  assign T217 = T218[2'h2:1'h1];
  assign T218 = T215[4'hb:4'h9];
  assign T219 = T220 & T211;
  assign T220 = T222 | T221;
  assign T221 = T217 == 2'h2;
  assign T222 = T226 & T223;
  assign T223 = T224 ^ 1'h1;
  assign T224 = T225 < 10'h2;
  assign T225 = T215[4'h9:1'h0];
  assign T226 = T217 == 2'h1;
  assign T227 = T228 & T211;
  assign T228 = T231 | T229;
  assign T229 = T230 & T224;
  assign T230 = T217 == 2'h1;
  assign T231 = T218 == 3'h1;
  assign T232 = {T235, T233};
  assign T233 = T234 & T211;
  assign T234 = T218 == 3'h0;
  assign T235 = T234 & T236;
  assign T236 = T211 ^ 1'h1;
  assign T237 = {T246, T238};
  assign T238 = {T244, T239};
  assign T239 = {T242, T240};
  assign T240 = T228 & T241;
  assign T241 = T211 ^ 1'h1;
  assign T242 = T220 & T243;
  assign T243 = T211 ^ 1'h1;
  assign T244 = T212 & T245;
  assign T245 = T211 ^ 1'h1;
  assign T246 = {T252, T247};
  assign T247 = T251 & T248;
  assign T248 = T249 ^ 1'h1;
  assign T249 = T250[6'h33:6'h33];
  assign T250 = in_in1[6'h33:1'h0];
  assign T251 = T218 == 3'h7;
  assign T252 = T251 & T253;
  assign T253 = T250[6'h33:6'h33];
  assign classify_s = {T284, T254};
  assign T254 = {T279, T255};
  assign T255 = {T274, T256};
  assign T256 = {T266, T257};
  assign T257 = T259 & T258;
  assign T258 = in_in1[6'h20:6'h20];
  assign T259 = T263 & T260;
  assign T260 = T261 ^ 1'h1;
  assign T261 = T262[3'h6:3'h6];
  assign T262 = in_in1[5'h1f:5'h17];
  assign T263 = T264 == 2'h3;
  assign T264 = T265[2'h2:1'h1];
  assign T265 = T262[4'h8:3'h6];
  assign T266 = T267 & T258;
  assign T267 = T269 | T268;
  assign T268 = T264 == 2'h2;
  assign T269 = T273 & T270;
  assign T270 = T271 ^ 1'h1;
  assign T271 = T272 < 7'h2;
  assign T272 = T262[3'h6:1'h0];
  assign T273 = T264 == 2'h1;
  assign T274 = T275 & T258;
  assign T275 = T278 | T276;
  assign T276 = T277 & T271;
  assign T277 = T264 == 2'h1;
  assign T278 = T265 == 3'h1;
  assign T279 = {T282, T280};
  assign T280 = T281 & T258;
  assign T281 = T265 == 3'h0;
  assign T282 = T281 & T283;
  assign T283 = T258 ^ 1'h1;
  assign T284 = {T293, T285};
  assign T285 = {T291, T286};
  assign T286 = {T289, T287};
  assign T287 = T275 & T288;
  assign T288 = T258 ^ 1'h1;
  assign T289 = T267 & T290;
  assign T290 = T258 ^ 1'h1;
  assign T291 = T259 & T292;
  assign T292 = T258 ^ 1'h1;
  assign T293 = {T299, T294};
  assign T294 = T298 & T295;
  assign T295 = T296 ^ 1'h1;
  assign T296 = T297[5'h16:5'h16];
  assign T297 = in_in1[5'h16:1'h0];
  assign T298 = T265 == 3'h7;
  assign T299 = T298 & T300;
  assign T300 = T297[5'h16:5'h16];
  assign T301 = in_rm[1'h0:1'h0];
  assign T338 = {63'h0, dcmp_out};
  assign dcmp_out = T302 != 3'h0;
  assign T302 = T304 & T339;
  assign T339 = {1'h0, T303};
  assign T303 = {dcmp_io_a_lt_b, dcmp_io_a_eq_b};
  assign T304 = ~ in_rm;
  assign T305 = T329 ? T308 : T340;
  assign T340 = {T341, T306};
  assign T306 = T307;
  assign T307 = T308[5'h1f:1'h0];
  assign T341 = T342 ? 32'hffffffff : 32'h0;
  assign T342 = T306[5'h1f:5'h1f];
  assign T308 = T58 ? T315 : T309;
  assign T309 = T310;
  assign T310 = T314 ? T313 : T311;
  assign T311 = T80 ? T312 : T69;
  assign T312 = ~ T69;
  assign T313 = T311 + 64'h1;
  assign T314 = T71 ^ T80;
  assign T315 = T327 ? 64'h8000000000000000 : T316;
  assign T316 = T325 ? 64'hffffffff80000000 : T317;
  assign T317 = T322 ? 64'h7fffffffffffffff : T343;
  assign T343 = {T344, T318};
  assign T318 = T319 ? 32'h7fffffff : 32'hffffffff;
  assign T319 = T321 & T320;
  assign T320 = T80 ^ 1'h1;
  assign T321 = T110 == 2'h1;
  assign T344 = T345 ? 32'hffffffff : 32'h0;
  assign T345 = T318[5'h1f:5'h1f];
  assign T322 = T324 & T323;
  assign T323 = T80 ^ 1'h1;
  assign T324 = T110 == 2'h3;
  assign T325 = T326 & T80;
  assign T326 = T110 == 2'h1;
  assign T327 = T328 & T80;
  assign T328 = T110 == 2'h3;
  assign T329 = in_typ[1'h1:1'h1];
  assign io_out_bits_store = unrec_out;
  assign io_out_bits_lt = dcmp_io_a_lt_b;
  assign io_out_valid = valid;
  recodedFloatNCompare dcmp(
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_a_eq_b( dcmp_io_a_eq_b ),
       .io_a_lt_b( dcmp_io_a_lt_b ),
       .io_a_eq_b_invalid( dcmp_io_a_eq_b_invalid ),
       .io_a_lt_b_invalid( dcmp_io_a_lt_b_invalid )
  );

  always @(posedge clk) begin
    if(T45) begin
      in_in2 <= T348;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(T45) begin
      in_in1 <= T25;
    end else if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      in_single <= io_in_bits_single;
    end
    valid <= io_in_valid;
  end
endmodule

module IntToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  reg [4:0] R0;
  wire[4:0] T1;
  reg [4:0] R2;
  wire[4:0] T3;
  wire[4:0] mux_exc;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[1:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[38:0] T12;
  wire[126:0] T13;
  wire[5:0] T14;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[5:0] T216;
  wire[5:0] T217;
  wire[5:0] T218;
  wire[5:0] T219;
  wire[5:0] T220;
  wire[5:0] T221;
  wire[5:0] T222;
  wire[5:0] T223;
  wire[5:0] T224;
  wire[5:0] T225;
  wire[5:0] T226;
  wire[5:0] T227;
  wire[5:0] T228;
  wire[5:0] T229;
  wire[5:0] T230;
  wire[5:0] T231;
  wire[5:0] T232;
  wire[5:0] T233;
  wire[5:0] T234;
  wire[5:0] T235;
  wire[5:0] T236;
  wire[5:0] T237;
  wire[5:0] T238;
  wire[4:0] T239;
  wire[4:0] T240;
  wire[4:0] T241;
  wire[4:0] T242;
  wire[4:0] T243;
  wire[4:0] T244;
  wire[4:0] T245;
  wire[4:0] T246;
  wire[4:0] T247;
  wire[4:0] T248;
  wire[4:0] T249;
  wire[4:0] T250;
  wire[4:0] T251;
  wire[4:0] T252;
  wire[4:0] T253;
  wire[4:0] T254;
  wire[3:0] T255;
  wire[3:0] T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[3:0] T262;
  wire[2:0] T263;
  wire[2:0] T264;
  wire[2:0] T265;
  wire[2:0] T266;
  wire[1:0] T267;
  wire[1:0] T268;
  wire T269;
  wire[63:0] T16;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[63:0] T17;
  wire[63:0] T332;
  wire[31:0] T18;
  wire[63:0] T19;
  wire[63:0] T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire[63:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  reg [1:0] R29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  reg  R38;
  wire T39;
  wire T40;
  wire[4:0] T41;
  reg [4:0] R42;
  wire[4:0] T43;
  wire[4:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire[2:0] T48;
  wire T49;
  wire[9:0] T50;
  wire[126:0] T51;
  wire[5:0] T52;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[5:0] T343;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[5:0] T349;
  wire[5:0] T350;
  wire[5:0] T351;
  wire[5:0] T352;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[5:0] T357;
  wire[5:0] T358;
  wire[5:0] T359;
  wire[5:0] T360;
  wire[5:0] T361;
  wire[5:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[4:0] T365;
  wire[4:0] T366;
  wire[4:0] T367;
  wire[4:0] T368;
  wire[4:0] T369;
  wire[4:0] T370;
  wire[4:0] T371;
  wire[4:0] T372;
  wire[4:0] T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire[4:0] T377;
  wire[4:0] T378;
  wire[4:0] T379;
  wire[4:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] T383;
  wire[3:0] T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[2:0] T389;
  wire[2:0] T390;
  wire[2:0] T391;
  wire[2:0] T392;
  wire[1:0] T393;
  wire[1:0] T394;
  wire T395;
  wire[63:0] T54;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire[63:0] T55;
  wire[63:0] T458;
  wire[31:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[1:0] T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T459;
  reg  R74;
  wire T460;
  reg [64:0] R75;
  wire[64:0] T76;
  reg [64:0] R77;
  wire[64:0] T78;
  wire[64:0] mux_data;
  wire[64:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[64:0] T82;
  wire[63:0] T83;
  wire[51:0] T84;
  wire[51:0] T85;
  wire[51:0] T86;
  wire[126:0] T87;
  wire[5:0] T88;
  wire[5:0] T461;
  wire[5:0] T462;
  wire[5:0] T463;
  wire[5:0] T464;
  wire[5:0] T465;
  wire[5:0] T466;
  wire[5:0] T467;
  wire[5:0] T468;
  wire[5:0] T469;
  wire[5:0] T470;
  wire[5:0] T471;
  wire[5:0] T472;
  wire[5:0] T473;
  wire[5:0] T474;
  wire[5:0] T475;
  wire[5:0] T476;
  wire[5:0] T477;
  wire[5:0] T478;
  wire[5:0] T479;
  wire[5:0] T480;
  wire[5:0] T481;
  wire[5:0] T482;
  wire[5:0] T483;
  wire[5:0] T484;
  wire[5:0] T485;
  wire[5:0] T486;
  wire[5:0] T487;
  wire[5:0] T488;
  wire[5:0] T489;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[5:0] T492;
  wire[4:0] T493;
  wire[4:0] T494;
  wire[4:0] T495;
  wire[4:0] T496;
  wire[4:0] T497;
  wire[4:0] T498;
  wire[4:0] T499;
  wire[4:0] T500;
  wire[4:0] T501;
  wire[4:0] T502;
  wire[4:0] T503;
  wire[4:0] T504;
  wire[4:0] T505;
  wire[4:0] T506;
  wire[4:0] T507;
  wire[4:0] T508;
  wire[3:0] T509;
  wire[3:0] T510;
  wire[3:0] T511;
  wire[3:0] T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[3:0] T516;
  wire[2:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire[2:0] T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire T523;
  wire[63:0] T90;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[63:0] T91;
  wire T92;
  wire[10:0] T93;
  wire[11:0] T94;
  wire[11:0] T586;
  wire[9:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[11:0] T101;
  wire[11:0] T587;
  wire[10:0] T102;
  wire[10:0] T103;
  wire[10:0] T588;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[11:0] T108;
  wire[11:0] T589;
  wire[11:0] T109;
  wire[11:0] T110;
  wire[5:0] T111;
  wire T112;
  wire[64:0] T113;
  wire[32:0] T114;
  wire[31:0] T115;
  wire[22:0] T116;
  wire[22:0] T117;
  wire[22:0] T118;
  wire[62:0] T119;
  wire[4:0] T120;
  wire[4:0] T590;
  wire[4:0] T591;
  wire[4:0] T592;
  wire[4:0] T593;
  wire[4:0] T594;
  wire[4:0] T595;
  wire[4:0] T596;
  wire[4:0] T597;
  wire[4:0] T598;
  wire[4:0] T599;
  wire[4:0] T600;
  wire[4:0] T601;
  wire[4:0] T602;
  wire[4:0] T603;
  wire[4:0] T604;
  wire[4:0] T605;
  wire[3:0] T606;
  wire[3:0] T607;
  wire[3:0] T608;
  wire[3:0] T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[3:0] T612;
  wire[3:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire[2:0] T616;
  wire[2:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire T620;
  wire[31:0] T122;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire[31:0] T123;
  wire T124;
  wire[7:0] T125;
  wire[8:0] T126;
  wire[8:0] T651;
  wire[6:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  wire[8:0] T133;
  wire[8:0] T652;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T653;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire[8:0] T140;
  wire[8:0] T654;
  wire[8:0] T141;
  wire[8:0] T142;
  wire[4:0] T143;
  wire T144;
  wire[64:0] T145;
  wire[32:0] T146;
  wire[31:0] T147;
  wire[22:0] T148;
  wire[24:0] T149;
  wire[24:0] T150;
  wire[23:0] T151;
  wire[24:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  reg [2:0] R159;
  wire[2:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire[1:0] T167;
  wire T168;
  wire[8:0] T169;
  wire[7:0] T170;
  wire[7:0] T171;
  wire[7:0] T655;
  wire T172;
  wire[7:0] T173;
  wire[6:0] T174;
  wire[5:0] T175;
  wire T176;
  wire[64:0] T177;
  wire[63:0] T178;
  wire[51:0] T179;
  wire[53:0] T180;
  wire[53:0] T181;
  wire[52:0] T182;
  wire[53:0] T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[1:0] T194;
  wire T195;
  wire[1:0] T196;
  wire T197;
  wire[11:0] T198;
  wire[10:0] T199;
  wire[10:0] T200;
  wire[10:0] T656;
  wire T201;
  wire[10:0] T202;
  wire[9:0] T203;
  wire[5:0] T204;
  wire T205;
  reg  R206;
  wire T657;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R2 = {1{$random}};
    R21 = {3{$random}};
    R29 = {1{$random}};
    R38 = {1{$random}};
    R42 = {1{$random}};
    R73 = {1{$random}};
    R74 = {1{$random}};
    R75 = {3{$random}};
    R77 = {3{$random}};
    R159 = {1{$random}};
    R206 = {1{$random}};
  end
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R74 ? R2 : R0;
  assign T3 = R73 ? mux_exc : R2;
  assign mux_exc = T4;
  assign T4 = T71 ? T44 : T5;
  assign T5 = T37 ? T6 : 5'h0;
  assign T6 = {3'h0, T7};
  assign T7 = {1'h0, T8};
  assign T8 = T9 != 2'h0;
  assign T9 = T10[1'h1:1'h0];
  assign T10 = {T36, T11};
  assign T11 = T12 != 39'h0;
  assign T12 = T13[6'h26:1'h0];
  assign T13 = T17 << T14;
  assign T14 = ~ T207;
  assign T207 = T331 ? 6'h3f : T208;
  assign T208 = T330 ? 6'h3e : T209;
  assign T209 = T329 ? 6'h3d : T210;
  assign T210 = T328 ? 6'h3c : T211;
  assign T211 = T327 ? 6'h3b : T212;
  assign T212 = T326 ? 6'h3a : T213;
  assign T213 = T325 ? 6'h39 : T214;
  assign T214 = T324 ? 6'h38 : T215;
  assign T215 = T323 ? 6'h37 : T216;
  assign T216 = T322 ? 6'h36 : T217;
  assign T217 = T321 ? 6'h35 : T218;
  assign T218 = T320 ? 6'h34 : T219;
  assign T219 = T319 ? 6'h33 : T220;
  assign T220 = T318 ? 6'h32 : T221;
  assign T221 = T317 ? 6'h31 : T222;
  assign T222 = T316 ? 6'h30 : T223;
  assign T223 = T315 ? 6'h2f : T224;
  assign T224 = T314 ? 6'h2e : T225;
  assign T225 = T313 ? 6'h2d : T226;
  assign T226 = T312 ? 6'h2c : T227;
  assign T227 = T311 ? 6'h2b : T228;
  assign T228 = T310 ? 6'h2a : T229;
  assign T229 = T309 ? 6'h29 : T230;
  assign T230 = T308 ? 6'h28 : T231;
  assign T231 = T307 ? 6'h27 : T232;
  assign T232 = T306 ? 6'h26 : T233;
  assign T233 = T305 ? 6'h25 : T234;
  assign T234 = T304 ? 6'h24 : T235;
  assign T235 = T303 ? 6'h23 : T236;
  assign T236 = T302 ? 6'h22 : T237;
  assign T237 = T301 ? 6'h21 : T238;
  assign T238 = T300 ? 6'h20 : T239;
  assign T239 = T299 ? 5'h1f : T240;
  assign T240 = T298 ? 5'h1e : T241;
  assign T241 = T297 ? 5'h1d : T242;
  assign T242 = T296 ? 5'h1c : T243;
  assign T243 = T295 ? 5'h1b : T244;
  assign T244 = T294 ? 5'h1a : T245;
  assign T245 = T293 ? 5'h19 : T246;
  assign T246 = T292 ? 5'h18 : T247;
  assign T247 = T291 ? 5'h17 : T248;
  assign T248 = T290 ? 5'h16 : T249;
  assign T249 = T289 ? 5'h15 : T250;
  assign T250 = T288 ? 5'h14 : T251;
  assign T251 = T287 ? 5'h13 : T252;
  assign T252 = T286 ? 5'h12 : T253;
  assign T253 = T285 ? 5'h11 : T254;
  assign T254 = T284 ? 5'h10 : T255;
  assign T255 = T283 ? 4'hf : T256;
  assign T256 = T282 ? 4'he : T257;
  assign T257 = T281 ? 4'hd : T258;
  assign T258 = T280 ? 4'hc : T259;
  assign T259 = T279 ? 4'hb : T260;
  assign T260 = T278 ? 4'ha : T261;
  assign T261 = T277 ? 4'h9 : T262;
  assign T262 = T276 ? 4'h8 : T263;
  assign T263 = T275 ? 3'h7 : T264;
  assign T264 = T274 ? 3'h6 : T265;
  assign T265 = T273 ? 3'h5 : T266;
  assign T266 = T272 ? 3'h4 : T267;
  assign T267 = T271 ? 2'h3 : T268;
  assign T268 = T270 ? 2'h2 : T269;
  assign T269 = T16[1'h1:1'h1];
  assign T16 = T17[6'h3f:1'h0];
  assign T270 = T16[2'h2:2'h2];
  assign T271 = T16[2'h3:2'h3];
  assign T272 = T16[3'h4:3'h4];
  assign T273 = T16[3'h5:3'h5];
  assign T274 = T16[3'h6:3'h6];
  assign T275 = T16[3'h7:3'h7];
  assign T276 = T16[4'h8:4'h8];
  assign T277 = T16[4'h9:4'h9];
  assign T278 = T16[4'ha:4'ha];
  assign T279 = T16[4'hb:4'hb];
  assign T280 = T16[4'hc:4'hc];
  assign T281 = T16[4'hd:4'hd];
  assign T282 = T16[4'he:4'he];
  assign T283 = T16[4'hf:4'hf];
  assign T284 = T16[5'h10:5'h10];
  assign T285 = T16[5'h11:5'h11];
  assign T286 = T16[5'h12:5'h12];
  assign T287 = T16[5'h13:5'h13];
  assign T288 = T16[5'h14:5'h14];
  assign T289 = T16[5'h15:5'h15];
  assign T290 = T16[5'h16:5'h16];
  assign T291 = T16[5'h17:5'h17];
  assign T292 = T16[5'h18:5'h18];
  assign T293 = T16[5'h19:5'h19];
  assign T294 = T16[5'h1a:5'h1a];
  assign T295 = T16[5'h1b:5'h1b];
  assign T296 = T16[5'h1c:5'h1c];
  assign T297 = T16[5'h1d:5'h1d];
  assign T298 = T16[5'h1e:5'h1e];
  assign T299 = T16[5'h1f:5'h1f];
  assign T300 = T16[6'h20:6'h20];
  assign T301 = T16[6'h21:6'h21];
  assign T302 = T16[6'h22:6'h22];
  assign T303 = T16[6'h23:6'h23];
  assign T304 = T16[6'h24:6'h24];
  assign T305 = T16[6'h25:6'h25];
  assign T306 = T16[6'h26:6'h26];
  assign T307 = T16[6'h27:6'h27];
  assign T308 = T16[6'h28:6'h28];
  assign T309 = T16[6'h29:6'h29];
  assign T310 = T16[6'h2a:6'h2a];
  assign T311 = T16[6'h2b:6'h2b];
  assign T312 = T16[6'h2c:6'h2c];
  assign T313 = T16[6'h2d:6'h2d];
  assign T314 = T16[6'h2e:6'h2e];
  assign T315 = T16[6'h2f:6'h2f];
  assign T316 = T16[6'h30:6'h30];
  assign T317 = T16[6'h31:6'h31];
  assign T318 = T16[6'h32:6'h32];
  assign T319 = T16[6'h33:6'h33];
  assign T320 = T16[6'h34:6'h34];
  assign T321 = T16[6'h35:6'h35];
  assign T322 = T16[6'h36:6'h36];
  assign T323 = T16[6'h37:6'h37];
  assign T324 = T16[6'h38:6'h38];
  assign T325 = T16[6'h39:6'h39];
  assign T326 = T16[6'h3a:6'h3a];
  assign T327 = T16[6'h3b:6'h3b];
  assign T328 = T16[6'h3c:6'h3c];
  assign T329 = T16[6'h3d:6'h3d];
  assign T330 = T16[6'h3e:6'h3e];
  assign T331 = T16[6'h3f:6'h3f];
  assign T17 = T33 ? T19 : T332;
  assign T332 = {32'h0, T18};
  assign T18 = T19[5'h1f:1'h0];
  assign T19 = T24 ? T23 : T20;
  assign T20 = R21[6'h3f:1'h0];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = 64'h0 - T20;
  assign T24 = T32 ? T31 : T25;
  assign T25 = T27 ? T26 : 1'h0;
  assign T26 = T20[6'h3f:6'h3f];
  assign T27 = T28 == 2'h3;
  assign T28 = R29 ^ 2'h1;
  assign T30 = io_in_valid ? io_in_bits_typ : R29;
  assign T31 = T20[5'h1f:5'h1f];
  assign T32 = T28 == 2'h1;
  assign T33 = T35 | T34;
  assign T34 = T28 == 2'h2;
  assign T35 = T28 == 2'h3;
  assign T36 = T13[6'h28:6'h27];
  assign T37 = T40 & R38;
  assign T39 = io_in_valid ? io_in_bits_single : R38;
  assign T40 = T41 == 5'h0;
  assign T41 = R42 & 5'h4;
  assign T43 = io_in_valid ? io_in_bits_cmd : R42;
  assign T44 = {3'h0, T45};
  assign T45 = {1'h0, T46};
  assign T46 = T47 != 2'h0;
  assign T47 = T48[1'h1:1'h0];
  assign T48 = {T70, T49};
  assign T49 = T50 != 10'h0;
  assign T50 = T51[4'h9:1'h0];
  assign T51 = T55 << T52;
  assign T52 = ~ T333;
  assign T333 = T457 ? 6'h3f : T334;
  assign T334 = T456 ? 6'h3e : T335;
  assign T335 = T455 ? 6'h3d : T336;
  assign T336 = T454 ? 6'h3c : T337;
  assign T337 = T453 ? 6'h3b : T338;
  assign T338 = T452 ? 6'h3a : T339;
  assign T339 = T451 ? 6'h39 : T340;
  assign T340 = T450 ? 6'h38 : T341;
  assign T341 = T449 ? 6'h37 : T342;
  assign T342 = T448 ? 6'h36 : T343;
  assign T343 = T447 ? 6'h35 : T344;
  assign T344 = T446 ? 6'h34 : T345;
  assign T345 = T445 ? 6'h33 : T346;
  assign T346 = T444 ? 6'h32 : T347;
  assign T347 = T443 ? 6'h31 : T348;
  assign T348 = T442 ? 6'h30 : T349;
  assign T349 = T441 ? 6'h2f : T350;
  assign T350 = T440 ? 6'h2e : T351;
  assign T351 = T439 ? 6'h2d : T352;
  assign T352 = T438 ? 6'h2c : T353;
  assign T353 = T437 ? 6'h2b : T354;
  assign T354 = T436 ? 6'h2a : T355;
  assign T355 = T435 ? 6'h29 : T356;
  assign T356 = T434 ? 6'h28 : T357;
  assign T357 = T433 ? 6'h27 : T358;
  assign T358 = T432 ? 6'h26 : T359;
  assign T359 = T431 ? 6'h25 : T360;
  assign T360 = T430 ? 6'h24 : T361;
  assign T361 = T429 ? 6'h23 : T362;
  assign T362 = T428 ? 6'h22 : T363;
  assign T363 = T427 ? 6'h21 : T364;
  assign T364 = T426 ? 6'h20 : T365;
  assign T365 = T425 ? 5'h1f : T366;
  assign T366 = T424 ? 5'h1e : T367;
  assign T367 = T423 ? 5'h1d : T368;
  assign T368 = T422 ? 5'h1c : T369;
  assign T369 = T421 ? 5'h1b : T370;
  assign T370 = T420 ? 5'h1a : T371;
  assign T371 = T419 ? 5'h19 : T372;
  assign T372 = T418 ? 5'h18 : T373;
  assign T373 = T417 ? 5'h17 : T374;
  assign T374 = T416 ? 5'h16 : T375;
  assign T375 = T415 ? 5'h15 : T376;
  assign T376 = T414 ? 5'h14 : T377;
  assign T377 = T413 ? 5'h13 : T378;
  assign T378 = T412 ? 5'h12 : T379;
  assign T379 = T411 ? 5'h11 : T380;
  assign T380 = T410 ? 5'h10 : T381;
  assign T381 = T409 ? 4'hf : T382;
  assign T382 = T408 ? 4'he : T383;
  assign T383 = T407 ? 4'hd : T384;
  assign T384 = T406 ? 4'hc : T385;
  assign T385 = T405 ? 4'hb : T386;
  assign T386 = T404 ? 4'ha : T387;
  assign T387 = T403 ? 4'h9 : T388;
  assign T388 = T402 ? 4'h8 : T389;
  assign T389 = T401 ? 3'h7 : T390;
  assign T390 = T400 ? 3'h6 : T391;
  assign T391 = T399 ? 3'h5 : T392;
  assign T392 = T398 ? 3'h4 : T393;
  assign T393 = T397 ? 2'h3 : T394;
  assign T394 = T396 ? 2'h2 : T395;
  assign T395 = T54[1'h1:1'h1];
  assign T54 = T55[6'h3f:1'h0];
  assign T396 = T54[2'h2:2'h2];
  assign T397 = T54[2'h3:2'h3];
  assign T398 = T54[3'h4:3'h4];
  assign T399 = T54[3'h5:3'h5];
  assign T400 = T54[3'h6:3'h6];
  assign T401 = T54[3'h7:3'h7];
  assign T402 = T54[4'h8:4'h8];
  assign T403 = T54[4'h9:4'h9];
  assign T404 = T54[4'ha:4'ha];
  assign T405 = T54[4'hb:4'hb];
  assign T406 = T54[4'hc:4'hc];
  assign T407 = T54[4'hd:4'hd];
  assign T408 = T54[4'he:4'he];
  assign T409 = T54[4'hf:4'hf];
  assign T410 = T54[5'h10:5'h10];
  assign T411 = T54[5'h11:5'h11];
  assign T412 = T54[5'h12:5'h12];
  assign T413 = T54[5'h13:5'h13];
  assign T414 = T54[5'h14:5'h14];
  assign T415 = T54[5'h15:5'h15];
  assign T416 = T54[5'h16:5'h16];
  assign T417 = T54[5'h17:5'h17];
  assign T418 = T54[5'h18:5'h18];
  assign T419 = T54[5'h19:5'h19];
  assign T420 = T54[5'h1a:5'h1a];
  assign T421 = T54[5'h1b:5'h1b];
  assign T422 = T54[5'h1c:5'h1c];
  assign T423 = T54[5'h1d:5'h1d];
  assign T424 = T54[5'h1e:5'h1e];
  assign T425 = T54[5'h1f:5'h1f];
  assign T426 = T54[6'h20:6'h20];
  assign T427 = T54[6'h21:6'h21];
  assign T428 = T54[6'h22:6'h22];
  assign T429 = T54[6'h23:6'h23];
  assign T430 = T54[6'h24:6'h24];
  assign T431 = T54[6'h25:6'h25];
  assign T432 = T54[6'h26:6'h26];
  assign T433 = T54[6'h27:6'h27];
  assign T434 = T54[6'h28:6'h28];
  assign T435 = T54[6'h29:6'h29];
  assign T436 = T54[6'h2a:6'h2a];
  assign T437 = T54[6'h2b:6'h2b];
  assign T438 = T54[6'h2c:6'h2c];
  assign T439 = T54[6'h2d:6'h2d];
  assign T440 = T54[6'h2e:6'h2e];
  assign T441 = T54[6'h2f:6'h2f];
  assign T442 = T54[6'h30:6'h30];
  assign T443 = T54[6'h31:6'h31];
  assign T444 = T54[6'h32:6'h32];
  assign T445 = T54[6'h33:6'h33];
  assign T446 = T54[6'h34:6'h34];
  assign T447 = T54[6'h35:6'h35];
  assign T448 = T54[6'h36:6'h36];
  assign T449 = T54[6'h37:6'h37];
  assign T450 = T54[6'h38:6'h38];
  assign T451 = T54[6'h39:6'h39];
  assign T452 = T54[6'h3a:6'h3a];
  assign T453 = T54[6'h3b:6'h3b];
  assign T454 = T54[6'h3c:6'h3c];
  assign T455 = T54[6'h3d:6'h3d];
  assign T456 = T54[6'h3e:6'h3e];
  assign T457 = T54[6'h3f:6'h3f];
  assign T55 = T67 ? T57 : T458;
  assign T458 = {32'h0, T56};
  assign T56 = T57[5'h1f:1'h0];
  assign T57 = T60 ? T59 : T58;
  assign T58 = R21[6'h3f:1'h0];
  assign T59 = 64'h0 - T58;
  assign T60 = T66 ? T65 : T61;
  assign T61 = T63 ? T62 : 1'h0;
  assign T62 = T58[6'h3f:6'h3f];
  assign T63 = T64 == 2'h3;
  assign T64 = R29 ^ 2'h1;
  assign T65 = T58[5'h1f:5'h1f];
  assign T66 = T64 == 2'h1;
  assign T67 = T69 | T68;
  assign T68 = T64 == 2'h2;
  assign T69 = T64 == 2'h3;
  assign T70 = T51[4'hb:4'ha];
  assign T71 = T40 & T72;
  assign T72 = R38 ^ 1'h1;
  assign T459 = reset ? 1'h0 : io_in_valid;
  assign T460 = reset ? 1'h0 : R73;
  assign io_out_bits_data = R75;
  assign T76 = R74 ? R77 : R75;
  assign T78 = R73 ? mux_data : R77;
  assign mux_data = T79;
  assign T79 = T71 ? T177 : T80;
  assign T80 = T37 ? T145 : T81;
  assign T81 = R38 ? T113 : T82;
  assign T82 = {T112, T83};
  assign T83 = {T94, T84};
  assign T84 = T92 ? T86 : T85;
  assign T85 = R21[6'h33:1'h0];
  assign T86 = T87[6'h3e:4'hb];
  assign T87 = T91 << T88;
  assign T88 = ~ T461;
  assign T461 = T585 ? 6'h3f : T462;
  assign T462 = T584 ? 6'h3e : T463;
  assign T463 = T583 ? 6'h3d : T464;
  assign T464 = T582 ? 6'h3c : T465;
  assign T465 = T581 ? 6'h3b : T466;
  assign T466 = T580 ? 6'h3a : T467;
  assign T467 = T579 ? 6'h39 : T468;
  assign T468 = T578 ? 6'h38 : T469;
  assign T469 = T577 ? 6'h37 : T470;
  assign T470 = T576 ? 6'h36 : T471;
  assign T471 = T575 ? 6'h35 : T472;
  assign T472 = T574 ? 6'h34 : T473;
  assign T473 = T573 ? 6'h33 : T474;
  assign T474 = T572 ? 6'h32 : T475;
  assign T475 = T571 ? 6'h31 : T476;
  assign T476 = T570 ? 6'h30 : T477;
  assign T477 = T569 ? 6'h2f : T478;
  assign T478 = T568 ? 6'h2e : T479;
  assign T479 = T567 ? 6'h2d : T480;
  assign T480 = T566 ? 6'h2c : T481;
  assign T481 = T565 ? 6'h2b : T482;
  assign T482 = T564 ? 6'h2a : T483;
  assign T483 = T563 ? 6'h29 : T484;
  assign T484 = T562 ? 6'h28 : T485;
  assign T485 = T561 ? 6'h27 : T486;
  assign T486 = T560 ? 6'h26 : T487;
  assign T487 = T559 ? 6'h25 : T488;
  assign T488 = T558 ? 6'h24 : T489;
  assign T489 = T557 ? 6'h23 : T490;
  assign T490 = T556 ? 6'h22 : T491;
  assign T491 = T555 ? 6'h21 : T492;
  assign T492 = T554 ? 6'h20 : T493;
  assign T493 = T553 ? 5'h1f : T494;
  assign T494 = T552 ? 5'h1e : T495;
  assign T495 = T551 ? 5'h1d : T496;
  assign T496 = T550 ? 5'h1c : T497;
  assign T497 = T549 ? 5'h1b : T498;
  assign T498 = T548 ? 5'h1a : T499;
  assign T499 = T547 ? 5'h19 : T500;
  assign T500 = T546 ? 5'h18 : T501;
  assign T501 = T545 ? 5'h17 : T502;
  assign T502 = T544 ? 5'h16 : T503;
  assign T503 = T543 ? 5'h15 : T504;
  assign T504 = T542 ? 5'h14 : T505;
  assign T505 = T541 ? 5'h13 : T506;
  assign T506 = T540 ? 5'h12 : T507;
  assign T507 = T539 ? 5'h11 : T508;
  assign T508 = T538 ? 5'h10 : T509;
  assign T509 = T537 ? 4'hf : T510;
  assign T510 = T536 ? 4'he : T511;
  assign T511 = T535 ? 4'hd : T512;
  assign T512 = T534 ? 4'hc : T513;
  assign T513 = T533 ? 4'hb : T514;
  assign T514 = T532 ? 4'ha : T515;
  assign T515 = T531 ? 4'h9 : T516;
  assign T516 = T530 ? 4'h8 : T517;
  assign T517 = T529 ? 3'h7 : T518;
  assign T518 = T528 ? 3'h6 : T519;
  assign T519 = T527 ? 3'h5 : T520;
  assign T520 = T526 ? 3'h4 : T521;
  assign T521 = T525 ? 2'h3 : T522;
  assign T522 = T524 ? 2'h2 : T523;
  assign T523 = T90[1'h1:1'h1];
  assign T90 = T91[6'h3f:1'h0];
  assign T524 = T90[2'h2:2'h2];
  assign T525 = T90[2'h3:2'h3];
  assign T526 = T90[3'h4:3'h4];
  assign T527 = T90[3'h5:3'h5];
  assign T528 = T90[3'h6:3'h6];
  assign T529 = T90[3'h7:3'h7];
  assign T530 = T90[4'h8:4'h8];
  assign T531 = T90[4'h9:4'h9];
  assign T532 = T90[4'ha:4'ha];
  assign T533 = T90[4'hb:4'hb];
  assign T534 = T90[4'hc:4'hc];
  assign T535 = T90[4'hd:4'hd];
  assign T536 = T90[4'he:4'he];
  assign T537 = T90[4'hf:4'hf];
  assign T538 = T90[5'h10:5'h10];
  assign T539 = T90[5'h11:5'h11];
  assign T540 = T90[5'h12:5'h12];
  assign T541 = T90[5'h13:5'h13];
  assign T542 = T90[5'h14:5'h14];
  assign T543 = T90[5'h15:5'h15];
  assign T544 = T90[5'h16:5'h16];
  assign T545 = T90[5'h17:5'h17];
  assign T546 = T90[5'h18:5'h18];
  assign T547 = T90[5'h19:5'h19];
  assign T548 = T90[5'h1a:5'h1a];
  assign T549 = T90[5'h1b:5'h1b];
  assign T550 = T90[5'h1c:5'h1c];
  assign T551 = T90[5'h1d:5'h1d];
  assign T552 = T90[5'h1e:5'h1e];
  assign T553 = T90[5'h1f:5'h1f];
  assign T554 = T90[6'h20:6'h20];
  assign T555 = T90[6'h21:6'h21];
  assign T556 = T90[6'h22:6'h22];
  assign T557 = T90[6'h23:6'h23];
  assign T558 = T90[6'h24:6'h24];
  assign T559 = T90[6'h25:6'h25];
  assign T560 = T90[6'h26:6'h26];
  assign T561 = T90[6'h27:6'h27];
  assign T562 = T90[6'h28:6'h28];
  assign T563 = T90[6'h29:6'h29];
  assign T564 = T90[6'h2a:6'h2a];
  assign T565 = T90[6'h2b:6'h2b];
  assign T566 = T90[6'h2c:6'h2c];
  assign T567 = T90[6'h2d:6'h2d];
  assign T568 = T90[6'h2e:6'h2e];
  assign T569 = T90[6'h2f:6'h2f];
  assign T570 = T90[6'h30:6'h30];
  assign T571 = T90[6'h31:6'h31];
  assign T572 = T90[6'h32:6'h32];
  assign T573 = T90[6'h33:6'h33];
  assign T574 = T90[6'h34:6'h34];
  assign T575 = T90[6'h35:6'h35];
  assign T576 = T90[6'h36:6'h36];
  assign T577 = T90[6'h37:6'h37];
  assign T578 = T90[6'h38:6'h38];
  assign T579 = T90[6'h39:6'h39];
  assign T580 = T90[6'h3a:6'h3a];
  assign T581 = T90[6'h3b:6'h3b];
  assign T582 = T90[6'h3c:6'h3c];
  assign T583 = T90[6'h3d:6'h3d];
  assign T584 = T90[6'h3e:6'h3e];
  assign T585 = T90[6'h3f:6'h3f];
  assign T91 = T85 << 4'hc;
  assign T92 = T93 == 11'h0;
  assign T93 = R21[6'h3e:6'h34];
  assign T94 = T101 | T586;
  assign T586 = {2'h0, T95};
  assign T95 = T96 << 4'h9;
  assign T96 = T99 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T85 == 52'h0;
  assign T99 = T100 == 2'h3;
  assign T100 = T101[4'hb:4'ha];
  assign T101 = T108 + T587;
  assign T587 = {1'h0, T102};
  assign T102 = T107 ? 11'h0 : T103;
  assign T103 = 11'h400 | T588;
  assign T588 = {9'h0, T104};
  assign T104 = T105 ? 2'h2 : 2'h1;
  assign T105 = T92 & T106;
  assign T106 = T98 ^ 1'h1;
  assign T107 = T92 & T98;
  assign T108 = T92 ? T109 : T589;
  assign T589 = {1'h0, T93};
  assign T109 = T98 ? 12'h0 : T110;
  assign T110 = {6'h3f, T111};
  assign T111 = ~ T88;
  assign T112 = R21[6'h3f:6'h3f];
  assign T113 = {32'hffffffff, T114};
  assign T114 = {T144, T115};
  assign T115 = {T126, T116};
  assign T116 = T124 ? T118 : T117;
  assign T117 = R21[5'h16:1'h0];
  assign T118 = T119[5'h1e:4'h8];
  assign T119 = T123 << T120;
  assign T120 = ~ T590;
  assign T590 = T650 ? 5'h1f : T591;
  assign T591 = T649 ? 5'h1e : T592;
  assign T592 = T648 ? 5'h1d : T593;
  assign T593 = T647 ? 5'h1c : T594;
  assign T594 = T646 ? 5'h1b : T595;
  assign T595 = T645 ? 5'h1a : T596;
  assign T596 = T644 ? 5'h19 : T597;
  assign T597 = T643 ? 5'h18 : T598;
  assign T598 = T642 ? 5'h17 : T599;
  assign T599 = T641 ? 5'h16 : T600;
  assign T600 = T640 ? 5'h15 : T601;
  assign T601 = T639 ? 5'h14 : T602;
  assign T602 = T638 ? 5'h13 : T603;
  assign T603 = T637 ? 5'h12 : T604;
  assign T604 = T636 ? 5'h11 : T605;
  assign T605 = T635 ? 5'h10 : T606;
  assign T606 = T634 ? 4'hf : T607;
  assign T607 = T633 ? 4'he : T608;
  assign T608 = T632 ? 4'hd : T609;
  assign T609 = T631 ? 4'hc : T610;
  assign T610 = T630 ? 4'hb : T611;
  assign T611 = T629 ? 4'ha : T612;
  assign T612 = T628 ? 4'h9 : T613;
  assign T613 = T627 ? 4'h8 : T614;
  assign T614 = T626 ? 3'h7 : T615;
  assign T615 = T625 ? 3'h6 : T616;
  assign T616 = T624 ? 3'h5 : T617;
  assign T617 = T623 ? 3'h4 : T618;
  assign T618 = T622 ? 2'h3 : T619;
  assign T619 = T621 ? 2'h2 : T620;
  assign T620 = T122[1'h1:1'h1];
  assign T122 = T123[5'h1f:1'h0];
  assign T621 = T122[2'h2:2'h2];
  assign T622 = T122[2'h3:2'h3];
  assign T623 = T122[3'h4:3'h4];
  assign T624 = T122[3'h5:3'h5];
  assign T625 = T122[3'h6:3'h6];
  assign T626 = T122[3'h7:3'h7];
  assign T627 = T122[4'h8:4'h8];
  assign T628 = T122[4'h9:4'h9];
  assign T629 = T122[4'ha:4'ha];
  assign T630 = T122[4'hb:4'hb];
  assign T631 = T122[4'hc:4'hc];
  assign T632 = T122[4'hd:4'hd];
  assign T633 = T122[4'he:4'he];
  assign T634 = T122[4'hf:4'hf];
  assign T635 = T122[5'h10:5'h10];
  assign T636 = T122[5'h11:5'h11];
  assign T637 = T122[5'h12:5'h12];
  assign T638 = T122[5'h13:5'h13];
  assign T639 = T122[5'h14:5'h14];
  assign T640 = T122[5'h15:5'h15];
  assign T641 = T122[5'h16:5'h16];
  assign T642 = T122[5'h17:5'h17];
  assign T643 = T122[5'h18:5'h18];
  assign T644 = T122[5'h19:5'h19];
  assign T645 = T122[5'h1a:5'h1a];
  assign T646 = T122[5'h1b:5'h1b];
  assign T647 = T122[5'h1c:5'h1c];
  assign T648 = T122[5'h1d:5'h1d];
  assign T649 = T122[5'h1e:5'h1e];
  assign T650 = T122[5'h1f:5'h1f];
  assign T123 = T117 << 4'h9;
  assign T124 = T125 == 8'h0;
  assign T125 = R21[5'h1e:5'h17];
  assign T126 = T133 | T651;
  assign T651 = {2'h0, T127};
  assign T127 = T128 << 3'h6;
  assign T128 = T131 & T129;
  assign T129 = T130 ^ 1'h1;
  assign T130 = T117 == 23'h0;
  assign T131 = T132 == 2'h3;
  assign T132 = T133[4'h8:3'h7];
  assign T133 = T140 + T652;
  assign T652 = {1'h0, T134};
  assign T134 = T139 ? 8'h0 : T135;
  assign T135 = 8'h80 | T653;
  assign T653 = {6'h0, T136};
  assign T136 = T137 ? 2'h2 : 2'h1;
  assign T137 = T124 & T138;
  assign T138 = T130 ^ 1'h1;
  assign T139 = T124 & T130;
  assign T140 = T124 ? T141 : T654;
  assign T654 = {1'h0, T125};
  assign T141 = T130 ? 9'h0 : T142;
  assign T142 = {4'hf, T143};
  assign T143 = ~ T120;
  assign T144 = R21[5'h1f:5'h1f];
  assign T145 = {32'hffffffff, T146};
  assign T146 = {T24, T147};
  assign T147 = {T169, T148};
  assign T148 = T149[5'h16:1'h0];
  assign T149 = T153 ? T152 : T150;
  assign T150 = {1'h0, T151};
  assign T151 = T13[6'h3f:6'h28];
  assign T152 = T150 + 25'h1;
  assign T153 = T168 ? T163 : T154;
  assign T154 = T162 ? T161 : T155;
  assign T155 = T158 ? T156 : 1'h0;
  assign T156 = T157 & T8;
  assign T157 = T24 ^ 1'h1;
  assign T158 = R159 == 3'h3;
  assign T160 = io_in_valid ? io_in_bits_rm : R159;
  assign T161 = T24 & T8;
  assign T162 = R159 == 3'h2;
  assign T163 = T166 | T164;
  assign T164 = T165 == 2'h3;
  assign T165 = T10[1'h1:1'h0];
  assign T166 = T167 == 2'h3;
  assign T167 = T10[2'h2:1'h1];
  assign T168 = R159 == 3'h0;
  assign T169 = {T176, T170};
  assign T170 = T171[3'h7:1'h0];
  assign T171 = T173 + T655;
  assign T655 = {7'h0, T172};
  assign T172 = T149[5'h18:5'h18];
  assign T173 = {1'h0, T174};
  assign T174 = {1'h0, T175};
  assign T175 = ~ T14;
  assign T176 = T13[6'h3f:6'h3f];
  assign T177 = {T60, T178};
  assign T178 = {T198, T179};
  assign T179 = T180[6'h33:1'h0];
  assign T180 = T184 ? T183 : T181;
  assign T181 = {1'h0, T182};
  assign T182 = T51[6'h3f:4'hb];
  assign T183 = T181 + 54'h1;
  assign T184 = T197 ? T192 : T185;
  assign T185 = T191 ? T190 : T186;
  assign T186 = T189 ? T187 : 1'h0;
  assign T187 = T188 & T46;
  assign T188 = T60 ^ 1'h1;
  assign T189 = R159 == 3'h3;
  assign T190 = T60 & T46;
  assign T191 = R159 == 3'h2;
  assign T192 = T195 | T193;
  assign T193 = T194 == 2'h3;
  assign T194 = T48[1'h1:1'h0];
  assign T195 = T196 == 2'h3;
  assign T196 = T48[2'h2:1'h1];
  assign T197 = R159 == 3'h0;
  assign T198 = {T205, T199};
  assign T199 = T200[4'ha:1'h0];
  assign T200 = T202 + T656;
  assign T656 = {10'h0, T201};
  assign T201 = T180[6'h35:6'h35];
  assign T202 = {1'h0, T203};
  assign T203 = {4'h0, T204};
  assign T204 = ~ T52;
  assign T205 = T51[6'h3f:6'h3f];
  assign io_out_valid = R206;
  assign T657 = reset ? 1'h0 : R74;

  always @(posedge clk) begin
    if(R74) begin
      R0 <= R2;
    end
    if(R73) begin
      R2 <= mux_exc;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R29 <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      R38 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R42 <= io_in_bits_cmd;
    end
    if(reset) begin
      R73 <= 1'h0;
    end else begin
      R73 <= io_in_valid;
    end
    if(reset) begin
      R74 <= 1'h0;
    end else begin
      R74 <= R73;
    end
    if(R74) begin
      R75 <= R77;
    end
    if(R73) begin
      R77 <= mux_data;
    end
    if(io_in_valid) begin
      R159 <= io_in_bits_rm;
    end
    if(reset) begin
      R206 <= 1'h0;
    end else begin
      R206 <= R74;
    end
  end
endmodule

module FPToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc,
    input  io_lt
);

  reg [4:0] R0;
  wire[4:0] T1;
  wire[4:0] mux_exc;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] minmax_exc;
  wire T5;
  wire issnan2;
  wire T6;
  wire T7;
  wire T8;
  reg [64:0] R9;
  wire[64:0] T10;
  wire T11;
  reg  R12;
  wire T13;
  wire isnan2;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire issnan1;
  wire T18;
  wire T19;
  wire T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire T23;
  wire isnan1;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire isSgnj;
  wire[4:0] T28;
  reg [4:0] R29;
  wire[4:0] T30;
  wire[4:0] T31;
  wire[2:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[2:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire[11:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[1:0] T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire[27:0] T56;
  wire[51:0] T57;
  wire T58;
  wire[23:0] T59;
  wire[48:0] T60;
  wire[4:0] T61;
  wire[11:0] T62;
  wire[11:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire[48:0] T67;
  wire[47:0] T68;
  wire[23:0] T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[24:0] T76;
  wire[24:0] T77;
  wire[24:0] T78;
  wire[24:0] T79;
  wire[55:0] T80;
  wire[4:0] T81;
  wire[24:0] T82;
  wire[22:0] T83;
  wire[24:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  reg [2:0] R92;
  wire[2:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[1:0] T98;
  wire T99;
  wire[1:0] T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire[4:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[22:0] T115;
  wire T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  reg  R120;
  wire T200;
  reg [64:0] R121;
  wire[64:0] T122;
  wire[64:0] mux_data;
  wire[64:0] T123;
  wire[64:0] T124;
  wire[64:0] T125;
  wire[64:0] fsgnj;
  wire[32:0] T126;
  wire[31:0] T127;
  wire sign_s;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire sign_d;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire isLHS;
  wire T150;
  wire T151;
  wire T152;
  wire isMax;
  wire[64:0] T153;
  wire[32:0] T154;
  wire[31:0] T155;
  wire[22:0] T156;
  wire[22:0] T157;
  wire[22:0] T158;
  wire[22:0] T159;
  wire[22:0] T160;
  wire[22:0] T201;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[22:0] T170;
  wire[22:0] T202;
  wire[8:0] T171;
  wire[8:0] T172;
  wire[8:0] T173;
  wire[8:0] T174;
  wire[8:0] T175;
  wire[8:0] T176;
  wire[8:0] T177;
  wire T178;
  wire[8:0] T203;
  wire[6:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire[64:0] T182;
  wire[63:0] T183;
  wire[51:0] T184;
  wire[51:0] T185;
  wire[51:0] T186;
  wire[51:0] T204;
  wire[11:0] T187;
  wire[11:0] T188;
  wire[11:0] T189;
  wire[11:0] T190;
  wire T191;
  wire[11:0] T192;
  wire[7:0] T196;
  wire T193;
  wire[11:0] T205;
  wire[10:0] T194;
  wire T195;
  wire[11:0] T206;
  wire T197;
  wire T198;
  reg  R199;
  wire T207;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R9 = {3{$random}};
    R12 = {1{$random}};
    R21 = {3{$random}};
    R29 = {1{$random}};
    R92 = {1{$random}};
    R120 = {1{$random}};
    R121 = {3{$random}};
    R199 = {1{$random}};
  end
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R120 ? mux_exc : R0;
  assign mux_exc = T2;
  assign T2 = T118 ? T111 : T3;
  assign T3 = T108 ? T31 : T4;
  assign T4 = isSgnj ? 5'h0 : minmax_exc;
  assign minmax_exc = {T5, 4'h0};
  assign T5 = issnan1 | issnan2;
  assign issnan2 = isnan2 & T6;
  assign T6 = ~ T7;
  assign T7 = R12 ? T11 : T8;
  assign T8 = R9[6'h33:6'h33];
  assign T10 = io_in_valid ? io_in_bits_in2 : R9;
  assign T11 = R9[5'h16:5'h16];
  assign T13 = io_in_valid ? io_in_bits_single : R12;
  assign isnan2 = R12 ? T16 : T14;
  assign T14 = T15 == 3'h7;
  assign T15 = R9[6'h3f:6'h3d];
  assign T16 = T17 == 3'h7;
  assign T17 = R9[5'h1f:5'h1d];
  assign issnan1 = isnan1 & T18;
  assign T18 = ~ T19;
  assign T19 = R12 ? T23 : T20;
  assign T20 = R21[6'h33:6'h33];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = R21[5'h16:5'h16];
  assign isnan1 = R12 ? T26 : T24;
  assign T24 = T25 == 3'h7;
  assign T25 = R21[6'h3f:6'h3d];
  assign T26 = T27 == 3'h7;
  assign T27 = R21[5'h1f:5'h1d];
  assign isSgnj = T28 == 5'h4;
  assign T28 = R29 & 5'h5;
  assign T30 = io_in_valid ? io_in_bits_cmd : R29;
  assign T31 = {T103, T32};
  assign T32 = {T73, T33};
  assign T33 = {T71, T34};
  assign T34 = T45 | T35;
  assign T35 = T43 & T36;
  assign T36 = T37 ^ 1'h1;
  assign T37 = T41 | T38;
  assign T38 = T39 == 2'h3;
  assign T39 = T40[2'h2:1'h1];
  assign T40 = R21[6'h3f:6'h3d];
  assign T41 = T42 ^ 1'h1;
  assign T42 = T40 != 3'h0;
  assign T43 = T44 < 12'h76a;
  assign T44 = R21[6'h3f:6'h34];
  assign T45 = T49 | T46;
  assign T46 = T48 & T47;
  assign T47 = T37 ^ 1'h1;
  assign T48 = 12'h87f < T44;
  assign T49 = T51 & T50;
  assign T50 = T37 ^ 1'h1;
  assign T51 = T52 != 2'h0;
  assign T52 = T53[1'h1:1'h0];
  assign T53 = {T70, T54};
  assign T54 = T58 | T55;
  assign T55 = T56 != 28'h0;
  assign T56 = T57[5'h1b:1'h0];
  assign T57 = R21[6'h33:1'h0];
  assign T58 = T59 != 24'h0;
  assign T59 = T60[5'h17:1'h0];
  assign T60 = T67 >> T61;
  assign T61 = T62[3'h4:1'h0];
  assign T62 = T64 ? T63 : 12'h0;
  assign T63 = 12'h782 - T44;
  assign T64 = T66 & T65;
  assign T65 = T44 <= 12'h781;
  assign T66 = 12'h76a <= T44;
  assign T67 = {1'h1, T68};
  assign T68 = {T69, 24'h0};
  assign T69 = T57[6'h33:5'h1c];
  assign T70 = T60[5'h19:5'h18];
  assign T71 = T35 | T72;
  assign T72 = T64 & T49;
  assign T73 = T46 | T74;
  assign T74 = T102 & T75;
  assign T75 = T76[5'h18:5'h18];
  assign T76 = T85 ? T84 : T77;
  assign T77 = T82 | T78;
  assign T78 = ~ T79;
  assign T79 = T80[5'h18:1'h0];
  assign T80 = 25'h1ffffff << T81;
  assign T81 = T61;
  assign T82 = {2'h1, T83};
  assign T83 = T57[6'h33:5'h1d];
  assign T84 = T77 + 25'h1;
  assign T85 = T101 ? T96 : T86;
  assign T86 = T95 ? T94 : T87;
  assign T87 = T91 ? T88 : 1'h0;
  assign T88 = T89 & T49;
  assign T89 = T90 ^ 1'h1;
  assign T90 = R21[7'h40:7'h40];
  assign T91 = R92 == 3'h3;
  assign T93 = io_in_valid ? io_in_bits_rm : R92;
  assign T94 = T90 & T49;
  assign T95 = R92 == 3'h2;
  assign T96 = T99 | T97;
  assign T97 = T98 == 2'h3;
  assign T98 = T53[2'h2:1'h1];
  assign T99 = T100 == 2'h3;
  assign T100 = T53[1'h1:1'h0];
  assign T101 = R92 == 3'h0;
  assign T102 = T44 == 12'h87f;
  assign T103 = {T104, 1'h0};
  assign T104 = T107 & T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = T57[6'h33:6'h33];
  assign T107 = T40 == 3'h7;
  assign T108 = T109 & R12;
  assign T109 = T110 == 5'h0;
  assign T110 = R29 & 5'h4;
  assign T111 = T112 << 3'h4;
  assign T112 = T116 & T113;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115[5'h16:5'h16];
  assign T115 = R21[5'h16:1'h0];
  assign T116 = T117 == 3'h7;
  assign T117 = R21[5'h1f:5'h1d];
  assign T118 = T109 & T119;
  assign T119 = R12 ^ 1'h1;
  assign T200 = reset ? 1'h0 : io_in_valid;
  assign io_out_bits_data = R121;
  assign T122 = R120 ? mux_data : R121;
  assign mux_data = T123;
  assign T123 = T118 ? T182 : T124;
  assign T124 = T108 ? T153 : T125;
  assign T125 = T149 ? fsgnj : R9;
  assign fsgnj = {T137, T126};
  assign T126 = {sign_s, T127};
  assign T127 = R21[5'h1f:1'h0];
  assign sign_s = T131 ^ T128;
  assign T128 = T130 & T129;
  assign T129 = R9[6'h20:6'h20];
  assign T130 = R12 & isSgnj;
  assign T131 = T134 ? T133 : T132;
  assign T132 = R92[1'h0:1'h0];
  assign T133 = R21[6'h20:6'h20];
  assign T134 = T136 | T135;
  assign T135 = T130 ^ 1'h1;
  assign T136 = R92[1'h1:1'h1];
  assign T137 = {sign_d, T138};
  assign T138 = R21[6'h3f:6'h21];
  assign sign_d = T143 ^ T139;
  assign T139 = T141 & T140;
  assign T140 = R9[7'h40:7'h40];
  assign T141 = T142 & isSgnj;
  assign T142 = R12 ^ 1'h1;
  assign T143 = T146 ? T145 : T144;
  assign T144 = R92[1'h0:1'h0];
  assign T145 = R21[7'h40:7'h40];
  assign T146 = T148 | T147;
  assign T147 = T141 ^ 1'h1;
  assign T148 = R92[1'h1:1'h1];
  assign T149 = isSgnj | isLHS;
  assign isLHS = isnan2 | T150;
  assign T150 = T152 & T151;
  assign T151 = isnan1 ^ 1'h1;
  assign T152 = isMax != io_lt;
  assign isMax = R92[1'h0:1'h0];
  assign T153 = {32'hffffffff, T154};
  assign T154 = {T90, T155};
  assign T155 = {T171, T156};
  assign T156 = T37 ? T170 : T157;
  assign T157 = T46 ? T160 : T158;
  assign T158 = T35 ? 23'h0 : T159;
  assign T159 = T76[5'h16:1'h0];
  assign T160 = 23'h0 - T201;
  assign T201 = {22'h0, T161};
  assign T161 = T162 ^ 1'h1;
  assign T162 = T164 | T163;
  assign T163 = R92 == 3'h0;
  assign T164 = T168 | T165;
  assign T165 = T167 & T166;
  assign T166 = T90 ^ 1'h1;
  assign T167 = R92 == 3'h3;
  assign T168 = T169 & T90;
  assign T169 = R92 == 3'h2;
  assign T170 = 23'h0 - T202;
  assign T202 = {22'h0, T107};
  assign T171 = T37 ? T181 : T172;
  assign T172 = T46 ? T180 : T173;
  assign T173 = T35 ? T203 : T174;
  assign T174 = T178 ? T177 : T175;
  assign T175 = T176 + 9'h100;
  assign T176 = T44[4'h8:1'h0];
  assign T177 = T175 + 9'h1;
  assign T178 = T76[5'h18:5'h18];
  assign T203 = {2'h0, T179};
  assign T179 = T164 ? 7'h6b : 7'h0;
  assign T180 = T162 ? 9'h180 : 9'h17f;
  assign T181 = T40 << 3'h6;
  assign T182 = {T198, T183};
  assign T183 = {T187, T184};
  assign T184 = T186 | T185;
  assign T185 = T115 << 5'h1d;
  assign T186 = 52'h0 - T204;
  assign T204 = {51'h0, T116};
  assign T187 = T197 ? T206 : T188;
  assign T188 = T195 ? T205 : T189;
  assign T189 = T193 ? T192 : T190;
  assign T190 = T191 ? 12'hc00 : 12'he00;
  assign T191 = T117 < 3'h7;
  assign T192 = {4'h8, T196};
  assign T196 = R21[5'h1e:5'h17];
  assign T193 = T117 < 3'h6;
  assign T205 = {1'h0, T194};
  assign T194 = {3'h7, T196};
  assign T195 = T117 < 3'h4;
  assign T206 = {4'h0, T196};
  assign T197 = T117 < 3'h1;
  assign T198 = R21[6'h20:6'h20];
  assign io_out_valid = R199;
  assign T207 = reset ? 1'h0 : R120;

  always @(posedge clk) begin
    if(R120) begin
      R0 <= mux_exc;
    end
    if(io_in_valid) begin
      R9 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      R12 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R29 <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      R92 <= io_in_bits_rm;
    end
    if(reset) begin
      R120 <= 1'h0;
    end else begin
      R120 <= io_in_valid;
    end
    if(R120) begin
      R121 <= mux_data;
    end
    if(reset) begin
      R199 <= 1'h0;
    end else begin
      R199 <= R120;
    end
  end
endmodule

module FPU(input clk, input reset,
    input  io_ctrl_valid,
    output io_ctrl_fcsr_rdy,
    output io_ctrl_nack_mem,
    output io_ctrl_illegal_rm,
    input  io_ctrl_killx,
    input  io_ctrl_killm,
    output[4:0] io_ctrl_dec_cmd,
    output io_ctrl_dec_ldst,
    output io_ctrl_dec_wen,
    output io_ctrl_dec_ren1,
    output io_ctrl_dec_ren2,
    output io_ctrl_dec_ren3,
    output io_ctrl_dec_swap23,
    output io_ctrl_dec_single,
    output io_ctrl_dec_fromint,
    output io_ctrl_dec_toint,
    output io_ctrl_dec_fastpipe,
    output io_ctrl_dec_fma,
    output io_ctrl_dec_round,
    output io_ctrl_sboard_set,
    output io_ctrl_sboard_clr,
    output[4:0] io_ctrl_sboard_clra,
    input [31:0] io_dpath_inst,
    input [63:0] io_dpath_fromint_data,
    input [2:0] io_dpath_fcsr_rm,
    output io_dpath_fcsr_flags_valid,
    output[4:0] io_dpath_fcsr_flags_bits,
    output[63:0] io_dpath_store_data,
    output[63:0] io_dpath_toint_data,
    input  io_dpath_dmem_resp_val,
    input [2:0] io_dpath_dmem_resp_type,
    input [4:0] io_dpath_dmem_resp_tag,
    input [63:0] io_dpath_dmem_resp_data
);

  wire[64:0] req_in3;
  wire[64:0] ex_rs3;
  reg [64:0] regfile [31:0];
  wire[64:0] T120;
  wire[64:0] T121;
  wire[96:0] wdata;
  wire[96:0] T122;
  wire[64:0] T123;
  wire T124;
  wire[1:0] T125;
  wire[1:0] wsrc;
  reg [6:0] winfo_0;
  wire[6:0] T5;
  wire[6:0] T6;
  reg [6:0] winfo_1;
  wire[6:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] memLatencyMask;
  wire[1:0] T11;
  wire T12;
  wire T13;
  reg  mem_ctrl_single;
  wire T14;
  reg  ex_ctrl_single;
  wire T15;
  reg  ex_reg_valid;
  wire T105;
  reg  mem_ctrl_fma;
  wire T16;
  reg  ex_ctrl_fma;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T106;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  reg  mem_ctrl_fromint;
  wire T22;
  reg  ex_ctrl_fromint;
  wire T23;
  wire[1:0] T107;
  reg  mem_ctrl_fastpipe;
  wire T24;
  reg  ex_ctrl_fastpipe;
  wire T25;
  wire T26;
  reg  write_port_busy;
  wire T27;
  wire T28;
  wire T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire[3:0] T35;
  wire[3:0] T108;
  wire[2:0] T36;
  wire T37;
  wire[3:0] T38;
  wire[3:0] T39;
  wire[3:0] T109;
  wire[2:0] T40;
  wire[3:0] T110;
  reg [1:0] wen;
  wire[1:0] T111;
  wire[1:0] T41;
  wire[1:0] T112;
  wire T42;
  wire[1:0] T43;
  wire[1:0] T113;
  wire T44;
  wire T45;
  wire T46;
  wire killm;
  wire T47;
  wire T48;
  wire[2:0] T49;
  wire[2:0] T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T114;
  wire[1:0] T55;
  wire T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T115;
  wire[1:0] T59;
  wire[2:0] T116;
  wire mem_wen;
  wire T60;
  wire T61;
  reg  mem_reg_valid;
  wire T117;
  wire T62;
  wire T63;
  wire T64;
  wire[6:0] mem_winfo;
  wire[4:0] T65;
  reg [31:0] mem_reg_inst;
  wire[31:0] T66;
  reg [31:0] ex_reg_inst;
  wire[31:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T118;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[96:0] T126;
  wire[96:0] T127;
  wire[96:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[4:0] T132;
  wire[4:0] waddr;
  wire[4:0] T93;
  wire[64:0] T133;
  wire[64:0] load_wb_data_recoded;
  wire[64:0] rec_d;
  wire[63:0] T134;
  wire[51:0] T135;
  wire[51:0] T136;
  reg [63:0] load_wb_data;
  wire[63:0] T137;
  wire[51:0] T138;
  wire[126:0] T139;
  wire[5:0] T140;
  wire[5:0] T141;
  wire[5:0] T142;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire[5:0] T146;
  wire[5:0] T147;
  wire[5:0] T148;
  wire[5:0] T149;
  wire[5:0] T150;
  wire[5:0] T151;
  wire[5:0] T152;
  wire[5:0] T153;
  wire[5:0] T154;
  wire[5:0] T155;
  wire[5:0] T156;
  wire[5:0] T157;
  wire[5:0] T158;
  wire[5:0] T159;
  wire[5:0] T160;
  wire[5:0] T161;
  wire[5:0] T162;
  wire[5:0] T163;
  wire[5:0] T164;
  wire[5:0] T165;
  wire[5:0] T166;
  wire[5:0] T167;
  wire[5:0] T168;
  wire[5:0] T169;
  wire[5:0] T170;
  wire[5:0] T171;
  wire[5:0] T172;
  wire[4:0] T173;
  wire[4:0] T174;
  wire[4:0] T175;
  wire[4:0] T176;
  wire[4:0] T177;
  wire[4:0] T178;
  wire[4:0] T179;
  wire[4:0] T180;
  wire[4:0] T181;
  wire[4:0] T182;
  wire[4:0] T183;
  wire[4:0] T184;
  wire[4:0] T185;
  wire[4:0] T186;
  wire[4:0] T187;
  wire[4:0] T188;
  wire[3:0] T189;
  wire[3:0] T190;
  wire[3:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[3:0] T195;
  wire[3:0] T196;
  wire[2:0] T197;
  wire[2:0] T198;
  wire[2:0] T199;
  wire[2:0] T200;
  wire[1:0] T201;
  wire[1:0] T202;
  wire T203;
  wire[63:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire[63:0] T267;
  wire T268;
  wire[10:0] T269;
  wire[11:0] T270;
  wire[11:0] T271;
  wire[9:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire[1:0] T277;
  wire[11:0] T278;
  wire[11:0] T279;
  wire[10:0] T280;
  wire[10:0] T281;
  wire[10:0] T282;
  wire[1:0] T283;
  wire T284;
  wire T285;
  wire T286;
  wire[11:0] T287;
  wire[11:0] T288;
  wire[11:0] T289;
  wire[11:0] T290;
  wire[5:0] T291;
  wire T292;
  wire[64:0] T293;
  wire[32:0] rec_s;
  wire[31:0] T294;
  wire[22:0] T295;
  wire[22:0] T296;
  wire[22:0] T297;
  wire[62:0] T298;
  wire[4:0] T299;
  wire[4:0] T300;
  wire[4:0] T301;
  wire[4:0] T302;
  wire[4:0] T303;
  wire[4:0] T304;
  wire[4:0] T305;
  wire[4:0] T306;
  wire[4:0] T307;
  wire[4:0] T308;
  wire[4:0] T309;
  wire[4:0] T310;
  wire[4:0] T311;
  wire[4:0] T312;
  wire[4:0] T313;
  wire[4:0] T314;
  wire[4:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[3:0] T318;
  wire[3:0] T319;
  wire[3:0] T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[2:0] T324;
  wire[2:0] T325;
  wire[2:0] T326;
  wire[2:0] T327;
  wire[1:0] T328;
  wire[1:0] T329;
  wire T330;
  wire[31:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire[31:0] T362;
  wire T363;
  wire[7:0] T364;
  wire[8:0] T365;
  wire[8:0] T366;
  wire[6:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[1:0] T372;
  wire[8:0] T373;
  wire[8:0] T374;
  wire[7:0] T375;
  wire[7:0] T376;
  wire[7:0] T377;
  wire[1:0] T378;
  wire T379;
  wire T380;
  wire T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire[8:0] T384;
  wire[8:0] T385;
  wire[4:0] T386;
  wire T387;
  reg  load_wb_single;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  reg  load_wb;
  reg [4:0] load_wb_tag;
  wire[4:0] T392;
  reg [4:0] ex_ra3;
  wire[4:0] T393;
  wire[4:0] T394;
  wire[4:0] T395;
  wire T396;
  wire[4:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire[64:0] req_in2;
  wire[64:0] ex_rs2;
  reg [4:0] ex_ra2;
  wire[4:0] T402;
  wire[4:0] T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[64:0] req_in1;
  wire[64:0] ex_rs1;
  reg [4:0] ex_ra1;
  wire[4:0] T408;
  wire[4:0] T409;
  wire[4:0] T410;
  wire T411;
  wire[4:0] T412;
  wire T413;
  wire[1:0] req_typ;
  wire[1:0] T414;
  wire[2:0] req_rm;
  wire[2:0] ex_rm;
  wire[2:0] T99;
  wire T100;
  wire[2:0] T101;
  wire req_round;
  reg  ex_ctrl_round;
  wire T97;
  wire req_fma;
  wire req_fastpipe;
  wire req_toint;
  reg  ex_ctrl_toint;
  wire T87;
  wire req_fromint;
  wire req_single;
  wire req_swap23;
  reg  ex_ctrl_swap23;
  wire T415;
  wire req_ren3;
  reg  ex_ctrl_ren3;
  wire T416;
  wire req_ren2;
  reg  ex_ctrl_ren2;
  wire T417;
  wire req_ren1;
  reg  ex_ctrl_ren1;
  wire T418;
  wire req_wen;
  reg  ex_ctrl_wen;
  wire T419;
  wire req_ldst;
  reg  ex_ctrl_ldst;
  wire T420;
  wire[4:0] req_cmd;
  reg [4:0] ex_ctrl_cmd;
  wire[4:0] T421;
  wire T422;
  wire[64:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[4:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] wexc;
  wire[4:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[4:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire[4:0] T84;
  reg [4:0] wb_toint_exc;
  wire[4:0] T85;
  reg  mem_ctrl_toint;
  wire T86;
  wire wb_toint_valid;
  reg  wb_ctrl_toint;
  wire T88;
  reg  wb_reg_valid;
  wire T119;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T94;
  reg  R95;
  wire T96;
  wire T98;
  wire T102;
  wire fp_inflight;
  wire T103;
  wire T104;
  wire[4:0] fp_decoder_io_sigs_cmd;
  wire fp_decoder_io_sigs_ldst;
  wire fp_decoder_io_sigs_wen;
  wire fp_decoder_io_sigs_ren1;
  wire fp_decoder_io_sigs_ren2;
  wire fp_decoder_io_sigs_ren3;
  wire fp_decoder_io_sigs_swap23;
  wire fp_decoder_io_sigs_single;
  wire fp_decoder_io_sigs_fromint;
  wire fp_decoder_io_sigs_toint;
  wire fp_decoder_io_sigs_fastpipe;
  wire fp_decoder_io_sigs_fma;
  wire fp_decoder_io_sigs_round;
  wire[64:0] ifpu_io_out_bits_data;
  wire[4:0] ifpu_io_out_bits_exc;
  wire[64:0] fpmu_io_out_bits_data;
  wire[4:0] fpmu_io_out_bits_exc;
  wire[64:0] sfma_io_out_bits_data;
  wire[4:0] sfma_io_out_bits_exc;
  wire[64:0] dfma_io_out_bits_data;
  wire[4:0] dfma_io_out_bits_exc;
  wire fpiu_io_out_bits_lt;
  wire[63:0] fpiu_io_out_bits_store;
  wire[63:0] fpiu_io_out_bits_toint;
  wire[4:0] fpiu_io_out_bits_exc;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 32; initvar = initvar+1)
      regfile[initvar] = {3{$random}};
    winfo_0 = {1{$random}};
    winfo_1 = {1{$random}};
    mem_ctrl_single = {1{$random}};
    ex_ctrl_single = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_ctrl_fma = {1{$random}};
    ex_ctrl_fma = {1{$random}};
    mem_ctrl_fromint = {1{$random}};
    ex_ctrl_fromint = {1{$random}};
    mem_ctrl_fastpipe = {1{$random}};
    ex_ctrl_fastpipe = {1{$random}};
    write_port_busy = {1{$random}};
    wen = {1{$random}};
    mem_reg_valid = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    load_wb_data = {2{$random}};
    load_wb_single = {1{$random}};
    load_wb = {1{$random}};
    load_wb_tag = {1{$random}};
    ex_ra3 = {1{$random}};
    ex_ra2 = {1{$random}};
    ex_ra1 = {1{$random}};
    ex_ctrl_round = {1{$random}};
    ex_ctrl_toint = {1{$random}};
    ex_ctrl_swap23 = {1{$random}};
    ex_ctrl_ren3 = {1{$random}};
    ex_ctrl_ren2 = {1{$random}};
    ex_ctrl_ren1 = {1{$random}};
    ex_ctrl_wen = {1{$random}};
    ex_ctrl_ldst = {1{$random}};
    ex_ctrl_cmd = {1{$random}};
    wb_toint_exc = {1{$random}};
    mem_ctrl_toint = {1{$random}};
    wb_ctrl_toint = {1{$random}};
    wb_reg_valid = {1{$random}};
    R95 = {1{$random}};
  end
`endif

  assign req_in3 = ex_rs3;
  assign ex_rs3 = regfile[ex_ra3];
  assign T121 = wdata[7'h40:1'h0];
  assign wdata = T130 ? T126 : T122;
  assign T122 = {32'h0, T123};
  assign T123 = T124 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data;
  assign T124 = T125[1'h0:1'h0];
  assign T125 = wsrc;
  assign wsrc = winfo_0 >> 3'h5;
  assign T5 = T76 ? mem_winfo : T6;
  assign T6 = T64 ? winfo_1 : winfo_0;
  assign T7 = T8 ? mem_winfo : winfo_1;
  assign T8 = mem_wen & T9;
  assign T9 = T26 & T10;
  assign T10 = memLatencyMask[1'h1:1'h1];
  assign memLatencyMask = T18 | T11;
  assign T11 = T12 ? 2'h2 : 2'h0;
  assign T12 = mem_ctrl_fma & T13;
  assign T13 = mem_ctrl_single ^ 1'h1;
  assign T14 = ex_reg_valid ? ex_ctrl_single : mem_ctrl_single;
  assign T15 = io_ctrl_valid ? fp_decoder_io_sigs_single : ex_ctrl_single;
  assign T105 = reset ? 1'h0 : io_ctrl_valid;
  assign T16 = ex_reg_valid ? ex_ctrl_fma : mem_ctrl_fma;
  assign T17 = io_ctrl_valid ? fp_decoder_io_sigs_fma : ex_ctrl_fma;
  assign T18 = T20 | T106;
  assign T106 = {1'h0, T19};
  assign T19 = mem_ctrl_fma & mem_ctrl_single;
  assign T20 = T107 | T21;
  assign T21 = mem_ctrl_fromint ? 2'h2 : 2'h0;
  assign T22 = ex_reg_valid ? ex_ctrl_fromint : mem_ctrl_fromint;
  assign T23 = io_ctrl_valid ? fp_decoder_io_sigs_fromint : ex_ctrl_fromint;
  assign T107 = {1'h0, mem_ctrl_fastpipe};
  assign T24 = ex_reg_valid ? ex_ctrl_fastpipe : mem_ctrl_fastpipe;
  assign T25 = io_ctrl_valid ? fp_decoder_io_sigs_fastpipe : ex_ctrl_fastpipe;
  assign T26 = write_port_busy ^ 1'h1;
  assign T27 = ex_reg_valid ? T28 : write_port_busy;
  assign T28 = T47 | T29;
  assign T29 = T30 != 4'h0;
  assign T30 = T110 & T31;
  assign T31 = T35 | T32;
  assign T32 = T33 ? 4'h8 : 4'h0;
  assign T33 = ex_ctrl_fma & T34;
  assign T34 = ex_ctrl_single ^ 1'h1;
  assign T35 = T38 | T108;
  assign T108 = {1'h0, T36};
  assign T36 = T37 ? 3'h4 : 3'h0;
  assign T37 = ex_ctrl_fma & ex_ctrl_single;
  assign T38 = T109 | T39;
  assign T39 = ex_ctrl_fromint ? 4'h8 : 4'h0;
  assign T109 = {1'h0, T40};
  assign T40 = ex_ctrl_fastpipe ? 3'h4 : 3'h0;
  assign T110 = {2'h0, wen};
  assign T111 = reset ? 2'h0 : T41;
  assign T41 = T45 ? T43 : T112;
  assign T112 = {1'h0, T42};
  assign T42 = wen >> 1'h1;
  assign T43 = T113 | memLatencyMask;
  assign T113 = {1'h0, T44};
  assign T44 = wen >> 1'h1;
  assign T45 = mem_wen & T46;
  assign T46 = killm ^ 1'h1;
  assign killm = io_ctrl_killm | io_ctrl_nack_mem;
  assign T47 = mem_wen & T48;
  assign T48 = T49 != 3'h0;
  assign T49 = T116 & T50;
  assign T50 = T54 | T51;
  assign T51 = T52 ? 3'h4 : 3'h0;
  assign T52 = ex_ctrl_fma & T53;
  assign T53 = ex_ctrl_single ^ 1'h1;
  assign T54 = T57 | T114;
  assign T114 = {1'h0, T55};
  assign T55 = T56 ? 2'h2 : 2'h0;
  assign T56 = ex_ctrl_fma & ex_ctrl_single;
  assign T57 = T115 | T58;
  assign T58 = ex_ctrl_fromint ? 3'h4 : 3'h0;
  assign T115 = {1'h0, T59};
  assign T59 = ex_ctrl_fastpipe ? 2'h2 : 2'h0;
  assign T116 = {1'h0, memLatencyMask};
  assign mem_wen = mem_reg_valid & T60;
  assign T60 = T61 | mem_ctrl_fromint;
  assign T61 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T117 = reset ? 1'h0 : T62;
  assign T62 = ex_reg_valid & T63;
  assign T63 = io_ctrl_killx ^ 1'h1;
  assign T64 = wen[1'h1:1'h1];
  assign mem_winfo = {T68, T65};
  assign T65 = mem_reg_inst[4'hb:3'h7];
  assign T66 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T67 = io_ctrl_valid ? io_dpath_inst : ex_reg_inst;
  assign T68 = T72 | T69;
  assign T69 = T70 ? 2'h3 : 2'h0;
  assign T70 = mem_ctrl_fma & T71;
  assign T71 = mem_ctrl_single ^ 1'h1;
  assign T72 = T118 | T73;
  assign T73 = T74 ? 2'h2 : 2'h0;
  assign T74 = mem_ctrl_fma & mem_ctrl_single;
  assign T118 = {1'h0, T75};
  assign T75 = 1'h0 | mem_ctrl_fromint;
  assign T76 = mem_wen & T77;
  assign T77 = T79 & T78;
  assign T78 = memLatencyMask[1'h0:1'h0];
  assign T79 = write_port_busy ^ 1'h1;
  assign T126 = T129 ? T128 : T127;
  assign T127 = {32'hffffffff, sfma_io_out_bits_data};
  assign T128 = {32'h0, dfma_io_out_bits_data};
  assign T129 = T125[1'h0:1'h0];
  assign T130 = T125[1'h1:1'h1];
  assign T131 = wen[1'h0:1'h0];
  assign T132 = waddr[3'h4:1'h0];
  assign waddr = T93;
  assign T93 = winfo_0[3'h4:1'h0];
  assign load_wb_data_recoded = load_wb_single ? T293 : rec_d;
  assign rec_d = {T292, T134};
  assign T134 = {T270, T135};
  assign T135 = T268 ? T138 : T136;
  assign T136 = load_wb_data[6'h33:1'h0];
  assign T137 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_data : load_wb_data;
  assign T138 = T139[6'h3e:4'hb];
  assign T139 = T267 << T140;
  assign T140 = ~ T141;
  assign T141 = T266 ? 6'h3f : T142;
  assign T142 = T265 ? 6'h3e : T143;
  assign T143 = T264 ? 6'h3d : T144;
  assign T144 = T263 ? 6'h3c : T145;
  assign T145 = T262 ? 6'h3b : T146;
  assign T146 = T261 ? 6'h3a : T147;
  assign T147 = T260 ? 6'h39 : T148;
  assign T148 = T259 ? 6'h38 : T149;
  assign T149 = T258 ? 6'h37 : T150;
  assign T150 = T257 ? 6'h36 : T151;
  assign T151 = T256 ? 6'h35 : T152;
  assign T152 = T255 ? 6'h34 : T153;
  assign T153 = T254 ? 6'h33 : T154;
  assign T154 = T253 ? 6'h32 : T155;
  assign T155 = T252 ? 6'h31 : T156;
  assign T156 = T251 ? 6'h30 : T157;
  assign T157 = T250 ? 6'h2f : T158;
  assign T158 = T249 ? 6'h2e : T159;
  assign T159 = T248 ? 6'h2d : T160;
  assign T160 = T247 ? 6'h2c : T161;
  assign T161 = T246 ? 6'h2b : T162;
  assign T162 = T245 ? 6'h2a : T163;
  assign T163 = T244 ? 6'h29 : T164;
  assign T164 = T243 ? 6'h28 : T165;
  assign T165 = T242 ? 6'h27 : T166;
  assign T166 = T241 ? 6'h26 : T167;
  assign T167 = T240 ? 6'h25 : T168;
  assign T168 = T239 ? 6'h24 : T169;
  assign T169 = T238 ? 6'h23 : T170;
  assign T170 = T237 ? 6'h22 : T171;
  assign T171 = T236 ? 6'h21 : T172;
  assign T172 = T235 ? 6'h20 : T173;
  assign T173 = T234 ? 5'h1f : T174;
  assign T174 = T233 ? 5'h1e : T175;
  assign T175 = T232 ? 5'h1d : T176;
  assign T176 = T231 ? 5'h1c : T177;
  assign T177 = T230 ? 5'h1b : T178;
  assign T178 = T229 ? 5'h1a : T179;
  assign T179 = T228 ? 5'h19 : T180;
  assign T180 = T227 ? 5'h18 : T181;
  assign T181 = T226 ? 5'h17 : T182;
  assign T182 = T225 ? 5'h16 : T183;
  assign T183 = T224 ? 5'h15 : T184;
  assign T184 = T223 ? 5'h14 : T185;
  assign T185 = T222 ? 5'h13 : T186;
  assign T186 = T221 ? 5'h12 : T187;
  assign T187 = T220 ? 5'h11 : T188;
  assign T188 = T219 ? 5'h10 : T189;
  assign T189 = T218 ? 4'hf : T190;
  assign T190 = T217 ? 4'he : T191;
  assign T191 = T216 ? 4'hd : T192;
  assign T192 = T215 ? 4'hc : T193;
  assign T193 = T214 ? 4'hb : T194;
  assign T194 = T213 ? 4'ha : T195;
  assign T195 = T212 ? 4'h9 : T196;
  assign T196 = T211 ? 4'h8 : T197;
  assign T197 = T210 ? 3'h7 : T198;
  assign T198 = T209 ? 3'h6 : T199;
  assign T199 = T208 ? 3'h5 : T200;
  assign T200 = T207 ? 3'h4 : T201;
  assign T201 = T206 ? 2'h3 : T202;
  assign T202 = T205 ? 2'h2 : T203;
  assign T203 = T204[1'h1:1'h1];
  assign T204 = T267[6'h3f:1'h0];
  assign T205 = T204[2'h2:2'h2];
  assign T206 = T204[2'h3:2'h3];
  assign T207 = T204[3'h4:3'h4];
  assign T208 = T204[3'h5:3'h5];
  assign T209 = T204[3'h6:3'h6];
  assign T210 = T204[3'h7:3'h7];
  assign T211 = T204[4'h8:4'h8];
  assign T212 = T204[4'h9:4'h9];
  assign T213 = T204[4'ha:4'ha];
  assign T214 = T204[4'hb:4'hb];
  assign T215 = T204[4'hc:4'hc];
  assign T216 = T204[4'hd:4'hd];
  assign T217 = T204[4'he:4'he];
  assign T218 = T204[4'hf:4'hf];
  assign T219 = T204[5'h10:5'h10];
  assign T220 = T204[5'h11:5'h11];
  assign T221 = T204[5'h12:5'h12];
  assign T222 = T204[5'h13:5'h13];
  assign T223 = T204[5'h14:5'h14];
  assign T224 = T204[5'h15:5'h15];
  assign T225 = T204[5'h16:5'h16];
  assign T226 = T204[5'h17:5'h17];
  assign T227 = T204[5'h18:5'h18];
  assign T228 = T204[5'h19:5'h19];
  assign T229 = T204[5'h1a:5'h1a];
  assign T230 = T204[5'h1b:5'h1b];
  assign T231 = T204[5'h1c:5'h1c];
  assign T232 = T204[5'h1d:5'h1d];
  assign T233 = T204[5'h1e:5'h1e];
  assign T234 = T204[5'h1f:5'h1f];
  assign T235 = T204[6'h20:6'h20];
  assign T236 = T204[6'h21:6'h21];
  assign T237 = T204[6'h22:6'h22];
  assign T238 = T204[6'h23:6'h23];
  assign T239 = T204[6'h24:6'h24];
  assign T240 = T204[6'h25:6'h25];
  assign T241 = T204[6'h26:6'h26];
  assign T242 = T204[6'h27:6'h27];
  assign T243 = T204[6'h28:6'h28];
  assign T244 = T204[6'h29:6'h29];
  assign T245 = T204[6'h2a:6'h2a];
  assign T246 = T204[6'h2b:6'h2b];
  assign T247 = T204[6'h2c:6'h2c];
  assign T248 = T204[6'h2d:6'h2d];
  assign T249 = T204[6'h2e:6'h2e];
  assign T250 = T204[6'h2f:6'h2f];
  assign T251 = T204[6'h30:6'h30];
  assign T252 = T204[6'h31:6'h31];
  assign T253 = T204[6'h32:6'h32];
  assign T254 = T204[6'h33:6'h33];
  assign T255 = T204[6'h34:6'h34];
  assign T256 = T204[6'h35:6'h35];
  assign T257 = T204[6'h36:6'h36];
  assign T258 = T204[6'h37:6'h37];
  assign T259 = T204[6'h38:6'h38];
  assign T260 = T204[6'h39:6'h39];
  assign T261 = T204[6'h3a:6'h3a];
  assign T262 = T204[6'h3b:6'h3b];
  assign T263 = T204[6'h3c:6'h3c];
  assign T264 = T204[6'h3d:6'h3d];
  assign T265 = T204[6'h3e:6'h3e];
  assign T266 = T204[6'h3f:6'h3f];
  assign T267 = T136 << 4'hc;
  assign T268 = T269 == 11'h0;
  assign T269 = load_wb_data[6'h3e:6'h34];
  assign T270 = T278 | T271;
  assign T271 = {2'h0, T272};
  assign T272 = T273 << 4'h9;
  assign T273 = T276 & T274;
  assign T274 = T275 ^ 1'h1;
  assign T275 = T136 == 52'h0;
  assign T276 = T277 == 2'h3;
  assign T277 = T278[4'hb:4'ha];
  assign T278 = T287 + T279;
  assign T279 = {1'h0, T280};
  assign T280 = T286 ? 11'h0 : T281;
  assign T281 = 11'h400 | T282;
  assign T282 = {9'h0, T283};
  assign T283 = T284 ? 2'h2 : 2'h1;
  assign T284 = T268 & T285;
  assign T285 = T275 ^ 1'h1;
  assign T286 = T268 & T275;
  assign T287 = T268 ? T289 : T288;
  assign T288 = {1'h0, T269};
  assign T289 = T275 ? 12'h0 : T290;
  assign T290 = {6'h3f, T291};
  assign T291 = ~ T140;
  assign T292 = load_wb_data[6'h3f:6'h3f];
  assign T293 = {32'hffffffff, rec_s};
  assign rec_s = {T387, T294};
  assign T294 = {T365, T295};
  assign T295 = T363 ? T297 : T296;
  assign T296 = load_wb_data[5'h16:1'h0];
  assign T297 = T298[5'h1e:4'h8];
  assign T298 = T362 << T299;
  assign T299 = ~ T300;
  assign T300 = T361 ? 5'h1f : T301;
  assign T301 = T360 ? 5'h1e : T302;
  assign T302 = T359 ? 5'h1d : T303;
  assign T303 = T358 ? 5'h1c : T304;
  assign T304 = T357 ? 5'h1b : T305;
  assign T305 = T356 ? 5'h1a : T306;
  assign T306 = T355 ? 5'h19 : T307;
  assign T307 = T354 ? 5'h18 : T308;
  assign T308 = T353 ? 5'h17 : T309;
  assign T309 = T352 ? 5'h16 : T310;
  assign T310 = T351 ? 5'h15 : T311;
  assign T311 = T350 ? 5'h14 : T312;
  assign T312 = T349 ? 5'h13 : T313;
  assign T313 = T348 ? 5'h12 : T314;
  assign T314 = T347 ? 5'h11 : T315;
  assign T315 = T346 ? 5'h10 : T316;
  assign T316 = T345 ? 4'hf : T317;
  assign T317 = T344 ? 4'he : T318;
  assign T318 = T343 ? 4'hd : T319;
  assign T319 = T342 ? 4'hc : T320;
  assign T320 = T341 ? 4'hb : T321;
  assign T321 = T340 ? 4'ha : T322;
  assign T322 = T339 ? 4'h9 : T323;
  assign T323 = T338 ? 4'h8 : T324;
  assign T324 = T337 ? 3'h7 : T325;
  assign T325 = T336 ? 3'h6 : T326;
  assign T326 = T335 ? 3'h5 : T327;
  assign T327 = T334 ? 3'h4 : T328;
  assign T328 = T333 ? 2'h3 : T329;
  assign T329 = T332 ? 2'h2 : T330;
  assign T330 = T331[1'h1:1'h1];
  assign T331 = T362[5'h1f:1'h0];
  assign T332 = T331[2'h2:2'h2];
  assign T333 = T331[2'h3:2'h3];
  assign T334 = T331[3'h4:3'h4];
  assign T335 = T331[3'h5:3'h5];
  assign T336 = T331[3'h6:3'h6];
  assign T337 = T331[3'h7:3'h7];
  assign T338 = T331[4'h8:4'h8];
  assign T339 = T331[4'h9:4'h9];
  assign T340 = T331[4'ha:4'ha];
  assign T341 = T331[4'hb:4'hb];
  assign T342 = T331[4'hc:4'hc];
  assign T343 = T331[4'hd:4'hd];
  assign T344 = T331[4'he:4'he];
  assign T345 = T331[4'hf:4'hf];
  assign T346 = T331[5'h10:5'h10];
  assign T347 = T331[5'h11:5'h11];
  assign T348 = T331[5'h12:5'h12];
  assign T349 = T331[5'h13:5'h13];
  assign T350 = T331[5'h14:5'h14];
  assign T351 = T331[5'h15:5'h15];
  assign T352 = T331[5'h16:5'h16];
  assign T353 = T331[5'h17:5'h17];
  assign T354 = T331[5'h18:5'h18];
  assign T355 = T331[5'h19:5'h19];
  assign T356 = T331[5'h1a:5'h1a];
  assign T357 = T331[5'h1b:5'h1b];
  assign T358 = T331[5'h1c:5'h1c];
  assign T359 = T331[5'h1d:5'h1d];
  assign T360 = T331[5'h1e:5'h1e];
  assign T361 = T331[5'h1f:5'h1f];
  assign T362 = T296 << 4'h9;
  assign T363 = T364 == 8'h0;
  assign T364 = load_wb_data[5'h1e:5'h17];
  assign T365 = T373 | T366;
  assign T366 = {2'h0, T367};
  assign T367 = T368 << 3'h6;
  assign T368 = T371 & T369;
  assign T369 = T370 ^ 1'h1;
  assign T370 = T296 == 23'h0;
  assign T371 = T372 == 2'h3;
  assign T372 = T373[4'h8:3'h7];
  assign T373 = T382 + T374;
  assign T374 = {1'h0, T375};
  assign T375 = T381 ? 8'h0 : T376;
  assign T376 = 8'h80 | T377;
  assign T377 = {6'h0, T378};
  assign T378 = T379 ? 2'h2 : 2'h1;
  assign T379 = T363 & T380;
  assign T380 = T370 ^ 1'h1;
  assign T381 = T363 & T370;
  assign T382 = T363 ? T384 : T383;
  assign T383 = {1'h0, T364};
  assign T384 = T370 ? 9'h0 : T385;
  assign T385 = {4'hf, T386};
  assign T386 = ~ T299;
  assign T387 = load_wb_data[5'h1f:5'h1f];
  assign T388 = io_dpath_dmem_resp_val ? T389 : load_wb_single;
  assign T389 = T391 | T390;
  assign T390 = io_dpath_dmem_resp_type == 3'h6;
  assign T391 = io_dpath_dmem_resp_type == 3'h2;
  assign T392 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_tag : load_wb_tag;
  assign T393 = T398 ? T397 : T394;
  assign T394 = T396 ? T395 : ex_ra3;
  assign T395 = io_dpath_inst[5'h1f:5'h1b];
  assign T396 = io_ctrl_valid & fp_decoder_io_sigs_ren3;
  assign T397 = io_dpath_inst[5'h18:5'h14];
  assign T398 = T401 & T399;
  assign T399 = T400 & fp_decoder_io_sigs_swap23;
  assign T400 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign T401 = io_ctrl_valid & fp_decoder_io_sigs_ren2;
  assign req_in2 = ex_rs2;
  assign ex_rs2 = regfile[ex_ra2];
  assign T402 = T404 ? T403 : ex_ra2;
  assign T403 = io_dpath_inst[5'h18:5'h14];
  assign T404 = T401 & T405;
  assign T405 = T407 & T406;
  assign T406 = fp_decoder_io_sigs_swap23 ^ 1'h1;
  assign T407 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign req_in1 = ex_rs1;
  assign ex_rs1 = regfile[ex_ra1];
  assign T408 = T413 ? T412 : T409;
  assign T409 = T411 ? T410 : ex_ra1;
  assign T410 = io_dpath_inst[5'h13:4'hf];
  assign T411 = io_ctrl_valid & fp_decoder_io_sigs_ren1;
  assign T412 = io_dpath_inst[5'h18:5'h14];
  assign T413 = T401 & fp_decoder_io_sigs_ldst;
  assign req_typ = T414;
  assign T414 = ex_reg_inst[5'h15:5'h14];
  assign req_rm = ex_rm;
  assign ex_rm = T100 ? io_dpath_fcsr_rm : T99;
  assign T99 = ex_reg_inst[4'he:4'hc];
  assign T100 = T101 == 3'h7;
  assign T101 = ex_reg_inst[4'he:4'hc];
  assign req_round = ex_ctrl_round;
  assign T97 = io_ctrl_valid ? fp_decoder_io_sigs_round : ex_ctrl_round;
  assign req_fma = ex_ctrl_fma;
  assign req_fastpipe = ex_ctrl_fastpipe;
  assign req_toint = ex_ctrl_toint;
  assign T87 = io_ctrl_valid ? fp_decoder_io_sigs_toint : ex_ctrl_toint;
  assign req_fromint = ex_ctrl_fromint;
  assign req_single = ex_ctrl_single;
  assign req_swap23 = ex_ctrl_swap23;
  assign T415 = io_ctrl_valid ? fp_decoder_io_sigs_swap23 : ex_ctrl_swap23;
  assign req_ren3 = ex_ctrl_ren3;
  assign T416 = io_ctrl_valid ? fp_decoder_io_sigs_ren3 : ex_ctrl_ren3;
  assign req_ren2 = ex_ctrl_ren2;
  assign T417 = io_ctrl_valid ? fp_decoder_io_sigs_ren2 : ex_ctrl_ren2;
  assign req_ren1 = ex_ctrl_ren1;
  assign T418 = io_ctrl_valid ? fp_decoder_io_sigs_ren1 : ex_ctrl_ren1;
  assign req_wen = ex_ctrl_wen;
  assign T419 = io_ctrl_valid ? fp_decoder_io_sigs_wen : ex_ctrl_wen;
  assign req_ldst = ex_ctrl_ldst;
  assign T420 = io_ctrl_valid ? fp_decoder_io_sigs_ldst : ex_ctrl_ldst;
  assign req_cmd = ex_ctrl_cmd;
  assign T421 = io_ctrl_valid ? fp_decoder_io_sigs_cmd : ex_ctrl_cmd;
  assign T422 = ex_reg_valid & ex_ctrl_fastpipe;
  assign T423 = {1'h0, io_dpath_fromint_data};
  assign T424 = ex_reg_valid & ex_ctrl_fromint;
  assign T425 = ex_reg_valid & T426;
  assign T426 = ex_ctrl_toint | T427;
  assign T427 = T428 == 5'h5;
  assign T428 = ex_ctrl_cmd & 5'hd;
  assign T429 = T431 & T430;
  assign T430 = ex_ctrl_single ^ 1'h1;
  assign T431 = ex_reg_valid & ex_ctrl_fma;
  assign T432 = T433 & ex_ctrl_single;
  assign T433 = ex_reg_valid & ex_ctrl_fma;
  assign io_dpath_toint_data = fpiu_io_out_bits_toint;
  assign io_dpath_store_data = fpiu_io_out_bits_store;
  assign io_dpath_fcsr_flags_bits = T0;
  assign T0 = T84 | T1;
  assign T1 = T83 ? wexc : 5'h0;
  assign wexc = T82 ? T80 : T2;
  assign T2 = T3 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = wsrc;
  assign T80 = T81 ? dfma_io_out_bits_exc : sfma_io_out_bits_exc;
  assign T81 = T4[1'h0:1'h0];
  assign T82 = T4[1'h1:1'h1];
  assign T83 = wen[1'h0:1'h0];
  assign T84 = wb_toint_valid ? wb_toint_exc : 5'h0;
  assign T85 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign T86 = ex_reg_valid ? ex_ctrl_toint : mem_ctrl_toint;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign T88 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign T119 = reset ? 1'h0 : T89;
  assign T89 = mem_reg_valid & T90;
  assign T90 = killm ^ 1'h1;
  assign io_dpath_fcsr_flags_valid = T91;
  assign T91 = wb_toint_valid | T92;
  assign T92 = wen[1'h0:1'h0];
  assign io_ctrl_sboard_clra = waddr;
  assign io_ctrl_sboard_clr = 1'h0;
  assign io_ctrl_sboard_set = T94;
  assign T94 = wb_reg_valid & R95;
  assign io_ctrl_dec_round = fp_decoder_io_sigs_round;
  assign io_ctrl_dec_fma = fp_decoder_io_sigs_fma;
  assign io_ctrl_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_ctrl_dec_toint = fp_decoder_io_sigs_toint;
  assign io_ctrl_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_ctrl_dec_single = fp_decoder_io_sigs_single;
  assign io_ctrl_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_ctrl_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_ctrl_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_ctrl_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_ctrl_dec_wen = fp_decoder_io_sigs_wen;
  assign io_ctrl_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_ctrl_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_ctrl_illegal_rm = T96;
  assign T96 = T98 & ex_ctrl_round;
  assign T98 = ex_rm[2'h2:2'h2];
  assign io_ctrl_nack_mem = write_port_busy;
  assign io_ctrl_fcsr_rdy = T102;
  assign T102 = fp_inflight ^ 1'h1;
  assign fp_inflight = T104 | T103;
  assign T103 = wen != 2'h0;
  assign T104 = wb_reg_valid & wb_ctrl_toint;
  FPUDecoder fp_decoder(
       .io_inst( io_dpath_inst ),
       .io_sigs_cmd( fp_decoder_io_sigs_cmd ),
       .io_sigs_ldst( fp_decoder_io_sigs_ldst ),
       .io_sigs_wen( fp_decoder_io_sigs_wen ),
       .io_sigs_ren1( fp_decoder_io_sigs_ren1 ),
       .io_sigs_ren2( fp_decoder_io_sigs_ren2 ),
       .io_sigs_ren3( fp_decoder_io_sigs_ren3 ),
       .io_sigs_swap23( fp_decoder_io_sigs_swap23 ),
       .io_sigs_single( fp_decoder_io_sigs_single ),
       .io_sigs_fromint( fp_decoder_io_sigs_fromint ),
       .io_sigs_toint( fp_decoder_io_sigs_toint ),
       .io_sigs_fastpipe( fp_decoder_io_sigs_fastpipe ),
       .io_sigs_fma( fp_decoder_io_sigs_fma ),
       .io_sigs_round( fp_decoder_io_sigs_round )
  );
  FPUFMAPipe_0 sfma(.clk(clk), .reset(reset),
       .io_in_valid( T432 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( sfma_io_out_bits_data ),
       .io_out_bits_exc( sfma_io_out_bits_exc )
  );
  FPUFMAPipe_1 dfma(.clk(clk), .reset(reset),
       .io_in_valid( T429 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( dfma_io_out_bits_data ),
       .io_out_bits_exc( dfma_io_out_bits_exc )
  );
  FPToInt fpiu(.clk(clk),
       .io_in_valid( T425 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_lt( fpiu_io_out_bits_lt ),
       .io_out_bits_store( fpiu_io_out_bits_store ),
       .io_out_bits_toint( fpiu_io_out_bits_toint ),
       .io_out_bits_exc( fpiu_io_out_bits_exc )
  );
  IntToFP ifpu(.clk(clk), .reset(reset),
       .io_in_valid( T424 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( T423 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( ifpu_io_out_bits_data ),
       .io_out_bits_exc( ifpu_io_out_bits_exc )
  );
  FPToFP fpmu(.clk(clk), .reset(reset),
       .io_in_valid( T422 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( fpmu_io_out_bits_data ),
       .io_out_bits_exc( fpmu_io_out_bits_exc ),
       .io_lt( fpiu_io_out_bits_lt )
  );

  always @(posedge clk) begin
    if (T131)
      regfile[T132] <= T121;
    if(T76) begin
      winfo_0 <= mem_winfo;
    end else if(T64) begin
      winfo_0 <= winfo_1;
    end
    if(T8) begin
      winfo_1 <= mem_winfo;
    end
    if(ex_reg_valid) begin
      mem_ctrl_single <= ex_ctrl_single;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_single <= fp_decoder_io_sigs_single;
    end
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_ctrl_valid;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fma <= ex_ctrl_fma;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fromint <= ex_ctrl_fromint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_ctrl_fastpipe;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if(ex_reg_valid) begin
      write_port_busy <= T28;
    end
    if(reset) begin
      wen <= 2'h0;
    end else if(T45) begin
      wen <= T43;
    end else begin
      wen <= T112;
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T62;
    end
    if(ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(io_ctrl_valid) begin
      ex_reg_inst <= io_dpath_inst;
    end
    if (load_wb)
      regfile[load_wb_tag] <= load_wb_data_recoded;
    if(io_dpath_dmem_resp_val) begin
      load_wb_data <= io_dpath_dmem_resp_data;
    end
    if(io_dpath_dmem_resp_val) begin
      load_wb_single <= T389;
    end
    load_wb <= io_dpath_dmem_resp_val;
    if(io_dpath_dmem_resp_val) begin
      load_wb_tag <= io_dpath_dmem_resp_tag;
    end
    if(T398) begin
      ex_ra3 <= T397;
    end else if(T396) begin
      ex_ra3 <= T395;
    end
    if(T404) begin
      ex_ra2 <= T403;
    end
    if(T413) begin
      ex_ra1 <= T412;
    end else if(T411) begin
      ex_ra1 <= T410;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_round <= fp_decoder_io_sigs_round;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren1 <= fp_decoder_io_sigs_ren1;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_wen <= fp_decoder_io_sigs_wen;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ldst <= fp_decoder_io_sigs_ldst;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_cmd <= fp_decoder_io_sigs_cmd;
    end
    if(mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if(ex_reg_valid) begin
      mem_ctrl_toint <= ex_ctrl_toint;
    end
    if(mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T89;
    end
    R95 <= 1'h0;
  end
endmodule

module Core(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[43:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_mispredict,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output[43:0] io_dmem_req_bits_addr,
    output[8:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [8:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [8:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    output io_rocc_resp_ready,
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [2:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [511:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[2:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready,
    output io_temac_sfp_tx_disable
);

  wire[2:0] ctrl_io_dpath_sel_pc;
  wire ctrl_io_dpath_killd;
  wire ctrl_io_dpath_ren_1;
  wire ctrl_io_dpath_ren_0;
  wire[2:0] ctrl_io_dpath_sel_alu2;
  wire[1:0] ctrl_io_dpath_sel_alu1;
  wire[2:0] ctrl_io_dpath_sel_imm;
  wire ctrl_io_dpath_fn_dw;
  wire[3:0] ctrl_io_dpath_fn_alu;
  wire ctrl_io_dpath_div_mul_val;
  wire ctrl_io_dpath_div_mul_kill;
  wire[2:0] ctrl_io_dpath_csr;
  wire ctrl_io_dpath_sret;
  wire ctrl_io_dpath_mem_load;
  wire ctrl_io_dpath_wb_load;
  wire ctrl_io_dpath_ex_fp_val;
  wire ctrl_io_dpath_mem_fp_val;
  wire ctrl_io_dpath_ex_wen;
  wire ctrl_io_dpath_ex_valid;
  wire ctrl_io_dpath_mem_jalr;
  wire ctrl_io_dpath_mem_branch;
  wire ctrl_io_dpath_mem_wen;
  wire ctrl_io_dpath_wb_wen;
  wire[2:0] ctrl_io_dpath_ex_mem_type;
  wire ctrl_io_dpath_ex_rs2_val;
  wire ctrl_io_dpath_ex_rocc_val;
  wire ctrl_io_dpath_mem_rocc_val;
  wire ctrl_io_dpath_bypass_1;
  wire ctrl_io_dpath_bypass_0;
  wire[1:0] ctrl_io_dpath_bypass_src_1;
  wire[1:0] ctrl_io_dpath_bypass_src_0;
  wire ctrl_io_dpath_ll_ready;
  wire ctrl_io_dpath_retire;
  wire ctrl_io_dpath_exception;
  wire[63:0] ctrl_io_dpath_cause;
  wire ctrl_io_dpath_badvaddr_wen;
  wire ctrl_io_imem_req_valid;
  wire ctrl_io_imem_resp_ready;
  wire ctrl_io_imem_btb_update_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  wire[42:0] ctrl_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire ctrl_io_imem_btb_update_bits_taken;
  wire ctrl_io_imem_btb_update_bits_isJump;
  wire ctrl_io_imem_btb_update_bits_isCall;
  wire ctrl_io_imem_btb_update_bits_isReturn;
  wire ctrl_io_imem_btb_update_bits_mispredict;
  wire ctrl_io_imem_invalidate;
  wire ctrl_io_dmem_req_valid;
  wire ctrl_io_dmem_req_bits_kill;
  wire[2:0] ctrl_io_dmem_req_bits_typ;
  wire ctrl_io_dmem_req_bits_phys;
  wire[4:0] ctrl_io_dmem_req_bits_cmd;
  wire ctrl_io_fpu_valid;
  wire ctrl_io_fpu_killx;
  wire ctrl_io_fpu_killm;
  wire ctrl_io_rocc_cmd_valid;
  wire ctrl_io_rocc_s;
  wire ctrl_io_rocc_exception;
  wire dpath_io_host_pcr_req_ready;
  wire dpath_io_host_pcr_rep_valid;
  wire[63:0] dpath_io_host_pcr_rep_bits;
  wire dpath_io_host_ipi_req_valid;
  wire dpath_io_host_ipi_req_bits;
  wire dpath_io_host_ipi_rep_ready;
  wire dpath_io_host_debug_stats_pcr;
  wire[31:0] dpath_io_ctrl_inst;
  wire dpath_io_ctrl_mem_br_taken;
  wire dpath_io_ctrl_mem_misprediction;
  wire dpath_io_ctrl_div_mul_rdy;
  wire dpath_io_ctrl_ll_wen;
  wire[4:0] dpath_io_ctrl_ll_waddr;
  wire[4:0] dpath_io_ctrl_ex_waddr;
  wire dpath_io_ctrl_mem_rs1_ra;
  wire[4:0] dpath_io_ctrl_mem_waddr;
  wire[4:0] dpath_io_ctrl_wb_waddr;
  wire[7:0] dpath_io_ctrl_status_ip;
  wire[7:0] dpath_io_ctrl_status_im;
  wire[6:0] dpath_io_ctrl_status_zero;
  wire dpath_io_ctrl_status_er;
  wire dpath_io_ctrl_status_vm;
  wire dpath_io_ctrl_status_s64;
  wire dpath_io_ctrl_status_u64;
  wire dpath_io_ctrl_status_ef;
  wire dpath_io_ctrl_status_pei;
  wire dpath_io_ctrl_status_ei;
  wire dpath_io_ctrl_status_ps;
  wire dpath_io_ctrl_status_s;
  wire dpath_io_ctrl_fp_sboard_clr;
  wire[4:0] dpath_io_ctrl_fp_sboard_clra;
  wire dpath_io_ctrl_csr_replay;
  wire[43:0] dpath_io_dmem_req_bits_addr;
  wire[8:0] dpath_io_dmem_req_bits_tag;
  wire[63:0] dpath_io_dmem_req_bits_data;
  wire[31:0] dpath_io_ptw_ptbr;
  wire dpath_io_ptw_invalidate;
  wire dpath_io_ptw_sret;
  wire[7:0] dpath_io_ptw_status_ip;
  wire[7:0] dpath_io_ptw_status_im;
  wire[6:0] dpath_io_ptw_status_zero;
  wire dpath_io_ptw_status_er;
  wire dpath_io_ptw_status_vm;
  wire dpath_io_ptw_status_s64;
  wire dpath_io_ptw_status_u64;
  wire dpath_io_ptw_status_ef;
  wire dpath_io_ptw_status_pei;
  wire dpath_io_ptw_status_ei;
  wire dpath_io_ptw_status_ps;
  wire dpath_io_ptw_status_s;
  wire[43:0] dpath_io_imem_req_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_target;
  wire[42:0] dpath_io_imem_btb_update_bits_returnAddr;
  wire[31:0] dpath_io_fpu_inst;
  wire[63:0] dpath_io_fpu_fromint_data;
  wire[2:0] dpath_io_fpu_fcsr_rm;
  wire dpath_io_fpu_dmem_resp_val;
  wire[2:0] dpath_io_fpu_dmem_resp_type;
  wire[4:0] dpath_io_fpu_dmem_resp_tag;
  wire[63:0] dpath_io_fpu_dmem_resp_data;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_funct;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs1;
  wire dpath_io_rocc_cmd_bits_inst_xd;
  wire dpath_io_rocc_cmd_bits_inst_xs1;
  wire dpath_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rd;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] dpath_io_rocc_cmd_bits_rs1;
  wire[63:0] dpath_io_rocc_cmd_bits_rs2;
  wire dpath_io_rocc_resp_ready;
  wire dpath_io_temac_rx_axis_fifo_tready;
  wire[7:0] dpath_io_temac_tx_axis_fifo_tdata;
  wire dpath_io_temac_tx_axis_fifo_tvalid;
  wire dpath_io_temac_tx_axis_fifo_tlast;
  wire[11:0] dpath_io_temac_s_axi_awaddr;
  wire dpath_io_temac_s_axi_awvalid;
  wire[31:0] dpath_io_temac_s_axi_wdata;
  wire dpath_io_temac_s_axi_wvalid;
  wire dpath_io_temac_s_axi_bready;
  wire[11:0] dpath_io_temac_s_axi_araddr;
  wire dpath_io_temac_s_axi_arvalid;
  wire dpath_io_temac_s_axi_rready;
  wire dpath_io_temac_sfp_tx_disable;
  wire FPU_io_ctrl_fcsr_rdy;
  wire FPU_io_ctrl_nack_mem;
  wire FPU_io_ctrl_illegal_rm;
  wire[4:0] FPU_io_ctrl_dec_cmd;
  wire FPU_io_ctrl_dec_ldst;
  wire FPU_io_ctrl_dec_wen;
  wire FPU_io_ctrl_dec_ren1;
  wire FPU_io_ctrl_dec_ren2;
  wire FPU_io_ctrl_dec_ren3;
  wire FPU_io_ctrl_dec_swap23;
  wire FPU_io_ctrl_dec_single;
  wire FPU_io_ctrl_dec_fromint;
  wire FPU_io_ctrl_dec_toint;
  wire FPU_io_ctrl_dec_fastpipe;
  wire FPU_io_ctrl_dec_fma;
  wire FPU_io_ctrl_dec_round;
  wire FPU_io_ctrl_sboard_set;
  wire FPU_io_ctrl_sboard_clr;
  wire[4:0] FPU_io_ctrl_sboard_clra;
  wire FPU_io_dpath_fcsr_flags_valid;
  wire[4:0] FPU_io_dpath_fcsr_flags_bits;
  wire[63:0] FPU_io_dpath_store_data;
  wire[63:0] FPU_io_dpath_toint_data;


  assign io_temac_sfp_tx_disable = dpath_io_temac_sfp_tx_disable;
  assign io_temac_s_axi_rready = dpath_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = dpath_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = dpath_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = dpath_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = dpath_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = dpath_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = dpath_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = dpath_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = dpath_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = dpath_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = dpath_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = dpath_io_temac_rx_axis_fifo_tready;
  assign io_rocc_exception = ctrl_io_rocc_exception;
  assign io_rocc_s = ctrl_io_rocc_s;
  assign io_rocc_resp_ready = dpath_io_rocc_resp_ready;
  assign io_rocc_cmd_bits_rs2 = dpath_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = dpath_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = dpath_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = dpath_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = dpath_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = dpath_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = dpath_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = dpath_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = dpath_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = dpath_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = ctrl_io_rocc_cmd_valid;
  assign io_ptw_status_s = dpath_io_ptw_status_s;
  assign io_ptw_status_ps = dpath_io_ptw_status_ps;
  assign io_ptw_status_ei = dpath_io_ptw_status_ei;
  assign io_ptw_status_pei = dpath_io_ptw_status_pei;
  assign io_ptw_status_ef = dpath_io_ptw_status_ef;
  assign io_ptw_status_u64 = dpath_io_ptw_status_u64;
  assign io_ptw_status_s64 = dpath_io_ptw_status_s64;
  assign io_ptw_status_vm = dpath_io_ptw_status_vm;
  assign io_ptw_status_er = dpath_io_ptw_status_er;
  assign io_ptw_status_zero = dpath_io_ptw_status_zero;
  assign io_ptw_status_im = dpath_io_ptw_status_im;
  assign io_ptw_status_ip = dpath_io_ptw_status_ip;
  assign io_ptw_sret = dpath_io_ptw_sret;
  assign io_ptw_invalidate = dpath_io_ptw_invalidate;
  assign io_ptw_ptbr = dpath_io_ptw_ptbr;
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_cmd = ctrl_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_tag = dpath_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_phys = ctrl_io_dmem_req_bits_phys;
  assign io_dmem_req_bits_typ = ctrl_io_dmem_req_bits_typ;
  assign io_dmem_req_bits_kill = ctrl_io_dmem_req_bits_kill;
  assign io_dmem_req_valid = ctrl_io_dmem_req_valid;
  assign io_imem_invalidate = ctrl_io_imem_invalidate;
  assign io_imem_btb_update_bits_mispredict = ctrl_io_imem_btb_update_bits_mispredict;
  assign io_imem_btb_update_bits_isReturn = ctrl_io_imem_btb_update_bits_isReturn;
  assign io_imem_btb_update_bits_isCall = ctrl_io_imem_btb_update_bits_isCall;
  assign io_imem_btb_update_bits_isJump = ctrl_io_imem_btb_update_bits_isJump;
  assign io_imem_btb_update_bits_taken = ctrl_io_imem_btb_update_bits_taken;
  assign io_imem_btb_update_bits_returnAddr = dpath_io_imem_btb_update_bits_returnAddr;
  assign io_imem_btb_update_bits_target = dpath_io_imem_btb_update_bits_target;
  assign io_imem_btb_update_bits_pc = dpath_io_imem_btb_update_bits_pc;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = ctrl_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = ctrl_io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_btb_update_bits_prediction_valid = ctrl_io_imem_btb_update_bits_prediction_valid;
  assign io_imem_btb_update_valid = ctrl_io_imem_btb_update_valid;
  assign io_imem_resp_ready = ctrl_io_imem_resp_ready;
  assign io_imem_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign io_imem_req_valid = ctrl_io_imem_req_valid;
  assign io_host_debug_stats_pcr = dpath_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = dpath_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = dpath_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = dpath_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = dpath_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = dpath_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = dpath_io_host_pcr_req_ready;
  Control ctrl(.clk(clk), .reset(reset),
       .io_dpath_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_dpath_killd( ctrl_io_dpath_killd ),
       .io_dpath_ren_1( ctrl_io_dpath_ren_1 ),
       .io_dpath_ren_0( ctrl_io_dpath_ren_0 ),
       .io_dpath_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_dpath_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_dpath_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_dpath_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_dpath_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_dpath_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_dpath_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_dpath_div_val(  )
       //.io_dpath_div_kill(  )
       .io_dpath_csr( ctrl_io_dpath_csr ),
       .io_dpath_sret( ctrl_io_dpath_sret ),
       .io_dpath_mem_load( ctrl_io_dpath_mem_load ),
       .io_dpath_wb_load( ctrl_io_dpath_wb_load ),
       .io_dpath_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_dpath_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_dpath_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_dpath_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_dpath_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_dpath_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_dpath_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_dpath_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_dpath_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_dpath_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_dpath_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_dpath_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_dpath_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_dpath_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_dpath_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_dpath_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_dpath_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_dpath_retire( ctrl_io_dpath_retire ),
       .io_dpath_exception( ctrl_io_dpath_exception ),
       .io_dpath_cause( ctrl_io_dpath_cause ),
       .io_dpath_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_dpath_inst( dpath_io_ctrl_inst ),
       //.io_dpath_jalr_eq(  )
       .io_dpath_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_dpath_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_dpath_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_dpath_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_dpath_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_dpath_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_dpath_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_dpath_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_dpath_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_dpath_status_ip( dpath_io_ctrl_status_ip ),
       .io_dpath_status_im( dpath_io_ctrl_status_im ),
       .io_dpath_status_zero( dpath_io_ctrl_status_zero ),
       .io_dpath_status_er( dpath_io_ctrl_status_er ),
       .io_dpath_status_vm( dpath_io_ctrl_status_vm ),
       .io_dpath_status_s64( dpath_io_ctrl_status_s64 ),
       .io_dpath_status_u64( dpath_io_ctrl_status_u64 ),
       .io_dpath_status_ef( dpath_io_ctrl_status_ef ),
       .io_dpath_status_pei( dpath_io_ctrl_status_pei ),
       .io_dpath_status_ei( dpath_io_ctrl_status_ei ),
       .io_dpath_status_ps( dpath_io_ctrl_status_ps ),
       .io_dpath_status_s( dpath_io_ctrl_status_s ),
       .io_dpath_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_dpath_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_dpath_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_imem_req_valid( ctrl_io_imem_req_valid ),
       //.io_imem_req_bits_pc(  )
       .io_imem_resp_ready( ctrl_io_imem_resp_ready ),
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( io_imem_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( ctrl_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( ctrl_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( ctrl_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( ctrl_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( ctrl_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( ctrl_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( ctrl_io_imem_btb_update_bits_prediction_bits_bht_value ),
       //.io_imem_btb_update_bits_pc(  )
       //.io_imem_btb_update_bits_target(  )
       //.io_imem_btb_update_bits_returnAddr(  )
       .io_imem_btb_update_bits_taken( ctrl_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( ctrl_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( ctrl_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( ctrl_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_mispredict( ctrl_io_imem_btb_update_bits_mispredict ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( ctrl_io_imem_invalidate ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       .io_dmem_req_valid( ctrl_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( ctrl_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( ctrl_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( ctrl_io_dmem_req_bits_phys ),
       //.io_dmem_req_bits_addr(  )
       //.io_dmem_req_bits_tag(  )
       .io_dmem_req_bits_cmd( ctrl_io_dmem_req_bits_cmd ),
       //.io_dmem_req_bits_data(  )
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_fpu_valid( ctrl_io_fpu_valid ),
       .io_fpu_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_fpu_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_fpu_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_fpu_killx( ctrl_io_fpu_killx ),
       .io_fpu_killm( ctrl_io_fpu_killm ),
       .io_fpu_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_fpu_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_fpu_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_fpu_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_fpu_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_fpu_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_fpu_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_fpu_dec_single( FPU_io_ctrl_dec_single ),
       .io_fpu_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_fpu_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_fpu_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_fpu_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_fpu_dec_round( FPU_io_ctrl_dec_round ),
       .io_fpu_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_fpu_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_fpu_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( ctrl_io_rocc_cmd_valid ),
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( ctrl_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( ctrl_io_rocc_exception )
  );
  Datapath dpath(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( dpath_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( dpath_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( dpath_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( dpath_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( dpath_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( dpath_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( dpath_io_host_debug_stats_pcr ),
       .io_ctrl_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_ctrl_killd( ctrl_io_dpath_killd ),
       .io_ctrl_ren_1( ctrl_io_dpath_ren_1 ),
       .io_ctrl_ren_0( ctrl_io_dpath_ren_0 ),
       .io_ctrl_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_ctrl_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_ctrl_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_ctrl_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_ctrl_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_ctrl_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_ctrl_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_ctrl_div_val(  )
       //.io_ctrl_div_kill(  )
       .io_ctrl_csr( ctrl_io_dpath_csr ),
       .io_ctrl_sret( ctrl_io_dpath_sret ),
       .io_ctrl_mem_load( ctrl_io_dpath_mem_load ),
       .io_ctrl_wb_load( ctrl_io_dpath_wb_load ),
       .io_ctrl_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_ctrl_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_ctrl_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_ctrl_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_ctrl_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_ctrl_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_ctrl_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_ctrl_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_ctrl_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_ctrl_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_ctrl_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_ctrl_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_ctrl_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_ctrl_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_ctrl_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_ctrl_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_ctrl_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_ctrl_retire( ctrl_io_dpath_retire ),
       .io_ctrl_exception( ctrl_io_dpath_exception ),
       .io_ctrl_cause( ctrl_io_dpath_cause ),
       .io_ctrl_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_ctrl_inst( dpath_io_ctrl_inst ),
       //.io_ctrl_jalr_eq(  )
       .io_ctrl_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_ctrl_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_ctrl_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_ctrl_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_ctrl_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_ctrl_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_ctrl_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_ctrl_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_ctrl_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_ctrl_status_ip( dpath_io_ctrl_status_ip ),
       .io_ctrl_status_im( dpath_io_ctrl_status_im ),
       .io_ctrl_status_zero( dpath_io_ctrl_status_zero ),
       .io_ctrl_status_er( dpath_io_ctrl_status_er ),
       .io_ctrl_status_vm( dpath_io_ctrl_status_vm ),
       .io_ctrl_status_s64( dpath_io_ctrl_status_s64 ),
       .io_ctrl_status_u64( dpath_io_ctrl_status_u64 ),
       .io_ctrl_status_ef( dpath_io_ctrl_status_ef ),
       .io_ctrl_status_pei( dpath_io_ctrl_status_pei ),
       .io_ctrl_status_ei( dpath_io_ctrl_status_ei ),
       .io_ctrl_status_ps( dpath_io_ctrl_status_ps ),
       .io_ctrl_status_s( dpath_io_ctrl_status_s ),
       .io_ctrl_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_ctrl_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_ctrl_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       //.io_dmem_req_valid(  )
       //.io_dmem_req_bits_kill(  )
       //.io_dmem_req_bits_typ(  )
       //.io_dmem_req_bits_phys(  )
       .io_dmem_req_bits_addr( dpath_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( dpath_io_dmem_req_bits_tag ),
       //.io_dmem_req_bits_cmd(  )
       .io_dmem_req_bits_data( dpath_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_ptw_ptbr( dpath_io_ptw_ptbr ),
       .io_ptw_invalidate( dpath_io_ptw_invalidate ),
       .io_ptw_sret( dpath_io_ptw_sret ),
       .io_ptw_status_ip( dpath_io_ptw_status_ip ),
       .io_ptw_status_im( dpath_io_ptw_status_im ),
       .io_ptw_status_zero( dpath_io_ptw_status_zero ),
       .io_ptw_status_er( dpath_io_ptw_status_er ),
       .io_ptw_status_vm( dpath_io_ptw_status_vm ),
       .io_ptw_status_s64( dpath_io_ptw_status_s64 ),
       .io_ptw_status_u64( dpath_io_ptw_status_u64 ),
       .io_ptw_status_ef( dpath_io_ptw_status_ef ),
       .io_ptw_status_pei( dpath_io_ptw_status_pei ),
       .io_ptw_status_ei( dpath_io_ptw_status_ei ),
       .io_ptw_status_ps( dpath_io_ptw_status_ps ),
       .io_ptw_status_s( dpath_io_ptw_status_s ),
       //.io_imem_req_valid(  )
       .io_imem_req_bits_pc( dpath_io_imem_req_bits_pc ),
       //.io_imem_resp_ready(  )
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( io_imem_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       //.io_imem_btb_update_valid(  )
       //.io_imem_btb_update_bits_prediction_valid(  )
       //.io_imem_btb_update_bits_prediction_bits_taken(  )
       //.io_imem_btb_update_bits_prediction_bits_target(  )
       //.io_imem_btb_update_bits_prediction_bits_entry(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_history(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_value(  )
       .io_imem_btb_update_bits_pc( dpath_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( dpath_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( dpath_io_imem_btb_update_bits_returnAddr ),
       //.io_imem_btb_update_bits_taken(  )
       //.io_imem_btb_update_bits_isJump(  )
       //.io_imem_btb_update_bits_isCall(  )
       //.io_imem_btb_update_bits_isReturn(  )
       //.io_imem_btb_update_bits_mispredict(  )
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       //.io_imem_invalidate(  )
       .io_fpu_inst( dpath_io_fpu_inst ),
       .io_fpu_fromint_data( dpath_io_fpu_fromint_data ),
       .io_fpu_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_fpu_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_fpu_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_fpu_store_data( FPU_io_dpath_store_data ),
       .io_fpu_toint_data( FPU_io_dpath_toint_data ),
       .io_fpu_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_fpu_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_fpu_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_fpu_dmem_resp_data( dpath_io_fpu_dmem_resp_data ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       .io_rocc_cmd_bits_inst_funct( dpath_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( dpath_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( dpath_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( dpath_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( dpath_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( dpath_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( dpath_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( dpath_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( dpath_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( dpath_io_rocc_cmd_bits_rs2 ),
       .io_rocc_resp_ready( dpath_io_rocc_resp_ready ),
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( dpath_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( dpath_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( dpath_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( dpath_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( dpath_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( dpath_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( dpath_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( dpath_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( dpath_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( dpath_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( dpath_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( dpath_io_temac_s_axi_rready ),
       .io_temac_sfp_tx_disable( dpath_io_temac_sfp_tx_disable )
  );
  FPU FPU(.clk(clk), .reset(reset),
       .io_ctrl_valid( ctrl_io_fpu_valid ),
       .io_ctrl_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_ctrl_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_ctrl_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_ctrl_killx( ctrl_io_fpu_killx ),
       .io_ctrl_killm( ctrl_io_fpu_killm ),
       .io_ctrl_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_ctrl_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_ctrl_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_ctrl_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_ctrl_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_ctrl_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_ctrl_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_ctrl_dec_single( FPU_io_ctrl_dec_single ),
       .io_ctrl_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_ctrl_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_ctrl_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_ctrl_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_ctrl_dec_round( FPU_io_ctrl_dec_round ),
       .io_ctrl_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_ctrl_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_ctrl_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_dpath_inst( dpath_io_fpu_inst ),
       .io_dpath_fromint_data( dpath_io_fpu_fromint_data ),
       .io_dpath_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_dpath_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_dpath_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_dpath_store_data( FPU_io_dpath_store_data ),
       .io_dpath_toint_data( FPU_io_dpath_toint_data ),
       .io_dpath_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_dpath_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_dpath_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_dpath_dmem_resp_data( dpath_io_fpu_dmem_resp_data )
  );
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_2_req_ready,
    input  io_requestor_2_req_valid,
    input  io_requestor_2_req_bits_kill,
    input [2:0] io_requestor_2_req_bits_typ,
    input  io_requestor_2_req_bits_phys,
    input [43:0] io_requestor_2_req_bits_addr,
    input [8:0] io_requestor_2_req_bits_tag,
    input [4:0] io_requestor_2_req_bits_cmd,
    input [63:0] io_requestor_2_req_bits_data,
    output io_requestor_2_resp_valid,
    output[63:0] io_requestor_2_resp_bits_data,
    output io_requestor_2_resp_bits_nack,
    output io_requestor_2_resp_bits_replay,
    output[2:0] io_requestor_2_resp_bits_typ,
    output io_requestor_2_resp_bits_has_data,
    output[63:0] io_requestor_2_resp_bits_data_subword,
    output[8:0] io_requestor_2_resp_bits_tag,
    output[3:0] io_requestor_2_resp_bits_cmd,
    output[43:0] io_requestor_2_resp_bits_addr,
    output[63:0] io_requestor_2_resp_bits_store_data,
    output io_requestor_2_replay_next_valid,
    output[8:0] io_requestor_2_replay_next_bits,
    output io_requestor_2_xcpt_ma_ld,
    output io_requestor_2_xcpt_ma_st,
    output io_requestor_2_xcpt_pf_ld,
    output io_requestor_2_xcpt_pf_st,
    //input  io_requestor_2_ptw_req_ready
    //output io_requestor_2_ptw_req_valid
    //output[29:0] io_requestor_2_ptw_req_bits
    //input  io_requestor_2_ptw_resp_valid
    //input  io_requestor_2_ptw_resp_bits_error
    //input [18:0] io_requestor_2_ptw_resp_bits_ppn
    //input [5:0] io_requestor_2_ptw_resp_bits_perm
    //input [7:0] io_requestor_2_ptw_status_ip
    //input [7:0] io_requestor_2_ptw_status_im
    //input [6:0] io_requestor_2_ptw_status_zero
    //input  io_requestor_2_ptw_status_er
    //input  io_requestor_2_ptw_status_vm
    //input  io_requestor_2_ptw_status_s64
    //input  io_requestor_2_ptw_status_u64
    //input  io_requestor_2_ptw_status_ef
    //input  io_requestor_2_ptw_status_pei
    //input  io_requestor_2_ptw_status_ei
    //input  io_requestor_2_ptw_status_ps
    //input  io_requestor_2_ptw_status_s
    //input  io_requestor_2_ptw_invalidate
    //input  io_requestor_2_ptw_sret
    output io_requestor_2_ordered,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input  io_requestor_1_req_bits_kill,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_phys,
    input [43:0] io_requestor_1_req_bits_addr,
    input [8:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    input [63:0] io_requestor_1_req_bits_data,
    output io_requestor_1_resp_valid,
    output[63:0] io_requestor_1_resp_bits_data,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output[2:0] io_requestor_1_resp_bits_typ,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[8:0] io_requestor_1_resp_bits_tag,
    output[3:0] io_requestor_1_resp_bits_cmd,
    output[43:0] io_requestor_1_resp_bits_addr,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[8:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    //input  io_requestor_1_ptw_req_ready
    //output io_requestor_1_ptw_req_valid
    //output[29:0] io_requestor_1_ptw_req_bits
    //input  io_requestor_1_ptw_resp_valid
    //input  io_requestor_1_ptw_resp_bits_error
    //input [18:0] io_requestor_1_ptw_resp_bits_ppn
    //input [5:0] io_requestor_1_ptw_resp_bits_perm
    //input [7:0] io_requestor_1_ptw_status_ip
    //input [7:0] io_requestor_1_ptw_status_im
    //input [6:0] io_requestor_1_ptw_status_zero
    //input  io_requestor_1_ptw_status_er
    //input  io_requestor_1_ptw_status_vm
    //input  io_requestor_1_ptw_status_s64
    //input  io_requestor_1_ptw_status_u64
    //input  io_requestor_1_ptw_status_ef
    //input  io_requestor_1_ptw_status_pei
    //input  io_requestor_1_ptw_status_ei
    //input  io_requestor_1_ptw_status_ps
    //input  io_requestor_1_ptw_status_s
    //input  io_requestor_1_ptw_invalidate
    //input  io_requestor_1_ptw_sret
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input  io_requestor_0_req_bits_kill,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_phys,
    input [43:0] io_requestor_0_req_bits_addr,
    input [8:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    input [63:0] io_requestor_0_req_bits_data,
    output io_requestor_0_resp_valid,
    output[63:0] io_requestor_0_resp_bits_data,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output[2:0] io_requestor_0_resp_bits_typ,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[8:0] io_requestor_0_resp_bits_tag,
    output[3:0] io_requestor_0_resp_bits_cmd,
    output[43:0] io_requestor_0_resp_bits_addr,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[8:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_ptw_req_ready
    //output io_requestor_0_ptw_req_valid
    //output[29:0] io_requestor_0_ptw_req_bits
    //input  io_requestor_0_ptw_resp_valid
    //input  io_requestor_0_ptw_resp_bits_error
    //input [18:0] io_requestor_0_ptw_resp_bits_ppn
    //input [5:0] io_requestor_0_ptw_resp_bits_perm
    //input [7:0] io_requestor_0_ptw_status_ip
    //input [7:0] io_requestor_0_ptw_status_im
    //input [6:0] io_requestor_0_ptw_status_zero
    //input  io_requestor_0_ptw_status_er
    //input  io_requestor_0_ptw_status_vm
    //input  io_requestor_0_ptw_status_s64
    //input  io_requestor_0_ptw_status_u64
    //input  io_requestor_0_ptw_status_ef
    //input  io_requestor_0_ptw_status_pei
    //input  io_requestor_0_ptw_status_ei
    //input  io_requestor_0_ptw_status_ps
    //input  io_requestor_0_ptw_status_s
    //input  io_requestor_0_ptw_invalidate
    //input  io_requestor_0_ptw_sret
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    output[8:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [8:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered
);

  wire[63:0] T0;
  wire[63:0] T1;
  reg  r_valid_1;
  reg  r_valid_0;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[8:0] T53;
  wire[10:0] T4;
  wire[10:0] T5;
  wire[10:0] T6;
  wire[10:0] T7;
  wire[10:0] T8;
  wire[43:0] T9;
  wire[43:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[8:0] T54;
  wire[6:0] T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire[8:0] T55;
  wire[6:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[8:0] T56;
  wire[6:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[8:0] T57;
  wire[6:0] T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[8:0] T58;
  wire[6:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[8:0] T59;
  wire[6:0] T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_valid_1 = {1{$random}};
    r_valid_0 = {1{$random}};
  end
`endif

  assign io_mem_req_bits_data = T0;
  assign T0 = r_valid_0 ? io_requestor_0_req_bits_data : T1;
  assign T1 = r_valid_1 ? io_requestor_1_req_bits_data : io_requestor_2_req_bits_data;
  assign io_mem_req_bits_cmd = T2;
  assign T2 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : T3;
  assign T3 = io_requestor_1_req_valid ? io_requestor_1_req_bits_cmd : io_requestor_2_req_bits_cmd;
  assign io_mem_req_bits_tag = T53;
  assign T53 = T4[4'h8:1'h0];
  assign T4 = io_requestor_0_req_valid ? T8 : T5;
  assign T5 = io_requestor_1_req_valid ? T7 : T6;
  assign T6 = {io_requestor_2_req_bits_tag, 2'h2};
  assign T7 = {io_requestor_1_req_bits_tag, 2'h1};
  assign T8 = {io_requestor_0_req_bits_tag, 2'h0};
  assign io_mem_req_bits_addr = T9;
  assign T9 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : T10;
  assign T10 = io_requestor_1_req_valid ? io_requestor_1_req_bits_addr : io_requestor_2_req_bits_addr;
  assign io_mem_req_bits_phys = T11;
  assign T11 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : T12;
  assign T12 = io_requestor_1_req_valid ? io_requestor_1_req_bits_phys : io_requestor_2_req_bits_phys;
  assign io_mem_req_bits_typ = T13;
  assign T13 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : T14;
  assign T14 = io_requestor_1_req_valid ? io_requestor_1_req_bits_typ : io_requestor_2_req_bits_typ;
  assign io_mem_req_bits_kill = T15;
  assign T15 = r_valid_0 ? io_requestor_0_req_bits_kill : T16;
  assign T16 = r_valid_1 ? io_requestor_1_req_bits_kill : io_requestor_2_req_bits_kill;
  assign io_mem_req_valid = T17;
  assign T17 = T18 | io_requestor_2_req_valid;
  assign T18 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T54;
  assign T54 = {2'h0, T19};
  assign T19 = io_mem_replay_next_bits >> 2'h2;
  assign io_requestor_0_replay_next_valid = T20;
  assign T20 = io_mem_replay_next_valid & T21;
  assign T21 = T22 == 2'h0;
  assign T22 = io_mem_replay_next_bits[1'h1:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T55;
  assign T55 = {2'h0, T23};
  assign T23 = io_mem_resp_bits_tag >> 2'h2;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_replay = T24;
  assign T24 = io_mem_resp_bits_replay & T25;
  assign T25 = T26 == 2'h0;
  assign T26 = io_mem_resp_bits_tag[1'h1:1'h0];
  assign io_requestor_0_resp_bits_nack = T27;
  assign T27 = io_mem_resp_bits_nack & T25;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_valid = T28;
  assign T28 = io_mem_resp_valid & T25;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T56;
  assign T56 = {2'h0, T29};
  assign T29 = io_mem_replay_next_bits >> 2'h2;
  assign io_requestor_1_replay_next_valid = T30;
  assign T30 = io_mem_replay_next_valid & T31;
  assign T31 = T32 == 2'h1;
  assign T32 = io_mem_replay_next_bits[1'h1:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T57;
  assign T57 = {2'h0, T33};
  assign T33 = io_mem_resp_bits_tag >> 2'h2;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_replay = T34;
  assign T34 = io_mem_resp_bits_replay & T35;
  assign T35 = T36 == 2'h1;
  assign T36 = io_mem_resp_bits_tag[1'h1:1'h0];
  assign io_requestor_1_resp_bits_nack = T37;
  assign T37 = io_mem_resp_bits_nack & T35;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_valid = T38;
  assign T38 = io_mem_resp_valid & T35;
  assign io_requestor_1_req_ready = T39;
  assign T39 = io_requestor_0_req_ready & T40;
  assign T40 = io_requestor_0_req_valid ^ 1'h1;
  assign io_requestor_2_ordered = io_mem_ordered;
  assign io_requestor_2_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_2_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_2_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_2_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_2_replay_next_bits = T58;
  assign T58 = {2'h0, T41};
  assign T41 = io_mem_replay_next_bits >> 2'h2;
  assign io_requestor_2_replay_next_valid = T42;
  assign T42 = io_mem_replay_next_valid & T43;
  assign T43 = T44 == 2'h2;
  assign T44 = io_mem_replay_next_bits[1'h1:1'h0];
  assign io_requestor_2_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_2_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_2_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_2_resp_bits_tag = T59;
  assign T59 = {2'h0, T45};
  assign T45 = io_mem_resp_bits_tag >> 2'h2;
  assign io_requestor_2_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_2_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_2_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_2_resp_bits_replay = T46;
  assign T46 = io_mem_resp_bits_replay & T47;
  assign T47 = T48 == 2'h2;
  assign T48 = io_mem_resp_bits_tag[1'h1:1'h0];
  assign io_requestor_2_resp_bits_nack = T49;
  assign T49 = io_mem_resp_bits_nack & T47;
  assign io_requestor_2_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_2_resp_valid = T50;
  assign T50 = io_mem_resp_valid & T47;
  assign io_requestor_2_req_ready = T51;
  assign T51 = io_requestor_1_req_ready & T52;
  assign T52 = io_requestor_1_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_1 <= io_requestor_1_req_valid;
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [511:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [511:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [511:0] io_in_0_bits_payload_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_a_type,
    output[511:0] io_out_bits_payload_subblock,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T81;
  wire[1:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire[511:0] T12;
  wire[511:0] T13;
  wire T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[511:0] T25;
  wire[511:0] T26;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire[25:0] T33;
  wire[25:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T10 ? 2'h1 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = io_in_0_valid ? 2'h0 : T4;
  assign T4 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T5 = io_in_2_valid & T6;
  assign T6 = R7 < 2'h2;
  assign T81 = reset ? 2'h0 : T8;
  assign T8 = T9 ? T0 : R7;
  assign T9 = io_out_ready & io_out_valid;
  assign T10 = io_in_1_valid & T11;
  assign T11 = R7 < 2'h1;
  assign io_out_bits_payload_subblock = T12;
  assign T12 = T16 ? io_in_2_bits_payload_subblock : T13;
  assign T13 = T14 ? io_in_1_bits_payload_subblock : io_in_0_bits_payload_subblock;
  assign T14 = T15[1'h0:1'h0];
  assign T15 = T0;
  assign T16 = T15[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T17;
  assign T17 = T20 ? io_in_2_bits_payload_a_type : T18;
  assign T18 = T19 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T19 = T15[1'h0:1'h0];
  assign T20 = T15[1'h1:1'h1];
  assign io_out_bits_payload_uncached = T21;
  assign T21 = T24 ? io_in_2_bits_payload_uncached : T22;
  assign T22 = T23 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T23 = T15[1'h0:1'h0];
  assign T24 = T15[1'h1:1'h1];
  assign io_out_bits_payload_data = T25;
  assign T25 = T28 ? io_in_2_bits_payload_data : T26;
  assign T26 = T27 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T27 = T15[1'h0:1'h0];
  assign T28 = T15[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T29;
  assign T29 = T32 ? io_in_2_bits_payload_client_xact_id : T30;
  assign T30 = T31 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T31 = T15[1'h0:1'h0];
  assign T32 = T15[1'h1:1'h1];
  assign io_out_bits_payload_addr = T33;
  assign T33 = T36 ? io_in_2_bits_payload_addr : T34;
  assign T34 = T35 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T35 = T15[1'h0:1'h0];
  assign T36 = T15[1'h1:1'h1];
  assign io_out_bits_header_dst = T37;
  assign T37 = T40 ? io_in_2_bits_header_dst : T38;
  assign T38 = T39 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T39 = T15[1'h0:1'h0];
  assign T40 = T15[1'h1:1'h1];
  assign io_out_bits_header_src = T41;
  assign T41 = T44 ? io_in_2_bits_header_src : T42;
  assign T42 = T43 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T43 = T15[1'h0:1'h0];
  assign T44 = T15[1'h1:1'h1];
  assign io_out_valid = T45;
  assign T45 = T48 ? io_in_2_valid : T46;
  assign T46 = T47 ? io_in_1_valid : io_in_0_valid;
  assign T47 = T15[1'h0:1'h0];
  assign T48 = T15[1'h1:1'h1];
  assign io_in_0_ready = T49;
  assign T49 = T50 & io_out_ready;
  assign T50 = T60 | T51;
  assign T51 = T52 ^ 1'h1;
  assign T52 = T55 | T53;
  assign T53 = io_in_2_valid & T54;
  assign T54 = R7 < 2'h2;
  assign T55 = T58 | T56;
  assign T56 = io_in_1_valid & T57;
  assign T57 = R7 < 2'h1;
  assign T58 = io_in_0_valid & T59;
  assign T59 = R7 < 2'h0;
  assign T60 = R7 < 2'h0;
  assign io_in_1_ready = T61;
  assign T61 = T62 & io_out_ready;
  assign T62 = T67 | T63;
  assign T63 = T64 ^ 1'h1;
  assign T64 = T65 | io_in_0_valid;
  assign T65 = T66 | T53;
  assign T66 = T58 | T56;
  assign T67 = T69 & T68;
  assign T68 = R7 < 2'h1;
  assign T69 = T58 ^ 1'h1;
  assign io_in_2_ready = T70;
  assign T70 = T71 & io_out_ready;
  assign T71 = T77 | T72;
  assign T72 = T73 ^ 1'h1;
  assign T73 = T74 | io_in_1_valid;
  assign T74 = T75 | io_in_0_valid;
  assign T75 = T76 | T53;
  assign T76 = T58 | T56;
  assign T77 = T79 & T78;
  assign T78 = R7 < 2'h2;
  assign T79 = T80 ^ 1'h1;
  assign T80 = T58 | T56;

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T9) begin
      R7 <= T0;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T61;
  wire[1:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T10 ? 2'h1 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = io_in_0_valid ? 2'h0 : T4;
  assign T4 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T5 = io_in_2_valid & T6;
  assign T6 = R7 < 2'h2;
  assign T61 = reset ? 2'h0 : T8;
  assign T8 = T9 ? T0 : R7;
  assign T9 = io_out_ready & io_out_valid;
  assign T10 = io_in_1_valid & T11;
  assign T11 = R7 < 2'h1;
  assign io_out_bits_payload_master_xact_id = T12;
  assign T12 = T16 ? io_in_2_bits_payload_master_xact_id : T13;
  assign T13 = T14 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T14 = T15[1'h0:1'h0];
  assign T15 = T0;
  assign T16 = T15[1'h1:1'h1];
  assign io_out_bits_header_dst = T17;
  assign T17 = T20 ? io_in_2_bits_header_dst : T18;
  assign T18 = T19 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T19 = T15[1'h0:1'h0];
  assign T20 = T15[1'h1:1'h1];
  assign io_out_bits_header_src = T21;
  assign T21 = T24 ? io_in_2_bits_header_src : T22;
  assign T22 = T23 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T23 = T15[1'h0:1'h0];
  assign T24 = T15[1'h1:1'h1];
  assign io_out_valid = T25;
  assign T25 = T28 ? io_in_2_valid : T26;
  assign T26 = T27 ? io_in_1_valid : io_in_0_valid;
  assign T27 = T15[1'h0:1'h0];
  assign T28 = T15[1'h1:1'h1];
  assign io_in_0_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = T40 | T31;
  assign T31 = T32 ^ 1'h1;
  assign T32 = T35 | T33;
  assign T33 = io_in_2_valid & T34;
  assign T34 = R7 < 2'h2;
  assign T35 = T38 | T36;
  assign T36 = io_in_1_valid & T37;
  assign T37 = R7 < 2'h1;
  assign T38 = io_in_0_valid & T39;
  assign T39 = R7 < 2'h0;
  assign T40 = R7 < 2'h0;
  assign io_in_1_ready = T41;
  assign T41 = T42 & io_out_ready;
  assign T42 = T47 | T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T45 | io_in_0_valid;
  assign T45 = T46 | T33;
  assign T46 = T38 | T36;
  assign T47 = T49 & T48;
  assign T48 = R7 < 2'h1;
  assign T49 = T38 ^ 1'h1;
  assign io_in_2_ready = T50;
  assign T50 = T51 & io_out_ready;
  assign T51 = T57 | T52;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T54 | io_in_1_valid;
  assign T54 = T55 | io_in_0_valid;
  assign T55 = T56 | T33;
  assign T56 = T38 | T36;
  assign T57 = T59 & T58;
  assign T58 = R7 < 2'h2;
  assign T59 = T60 ^ 1'h1;
  assign T60 = T38 | T36;

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T9) begin
      R7 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatAppendsArbiterId(input clk, input reset,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [2:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_2_acquire_bits_payload_data,
    input  io_in_2_acquire_bits_payload_uncached,
    input [1:0] io_in_2_acquire_bits_payload_a_type,
    input [511:0] io_in_2_acquire_bits_payload_subblock,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[511:0] io_in_2_grant_bits_payload_data,
    output[2:0] io_in_2_grant_bits_payload_client_xact_id,
    output[2:0] io_in_2_grant_bits_payload_master_xact_id,
    output io_in_2_grant_bits_payload_uncached,
    output[1:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input [2:0] io_in_2_finish_bits_payload_master_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [2:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input  io_in_1_acquire_bits_payload_uncached,
    input [1:0] io_in_1_acquire_bits_payload_a_type,
    input [511:0] io_in_1_acquire_bits_payload_subblock,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[2:0] io_in_1_grant_bits_payload_client_xact_id,
    output[2:0] io_in_1_grant_bits_payload_master_xact_id,
    output io_in_1_grant_bits_payload_uncached,
    output[1:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [2:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [2:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input  io_in_0_acquire_bits_payload_uncached,
    input [1:0] io_in_0_acquire_bits_payload_a_type,
    input [511:0] io_in_0_acquire_bits_payload_subblock,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[2:0] io_in_0_grant_bits_payload_client_xact_id,
    output[2:0] io_in_0_grant_bits_payload_master_xact_id,
    output io_in_0_grant_bits_payload_uncached,
    output[1:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [2:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[2:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output io_out_acquire_bits_payload_uncached,
    output[1:0] io_out_acquire_bits_payload_a_type,
    output[511:0] io_out_acquire_bits_payload_subblock,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [2:0] io_out_grant_bits_payload_client_xact_id,
    input [2:0] io_out_grant_bits_payload_master_xact_id,
    input  io_out_grant_bits_payload_uncached,
    input [1:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[2:0] io_out_finish_bits_payload_master_xact_id
);

  wire[2:0] T21;
  wire[4:0] T22;
  wire[2:0] T23;
  wire[4:0] T24;
  wire[2:0] T25;
  wire[4:0] T26;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[2:0] T18;
  wire T12;
  wire T13;
  wire[2:0] T19;
  wire T14;
  wire T15;
  wire[2:0] T20;
  wire T16;
  wire T17;
  wire RRArbiter_0_io_in_2_ready;
  wire RRArbiter_0_io_in_1_ready;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_0_io_out_valid;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[2:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire RRArbiter_0_io_out_bits_payload_uncached;
  wire[1:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] RRArbiter_0_io_out_bits_payload_subblock;
  wire RRArbiter_1_io_in_2_ready;
  wire RRArbiter_1_io_in_1_ready;
  wire RRArbiter_1_io_in_0_ready;
  wire RRArbiter_1_io_out_valid;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[2:0] RRArbiter_1_io_out_bits_payload_master_xact_id;


  assign T21 = T22[2'h2:1'h0];
  assign T22 = {io_in_0_acquire_bits_payload_client_xact_id, 2'h0};
  assign T23 = T24[2'h2:1'h0];
  assign T24 = {io_in_1_acquire_bits_payload_client_xact_id, 2'h1};
  assign T25 = T26[2'h2:1'h0];
  assign T26 = {io_in_2_acquire_bits_payload_client_xact_id, 2'h2};
  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T9 ? io_in_2_grant_ready : T1;
  assign T1 = T6 ? io_in_1_grant_ready : T2;
  assign T2 = T3 ? io_in_0_grant_ready : 1'h0;
  assign T3 = T4 == 2'h0;
  assign T4 = T5;
  assign T5 = io_out_grant_bits_payload_client_xact_id[1'h1:1'h0];
  assign T6 = T7 == 2'h1;
  assign T7 = T8;
  assign T8 = io_out_grant_bits_payload_client_xact_id[1'h1:1'h0];
  assign T9 = T10 == 2'h2;
  assign T10 = T11;
  assign T11 = io_out_grant_bits_payload_client_xact_id[1'h1:1'h0];
  assign io_out_acquire_bits_payload_subblock = RRArbiter_0_io_out_bits_payload_subblock;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_uncached = RRArbiter_0_io_out_bits_payload_uncached;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = T18;
  assign T18 = {2'h0, T12};
  assign T12 = io_out_grant_bits_payload_client_xact_id >> 2'h2;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T13;
  assign T13 = T3 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = T19;
  assign T19 = {2'h0, T14};
  assign T14 = io_out_grant_bits_payload_client_xact_id >> 2'h2;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T15;
  assign T15 = T6 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  assign io_in_2_finish_ready = RRArbiter_1_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_2_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = T20;
  assign T20 = {2'h0, T16};
  assign T16 = io_out_grant_bits_payload_client_xact_id >> 2'h2;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = RRArbiter_0_io_in_2_ready;
  RRArbiter_1 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( RRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( T25 ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_acquire_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_acquire_bits_payload_subblock ),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T23 ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_acquire_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_acquire_bits_payload_subblock ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T21 ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_acquire_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_acquire_bits_payload_subblock ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( RRArbiter_0_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( RRArbiter_0_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  RRArbiter_2 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( RRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_finish_bits_payload_master_xact_id ),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [8:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[8:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[63:0] io_deq_bits_data,
    output io_count
);

  wire T33;
  wire[1:0] T0;
  reg  full;
  wire T34;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_flow;
  wire empty;
  wire T3;
  wire T4;
  wire do_deq;
  wire T5;
  wire T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[126:0] T9;
  reg [126:0] ram [0:0];
  wire[126:0] T10;
  wire[126:0] T11;
  wire[126:0] T12;
  wire[121:0] T13;
  wire[68:0] T14;
  wire[52:0] T15;
  wire[4:0] T16;
  wire[3:0] T17;
  wire[4:0] T18;
  wire[4:0] T19;
  wire[8:0] T20;
  wire[8:0] T21;
  wire[43:0] T22;
  wire[43:0] T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T33;
  assign T33 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T34 = reset ? 1'h0 : T1;
  assign T1 = T4 ? do_enq : full;
  assign do_enq = T3 & T2;
  assign T2 = do_flow ^ 1'h1;
  assign do_flow = empty & io_deq_ready;
  assign empty = full ^ 1'h1;
  assign T3 = io_enq_ready & io_enq_valid;
  assign T4 = do_enq != do_deq;
  assign do_deq = T6 & T5;
  assign T5 = do_flow ^ 1'h1;
  assign T6 = io_deq_ready & io_deq_valid;
  assign io_deq_bits_data = T7;
  assign T7 = empty ? io_enq_bits_data : T8;
  assign T8 = T9[6'h3f:1'h0];
  assign T9 = ram[1'h0];
  assign T11 = T12;
  assign T12 = {T16, T13};
  assign T13 = {T15, T14};
  assign T14 = {io_enq_bits_cmd, io_enq_bits_data};
  assign T15 = {io_enq_bits_addr, io_enq_bits_tag};
  assign T16 = {io_enq_bits_kill, T17};
  assign T17 = {io_enq_bits_typ, io_enq_bits_phys};
  assign io_deq_bits_cmd = T18;
  assign T18 = empty ? io_enq_bits_cmd : T19;
  assign T19 = T9[7'h44:7'h40];
  assign io_deq_bits_tag = T20;
  assign T20 = empty ? io_enq_bits_tag : T21;
  assign T21 = T9[7'h4d:7'h45];
  assign io_deq_bits_addr = T22;
  assign T22 = empty ? io_enq_bits_addr : T23;
  assign T23 = T9[7'h79:7'h4e];
  assign io_deq_bits_phys = T24;
  assign T24 = empty ? io_enq_bits_phys : T25;
  assign T25 = T9[7'h7a:7'h7a];
  assign io_deq_bits_typ = T26;
  assign T26 = empty ? io_enq_bits_typ : T27;
  assign T27 = T9[7'h7d:7'h7b];
  assign io_deq_bits_kill = T28;
  assign T28 = empty ? io_enq_bits_kill : T29;
  assign T29 = T9[7'h7e:7'h7e];
  assign io_deq_valid = T30;
  assign T30 = T31 | io_enq_valid;
  assign T31 = empty ^ 1'h1;
  assign io_enq_ready = T32;
  assign T32 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T4) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T11;
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [8:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[8:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[63:0] io_deq_bits_data,
    output io_count
);

  wire T21;
  wire[1:0] T0;
  reg  full;
  wire T22;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[63:0] T3;
  wire[126:0] T4;
  reg [126:0] ram [0:0];
  wire[126:0] T5;
  wire[126:0] T6;
  wire[126:0] T7;
  wire[121:0] T8;
  wire[68:0] T9;
  wire[52:0] T10;
  wire[4:0] T11;
  wire[3:0] T12;
  wire[4:0] T13;
  wire[8:0] T14;
  wire[43:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire empty;
  wire T20;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T21;
  assign T21 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T22 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_data = T3;
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_cmd, io_enq_bits_data};
  assign T10 = {io_enq_bits_addr, io_enq_bits_tag};
  assign T11 = {io_enq_bits_kill, T12};
  assign T12 = {io_enq_bits_typ, io_enq_bits_phys};
  assign io_deq_bits_cmd = T13;
  assign T13 = T4[7'h44:7'h40];
  assign io_deq_bits_tag = T14;
  assign T14 = T4[7'h4d:7'h45];
  assign io_deq_bits_addr = T15;
  assign T15 = T4[7'h79:7'h4e];
  assign io_deq_bits_phys = T16;
  assign T16 = T4[7'h7a:7'h7a];
  assign io_deq_bits_typ = T17;
  assign T17 = T4[7'h7d:7'h7b];
  assign io_deq_bits_kill = T18;
  assign T18 = T4[7'h7e:7'h7e];
  assign io_deq_valid = T19;
  assign T19 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [8:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [8:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[2:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[8:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[63:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[8:0] T5;
  wire[43:0] T6;
  wire T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T2;
  assign T2 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T3 = T0;
  assign io_out_bits_cmd = T4;
  assign T4 = T3 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T5;
  assign T5 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T6;
  assign T6 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T7;
  assign T7 = T3 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T8;
  assign T8 = T3 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T9;
  assign T9 = T3 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T10;
  assign T10 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module SimpleHellaCacheIF(input clk, input reset,
    output io_requestor_req_ready,
    input  io_requestor_req_valid,
    input  io_requestor_req_bits_kill,
    input [2:0] io_requestor_req_bits_typ,
    input  io_requestor_req_bits_phys,
    input [43:0] io_requestor_req_bits_addr,
    input [8:0] io_requestor_req_bits_tag,
    input [4:0] io_requestor_req_bits_cmd,
    input [63:0] io_requestor_req_bits_data,
    output io_requestor_resp_valid,
    output[63:0] io_requestor_resp_bits_data,
    output io_requestor_resp_bits_nack,
    output io_requestor_resp_bits_replay,
    output[2:0] io_requestor_resp_bits_typ,
    output io_requestor_resp_bits_has_data,
    output[63:0] io_requestor_resp_bits_data_subword,
    output[8:0] io_requestor_resp_bits_tag,
    output[3:0] io_requestor_resp_bits_cmd,
    output[43:0] io_requestor_resp_bits_addr,
    output[63:0] io_requestor_resp_bits_store_data,
    //output io_requestor_replay_next_valid
    //output[8:0] io_requestor_replay_next_bits
    //output io_requestor_xcpt_ma_ld
    //output io_requestor_xcpt_ma_st
    //output io_requestor_xcpt_pf_ld
    //output io_requestor_xcpt_pf_st
    input  io_requestor_ptw_req_ready,
    //output io_requestor_ptw_req_valid
    //output[29:0] io_requestor_ptw_req_bits
    input  io_requestor_ptw_resp_valid,
    input  io_requestor_ptw_resp_bits_error,
    input [18:0] io_requestor_ptw_resp_bits_ppn,
    input [5:0] io_requestor_ptw_resp_bits_perm,
    input [7:0] io_requestor_ptw_status_ip,
    input [7:0] io_requestor_ptw_status_im,
    input [6:0] io_requestor_ptw_status_zero,
    input  io_requestor_ptw_status_er,
    input  io_requestor_ptw_status_vm,
    input  io_requestor_ptw_status_s64,
    input  io_requestor_ptw_status_u64,
    input  io_requestor_ptw_status_ef,
    input  io_requestor_ptw_status_pei,
    input  io_requestor_ptw_status_ei,
    input  io_requestor_ptw_status_ps,
    input  io_requestor_ptw_status_s,
    input  io_requestor_ptw_invalidate,
    input  io_requestor_ptw_sret,
    //output io_requestor_ordered
    input  io_cache_req_ready,
    output io_cache_req_valid,
    output io_cache_req_bits_kill,
    output[2:0] io_cache_req_bits_typ,
    output io_cache_req_bits_phys,
    output[43:0] io_cache_req_bits_addr,
    output[8:0] io_cache_req_bits_tag,
    output[4:0] io_cache_req_bits_cmd,
    output[63:0] io_cache_req_bits_data,
    input  io_cache_resp_valid,
    input [63:0] io_cache_resp_bits_data,
    input  io_cache_resp_bits_nack,
    input  io_cache_resp_bits_replay,
    input [2:0] io_cache_resp_bits_typ,
    input  io_cache_resp_bits_has_data,
    input [63:0] io_cache_resp_bits_data_subword,
    input [8:0] io_cache_resp_bits_tag,
    input [3:0] io_cache_resp_bits_cmd,
    input [43:0] io_cache_resp_bits_addr,
    input [63:0] io_cache_resp_bits_store_data,
    input  io_cache_replay_next_valid,
    input [8:0] io_cache_replay_next_bits,
    input  io_cache_xcpt_ma_ld,
    input  io_cache_xcpt_ma_st,
    input  io_cache_xcpt_pf_ld,
    input  io_cache_xcpt_pf_st,
    //output io_cache_ptw_req_ready
    //input  io_cache_ptw_req_valid
    //input [29:0] io_cache_ptw_req_bits
    //output io_cache_ptw_resp_valid
    //output io_cache_ptw_resp_bits_error
    //output[18:0] io_cache_ptw_resp_bits_ppn
    //output[5:0] io_cache_ptw_resp_bits_perm
    //output[7:0] io_cache_ptw_status_ip
    //output[7:0] io_cache_ptw_status_im
    //output[6:0] io_cache_ptw_status_zero
    //output io_cache_ptw_status_er
    //output io_cache_ptw_status_vm
    //output io_cache_ptw_status_s64
    //output io_cache_ptw_status_u64
    //output io_cache_ptw_status_ef
    //output io_cache_ptw_status_pei
    //output io_cache_ptw_status_ei
    //output io_cache_ptw_status_ps
    //output io_cache_ptw_status_s
    //output io_cache_ptw_invalidate
    //output io_cache_ptw_sret
    input  io_cache_ordered
);

  wire T14;
  wire T15;
  wire replaying_cmb;
  wire T4;
  wire T5;
  reg  replaying;
  wire T13;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg  R11;
  reg  R12;
  reg  s2_req_fire;
  reg  s1_req_fire;
  wire s0_req_fire;
  wire T16;
  wire[4:0] T17;
  wire T18;
  reg  s3_nack;
  wire[63:0] T19;
  wire[4:0] T20;
  wire[4:0] T21;
  wire[8:0] T22;
  wire[43:0] T23;
  wire[2:0] T24;
  wire T25;
  reg [63:0] R0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  wire replayq1_io_deq_valid;
  wire replayq1_io_deq_bits_kill;
  wire[2:0] replayq1_io_deq_bits_typ;
  wire replayq1_io_deq_bits_phys;
  wire[43:0] replayq1_io_deq_bits_addr;
  wire[8:0] replayq1_io_deq_bits_tag;
  wire[4:0] replayq1_io_deq_bits_cmd;
  wire[63:0] replayq1_io_deq_bits_data;
  wire replayq2_io_deq_valid;
  wire[2:0] replayq2_io_deq_bits_typ;
  wire[43:0] replayq2_io_deq_bits_addr;
  wire[8:0] replayq2_io_deq_bits_tag;
  wire[4:0] replayq2_io_deq_bits_cmd;
  wire[63:0] replayq2_io_deq_bits_data;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire[2:0] req_arb_io_out_bits_typ;
  wire[43:0] req_arb_io_out_bits_addr;
  wire[8:0] req_arb_io_out_bits_tag;
  wire[4:0] req_arb_io_out_bits_cmd;
  wire[63:0] req_arb_io_out_bits_data;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    replaying = {1{$random}};
    R11 = {1{$random}};
    R12 = {1{$random}};
    s2_req_fire = {1{$random}};
    s1_req_fire = {1{$random}};
    s3_nack = {1{$random}};
    R0 = {2{$random}};
  end
`endif

  assign T14 = T15 & io_requestor_req_valid;
  assign T15 = replaying_cmb ^ 1'h1;
  assign replaying_cmb = T4;
  assign T4 = T6 ? 1'h0 : T5;
  assign T5 = io_cache_resp_bits_nack ? 1'h1 : replaying;
  assign T13 = reset ? 1'h0 : replaying_cmb;
  assign T6 = T8 & T7;
  assign T7 = replayq2_io_deq_valid ^ 1'h1;
  assign T8 = T10 & T9;
  assign T9 = io_cache_resp_bits_nack ^ 1'h1;
  assign T10 = s2_req_fire & R11;
  assign s0_req_fire = io_cache_req_ready & io_cache_req_valid;
  assign T16 = T8 & replayq2_io_deq_valid;
  assign T17 = {1'h0, io_cache_resp_bits_cmd};
  assign T18 = s2_req_fire & s3_nack;
  assign T19 = T16 ? replayq2_io_deq_bits_data : io_cache_resp_bits_store_data;
  assign T20 = T16 ? replayq2_io_deq_bits_cmd : T21;
  assign T21 = {1'h0, io_cache_resp_bits_cmd};
  assign T22 = T16 ? replayq2_io_deq_bits_tag : io_cache_resp_bits_tag;
  assign T23 = T16 ? replayq2_io_deq_bits_addr : io_cache_resp_bits_addr;
  assign T24 = T16 ? replayq2_io_deq_bits_typ : io_cache_resp_bits_typ;
  assign T25 = T16 ? 1'h1 : io_cache_resp_bits_nack;
  assign io_cache_req_bits_data = R0;
  assign T1 = s0_req_fire ? req_arb_io_out_bits_data : R0;
  assign io_cache_req_bits_cmd = req_arb_io_out_bits_cmd;
  assign io_cache_req_bits_tag = req_arb_io_out_bits_tag;
  assign io_cache_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_cache_req_bits_phys = 1'h1;
  assign io_cache_req_bits_typ = req_arb_io_out_bits_typ;
  assign io_cache_req_bits_kill = io_cache_resp_bits_nack;
  assign io_cache_req_valid = req_arb_io_out_valid;
  assign io_requestor_resp_bits_store_data = io_cache_resp_bits_store_data;
  assign io_requestor_resp_bits_addr = io_cache_resp_bits_addr;
  assign io_requestor_resp_bits_cmd = io_cache_resp_bits_cmd;
  assign io_requestor_resp_bits_tag = io_cache_resp_bits_tag;
  assign io_requestor_resp_bits_data_subword = io_cache_resp_bits_data_subword;
  assign io_requestor_resp_bits_has_data = io_cache_resp_bits_has_data;
  assign io_requestor_resp_bits_typ = io_cache_resp_bits_typ;
  assign io_requestor_resp_bits_replay = io_cache_resp_bits_replay;
  assign io_requestor_resp_bits_nack = io_cache_resp_bits_nack;
  assign io_requestor_resp_bits_data = io_cache_resp_bits_data;
  assign io_requestor_resp_valid = io_cache_resp_valid;
  assign io_requestor_req_ready = T2;
  assign T2 = T3 & req_arb_io_in_1_ready;
  assign T3 = replaying_cmb ^ 1'h1;
  Queue_11 replayq1(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( T25 ),
       //.io_enq_bits_kill(  )
       .io_enq_bits_typ( T24 ),
       //.io_enq_bits_phys(  )
       .io_enq_bits_addr( T23 ),
       .io_enq_bits_tag( T22 ),
       .io_enq_bits_cmd( T20 ),
       .io_enq_bits_data( T19 ),
       .io_deq_ready( req_arb_io_in_0_ready ),
       .io_deq_valid( replayq1_io_deq_valid ),
       .io_deq_bits_kill( replayq1_io_deq_bits_kill ),
       .io_deq_bits_typ( replayq1_io_deq_bits_typ ),
       .io_deq_bits_phys( replayq1_io_deq_bits_phys ),
       .io_deq_bits_addr( replayq1_io_deq_bits_addr ),
       .io_deq_bits_tag( replayq1_io_deq_bits_tag ),
       .io_deq_bits_cmd( replayq1_io_deq_bits_cmd ),
       .io_deq_bits_data( replayq1_io_deq_bits_data )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign replayq1.io_enq_bits_kill = {1{$random}};
    assign replayq1.io_enq_bits_phys = {1{$random}};
  `endif
  Queue_12 replayq2(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( T18 ),
       //.io_enq_bits_kill(  )
       .io_enq_bits_typ( io_cache_resp_bits_typ ),
       //.io_enq_bits_phys(  )
       .io_enq_bits_addr( io_cache_resp_bits_addr ),
       .io_enq_bits_tag( io_cache_resp_bits_tag ),
       .io_enq_bits_cmd( T17 ),
       .io_enq_bits_data( io_cache_resp_bits_store_data ),
       .io_deq_ready( T16 ),
       .io_deq_valid( replayq2_io_deq_valid ),
       //.io_deq_bits_kill(  )
       .io_deq_bits_typ( replayq2_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( replayq2_io_deq_bits_addr ),
       .io_deq_bits_tag( replayq2_io_deq_bits_tag ),
       .io_deq_bits_cmd( replayq2_io_deq_bits_cmd ),
       .io_deq_bits_data( replayq2_io_deq_bits_data )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign replayq2.io_enq_bits_kill = {1{$random}};
    assign replayq2.io_enq_bits_phys = {1{$random}};
  `endif
  Arbiter_6 req_arb(
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_kill( io_requestor_req_bits_kill ),
       .io_in_1_bits_typ( io_requestor_req_bits_typ ),
       .io_in_1_bits_phys( io_requestor_req_bits_phys ),
       .io_in_1_bits_addr( io_requestor_req_bits_addr ),
       .io_in_1_bits_tag( io_requestor_req_bits_tag ),
       .io_in_1_bits_cmd( io_requestor_req_bits_cmd ),
       .io_in_1_bits_data( io_requestor_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( replayq1_io_deq_valid ),
       .io_in_0_bits_kill( replayq1_io_deq_bits_kill ),
       .io_in_0_bits_typ( replayq1_io_deq_bits_typ ),
       .io_in_0_bits_phys( replayq1_io_deq_bits_phys ),
       .io_in_0_bits_addr( replayq1_io_deq_bits_addr ),
       .io_in_0_bits_tag( replayq1_io_deq_bits_tag ),
       .io_in_0_bits_cmd( replayq1_io_deq_bits_cmd ),
       .io_in_0_bits_data( replayq1_io_deq_bits_data ),
       .io_out_ready( io_cache_req_ready ),
       .io_out_valid( req_arb_io_out_valid ),
       //.io_out_bits_kill(  )
       .io_out_bits_typ( req_arb_io_out_bits_typ ),
       //.io_out_bits_phys(  )
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_tag( req_arb_io_out_bits_tag ),
       .io_out_bits_cmd( req_arb_io_out_bits_cmd ),
       .io_out_bits_data( req_arb_io_out_bits_data )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      replaying <= 1'h0;
    end else begin
      replaying <= replaying_cmb;
    end
    R11 <= R12;
    R12 <= replaying_cmb;
    s2_req_fire <= s1_req_fire;
    s1_req_fire <= s0_req_fire;
    s3_nack <= io_cache_resp_bits_nack;
    if(s0_req_fire) begin
      R0 <= req_arb_io_out_bits_data;
    end
  end
endmodule

module RocketTile(input clk, input reset,
    input  io_tilelink_acquire_ready,
    output io_tilelink_acquire_valid,
    output[1:0] io_tilelink_acquire_bits_header_src,
    output[1:0] io_tilelink_acquire_bits_header_dst,
    output[25:0] io_tilelink_acquire_bits_payload_addr,
    output[2:0] io_tilelink_acquire_bits_payload_client_xact_id,
    output[511:0] io_tilelink_acquire_bits_payload_data,
    output io_tilelink_acquire_bits_payload_uncached,
    output[1:0] io_tilelink_acquire_bits_payload_a_type,
    output[511:0] io_tilelink_acquire_bits_payload_subblock,
    output io_tilelink_grant_ready,
    input  io_tilelink_grant_valid,
    input [1:0] io_tilelink_grant_bits_header_src,
    input [1:0] io_tilelink_grant_bits_header_dst,
    input [511:0] io_tilelink_grant_bits_payload_data,
    input [2:0] io_tilelink_grant_bits_payload_client_xact_id,
    input [2:0] io_tilelink_grant_bits_payload_master_xact_id,
    input  io_tilelink_grant_bits_payload_uncached,
    input [1:0] io_tilelink_grant_bits_payload_g_type,
    input  io_tilelink_finish_ready,
    output io_tilelink_finish_valid,
    output[1:0] io_tilelink_finish_bits_header_src,
    output[1:0] io_tilelink_finish_bits_header_dst,
    output[2:0] io_tilelink_finish_bits_payload_master_xact_id,
    output io_tilelink_probe_ready,
    input  io_tilelink_probe_valid,
    input [1:0] io_tilelink_probe_bits_header_src,
    input [1:0] io_tilelink_probe_bits_header_dst,
    input [25:0] io_tilelink_probe_bits_payload_addr,
    input [1:0] io_tilelink_probe_bits_payload_p_type,
    input  io_tilelink_release_ready,
    output io_tilelink_release_valid,
    output[1:0] io_tilelink_release_bits_header_src,
    output[1:0] io_tilelink_release_bits_header_dst,
    output[25:0] io_tilelink_release_bits_payload_addr,
    output[2:0] io_tilelink_release_bits_payload_client_xact_id,
    output[511:0] io_tilelink_release_bits_payload_data,
    output[2:0] io_tilelink_release_bits_payload_r_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready,
    output io_temac_sfp_tx_disable,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    output io_rocc_resp_ready,
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    output io_rocc_mem_req_ready,
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    output io_rocc_mem_resp_valid,
    output[63:0] io_rocc_mem_resp_bits_data,
    output io_rocc_mem_resp_bits_nack,
    output io_rocc_mem_resp_bits_replay,
    output[2:0] io_rocc_mem_resp_bits_typ,
    output io_rocc_mem_resp_bits_has_data,
    output[63:0] io_rocc_mem_resp_bits_data_subword,
    output[8:0] io_rocc_mem_resp_bits_tag,
    output[3:0] io_rocc_mem_resp_bits_cmd,
    output[43:0] io_rocc_mem_resp_bits_addr,
    output[63:0] io_rocc_mem_resp_bits_store_data,
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    output io_rocc_imem_acquire_ready,
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [2:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [511:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    output io_rocc_imem_grant_valid,
    output[1:0] io_rocc_imem_grant_bits_header_src,
    output[1:0] io_rocc_imem_grant_bits_header_dst,
    output[511:0] io_rocc_imem_grant_bits_payload_data,
    output[2:0] io_rocc_imem_grant_bits_payload_client_xact_id,
    output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id,
    output io_rocc_imem_grant_bits_payload_uncached,
    output[1:0] io_rocc_imem_grant_bits_payload_g_type,
    output io_rocc_imem_finish_ready,
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    output io_rocc_iptw_req_ready,
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    output io_rocc_iptw_resp_valid,
    output io_rocc_iptw_resp_bits_error,
    output[18:0] io_rocc_iptw_resp_bits_ppn,
    output[5:0] io_rocc_iptw_resp_bits_perm,
    output[7:0] io_rocc_iptw_status_ip,
    output[7:0] io_rocc_iptw_status_im,
    output[6:0] io_rocc_iptw_status_zero,
    output io_rocc_iptw_status_er,
    output io_rocc_iptw_status_vm,
    output io_rocc_iptw_status_s64,
    output io_rocc_iptw_status_u64,
    output io_rocc_iptw_status_ef,
    output io_rocc_iptw_status_pei,
    output io_rocc_iptw_status_ei,
    output io_rocc_iptw_status_ps,
    output io_rocc_iptw_status_s,
    output io_rocc_iptw_invalidate,
    output io_rocc_iptw_sret,
    output io_rocc_dptw_req_ready,
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    output io_rocc_dptw_resp_valid,
    output io_rocc_dptw_resp_bits_error,
    output[18:0] io_rocc_dptw_resp_bits_ppn,
    output[5:0] io_rocc_dptw_resp_bits_perm,
    output[7:0] io_rocc_dptw_status_ip,
    output[7:0] io_rocc_dptw_status_im,
    output[6:0] io_rocc_dptw_status_zero,
    output io_rocc_dptw_status_er,
    output io_rocc_dptw_status_vm,
    output io_rocc_dptw_status_s64,
    output io_rocc_dptw_status_u64,
    output io_rocc_dptw_status_ef,
    output io_rocc_dptw_status_pei,
    output io_rocc_dptw_status_ei,
    output io_rocc_dptw_status_ps,
    output io_rocc_dptw_status_s,
    output io_rocc_dptw_invalidate,
    output io_rocc_dptw_sret,
    output io_rocc_pptw_req_ready,
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    output io_rocc_pptw_resp_valid,
    output io_rocc_pptw_resp_bits_error,
    output[18:0] io_rocc_pptw_resp_bits_ppn,
    output[5:0] io_rocc_pptw_resp_bits_perm,
    output[7:0] io_rocc_pptw_status_ip,
    output[7:0] io_rocc_pptw_status_im,
    output[6:0] io_rocc_pptw_status_zero,
    output io_rocc_pptw_status_er,
    output io_rocc_pptw_status_vm,
    output io_rocc_pptw_status_s64,
    output io_rocc_pptw_status_u64,
    output io_rocc_pptw_status_ef,
    output io_rocc_pptw_status_pei,
    output io_rocc_pptw_status_ei,
    output io_rocc_pptw_status_ps,
    output io_rocc_pptw_status_s,
    output io_rocc_pptw_invalidate,
    output io_rocc_pptw_sret,
    output io_rocc_exception
);

  wire[2:0] T1;
  wire[4:0] T0;
  wire dcArb_io_requestor_2_req_ready;
  wire dcArb_io_requestor_2_resp_valid;
  wire[63:0] dcArb_io_requestor_2_resp_bits_data;
  wire dcArb_io_requestor_2_resp_bits_nack;
  wire dcArb_io_requestor_2_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_2_resp_bits_typ;
  wire dcArb_io_requestor_2_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_2_resp_bits_data_subword;
  wire[8:0] dcArb_io_requestor_2_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_2_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_2_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_2_resp_bits_store_data;
  wire dcArb_io_requestor_2_replay_next_valid;
  wire[8:0] dcArb_io_requestor_2_replay_next_bits;
  wire dcArb_io_requestor_2_xcpt_ma_ld;
  wire dcArb_io_requestor_2_xcpt_ma_st;
  wire dcArb_io_requestor_2_xcpt_pf_ld;
  wire dcArb_io_requestor_2_xcpt_pf_st;
  wire dcArb_io_requestor_2_ordered;
  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_subword;
  wire[8:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[8:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_subword;
  wire[8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[8:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire dcArb_io_mem_req_bits_kill;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_phys;
  wire[43:0] dcArb_io_mem_req_bits_addr;
  wire[8:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire ptw_io_requestor_4_req_ready;
  wire ptw_io_requestor_4_resp_valid;
  wire ptw_io_requestor_4_resp_bits_error;
  wire[18:0] ptw_io_requestor_4_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_4_resp_bits_perm;
  wire[7:0] ptw_io_requestor_4_status_ip;
  wire[7:0] ptw_io_requestor_4_status_im;
  wire[6:0] ptw_io_requestor_4_status_zero;
  wire ptw_io_requestor_4_status_er;
  wire ptw_io_requestor_4_status_vm;
  wire ptw_io_requestor_4_status_s64;
  wire ptw_io_requestor_4_status_u64;
  wire ptw_io_requestor_4_status_ef;
  wire ptw_io_requestor_4_status_pei;
  wire ptw_io_requestor_4_status_ei;
  wire ptw_io_requestor_4_status_ps;
  wire ptw_io_requestor_4_status_s;
  wire ptw_io_requestor_4_invalidate;
  wire ptw_io_requestor_4_sret;
  wire ptw_io_requestor_3_req_ready;
  wire ptw_io_requestor_3_resp_valid;
  wire ptw_io_requestor_3_resp_bits_error;
  wire[18:0] ptw_io_requestor_3_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_3_resp_bits_perm;
  wire[7:0] ptw_io_requestor_3_status_ip;
  wire[7:0] ptw_io_requestor_3_status_im;
  wire[6:0] ptw_io_requestor_3_status_zero;
  wire ptw_io_requestor_3_status_er;
  wire ptw_io_requestor_3_status_vm;
  wire ptw_io_requestor_3_status_s64;
  wire ptw_io_requestor_3_status_u64;
  wire ptw_io_requestor_3_status_ef;
  wire ptw_io_requestor_3_status_pei;
  wire ptw_io_requestor_3_status_ei;
  wire ptw_io_requestor_3_status_ps;
  wire ptw_io_requestor_3_status_s;
  wire ptw_io_requestor_3_invalidate;
  wire ptw_io_requestor_3_sret;
  wire ptw_io_requestor_2_req_ready;
  wire ptw_io_requestor_2_resp_valid;
  wire ptw_io_requestor_2_resp_bits_error;
  wire[18:0] ptw_io_requestor_2_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_2_resp_bits_perm;
  wire[7:0] ptw_io_requestor_2_status_ip;
  wire[7:0] ptw_io_requestor_2_status_im;
  wire[6:0] ptw_io_requestor_2_status_zero;
  wire ptw_io_requestor_2_status_er;
  wire ptw_io_requestor_2_status_vm;
  wire ptw_io_requestor_2_status_s64;
  wire ptw_io_requestor_2_status_u64;
  wire ptw_io_requestor_2_status_ef;
  wire ptw_io_requestor_2_status_pei;
  wire ptw_io_requestor_2_status_ei;
  wire ptw_io_requestor_2_status_ps;
  wire ptw_io_requestor_2_status_s;
  wire ptw_io_requestor_2_invalidate;
  wire ptw_io_requestor_2_sret;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[18:0] ptw_io_requestor_1_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_1_resp_bits_perm;
  wire[7:0] ptw_io_requestor_1_status_ip;
  wire[7:0] ptw_io_requestor_1_status_im;
  wire[6:0] ptw_io_requestor_1_status_zero;
  wire ptw_io_requestor_1_status_er;
  wire ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_s64;
  wire ptw_io_requestor_1_status_u64;
  wire ptw_io_requestor_1_status_ef;
  wire ptw_io_requestor_1_status_pei;
  wire ptw_io_requestor_1_status_ei;
  wire ptw_io_requestor_1_status_ps;
  wire ptw_io_requestor_1_status_s;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_1_sret;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[18:0] ptw_io_requestor_0_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_0_resp_bits_perm;
  wire[7:0] ptw_io_requestor_0_status_ip;
  wire[7:0] ptw_io_requestor_0_status_im;
  wire[6:0] ptw_io_requestor_0_status_zero;
  wire ptw_io_requestor_0_status_er;
  wire ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_s64;
  wire ptw_io_requestor_0_status_u64;
  wire ptw_io_requestor_0_status_ef;
  wire ptw_io_requestor_0_status_pei;
  wire ptw_io_requestor_0_status_ei;
  wire ptw_io_requestor_0_status_ps;
  wire ptw_io_requestor_0_status_s;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_requestor_0_sret;
  wire ptw_io_mem_req_valid;
  wire ptw_io_mem_req_bits_kill;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_phys;
  wire[43:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire memArb_io_in_2_acquire_ready;
  wire memArb_io_in_2_grant_valid;
  wire[1:0] memArb_io_in_2_grant_bits_header_src;
  wire[1:0] memArb_io_in_2_grant_bits_header_dst;
  wire[511:0] memArb_io_in_2_grant_bits_payload_data;
  wire[2:0] memArb_io_in_2_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_2_grant_bits_payload_master_xact_id;
  wire memArb_io_in_2_grant_bits_payload_uncached;
  wire[1:0] memArb_io_in_2_grant_bits_payload_g_type;
  wire memArb_io_in_2_finish_ready;
  wire memArb_io_in_1_acquire_ready;
  wire memArb_io_in_1_grant_valid;
  wire[1:0] memArb_io_in_1_grant_bits_header_src;
  wire[1:0] memArb_io_in_1_grant_bits_header_dst;
  wire[511:0] memArb_io_in_1_grant_bits_payload_data;
  wire[2:0] memArb_io_in_1_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_1_grant_bits_payload_master_xact_id;
  wire memArb_io_in_1_grant_bits_payload_uncached;
  wire[1:0] memArb_io_in_1_grant_bits_payload_g_type;
  wire memArb_io_in_1_finish_ready;
  wire memArb_io_in_0_acquire_ready;
  wire memArb_io_in_0_grant_valid;
  wire[1:0] memArb_io_in_0_grant_bits_header_src;
  wire[1:0] memArb_io_in_0_grant_bits_header_dst;
  wire[511:0] memArb_io_in_0_grant_bits_payload_data;
  wire[2:0] memArb_io_in_0_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_0_grant_bits_payload_master_xact_id;
  wire memArb_io_in_0_grant_bits_payload_uncached;
  wire[1:0] memArb_io_in_0_grant_bits_payload_g_type;
  wire memArb_io_in_0_finish_ready;
  wire memArb_io_out_acquire_valid;
  wire[1:0] memArb_io_out_acquire_bits_header_src;
  wire[1:0] memArb_io_out_acquire_bits_header_dst;
  wire[25:0] memArb_io_out_acquire_bits_payload_addr;
  wire[2:0] memArb_io_out_acquire_bits_payload_client_xact_id;
  wire[511:0] memArb_io_out_acquire_bits_payload_data;
  wire memArb_io_out_acquire_bits_payload_uncached;
  wire[1:0] memArb_io_out_acquire_bits_payload_a_type;
  wire[511:0] memArb_io_out_acquire_bits_payload_subblock;
  wire memArb_io_out_grant_ready;
  wire memArb_io_out_finish_valid;
  wire[1:0] memArb_io_out_finish_bits_header_src;
  wire[1:0] memArb_io_out_finish_bits_header_dst;
  wire[2:0] memArb_io_out_finish_bits_payload_master_xact_id;
  wire SimpleHellaCacheIF_io_requestor_req_ready;
  wire SimpleHellaCacheIF_io_requestor_resp_valid;
  wire[63:0] SimpleHellaCacheIF_io_requestor_resp_bits_data;
  wire SimpleHellaCacheIF_io_requestor_resp_bits_nack;
  wire SimpleHellaCacheIF_io_requestor_resp_bits_replay;
  wire[2:0] SimpleHellaCacheIF_io_requestor_resp_bits_typ;
  wire SimpleHellaCacheIF_io_requestor_resp_bits_has_data;
  wire[63:0] SimpleHellaCacheIF_io_requestor_resp_bits_data_subword;
  wire[8:0] SimpleHellaCacheIF_io_requestor_resp_bits_tag;
  wire[3:0] SimpleHellaCacheIF_io_requestor_resp_bits_cmd;
  wire[43:0] SimpleHellaCacheIF_io_requestor_resp_bits_addr;
  wire[63:0] SimpleHellaCacheIF_io_requestor_resp_bits_store_data;
  wire SimpleHellaCacheIF_io_cache_req_valid;
  wire SimpleHellaCacheIF_io_cache_req_bits_kill;
  wire[2:0] SimpleHellaCacheIF_io_cache_req_bits_typ;
  wire SimpleHellaCacheIF_io_cache_req_bits_phys;
  wire[43:0] SimpleHellaCacheIF_io_cache_req_bits_addr;
  wire[8:0] SimpleHellaCacheIF_io_cache_req_bits_tag;
  wire[4:0] SimpleHellaCacheIF_io_cache_req_bits_cmd;
  wire[63:0] SimpleHellaCacheIF_io_cache_req_bits_data;
  wire icache_io_cpu_resp_valid;
  wire[43:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data;
  wire icache_io_cpu_resp_bits_xcpt_ma;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire[42:0] icache_io_cpu_btb_resp_bits_target;
  wire[5:0] icache_io_cpu_btb_resp_bits_entry;
  wire[6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire icache_io_cpu_ptw_req_valid;
  wire[29:0] icache_io_cpu_ptw_req_bits;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[2:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire icache_io_mem_acquire_bits_payload_uncached;
  wire[1:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] icache_io_mem_acquire_bits_payload_subblock;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[8:0] dcache_io_cpu_resp_bits_tag;
  wire[3:0] dcache_io_cpu_resp_bits_cmd;
  wire[43:0] dcache_io_cpu_resp_bits_addr;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[8:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ptw_req_valid;
  wire[29:0] dcache_io_cpu_ptw_req_bits;
  wire dcache_io_cpu_ordered;
  wire dcache_io_mem_acquire_valid;
  wire[1:0] dcache_io_mem_acquire_bits_header_src;
  wire[1:0] dcache_io_mem_acquire_bits_header_dst;
  wire[25:0] dcache_io_mem_acquire_bits_payload_addr;
  wire[2:0] dcache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] dcache_io_mem_acquire_bits_payload_data;
  wire dcache_io_mem_acquire_bits_payload_uncached;
  wire[1:0] dcache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] dcache_io_mem_acquire_bits_payload_subblock;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_finish_valid;
  wire[1:0] dcache_io_mem_finish_bits_header_src;
  wire[1:0] dcache_io_mem_finish_bits_header_dst;
  wire[2:0] dcache_io_mem_finish_bits_payload_master_xact_id;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_header_src;
  wire[1:0] dcache_io_mem_release_bits_header_dst;
  wire[25:0] dcache_io_mem_release_bits_payload_addr;
  wire[2:0] dcache_io_mem_release_bits_payload_client_xact_id;
  wire[511:0] dcache_io_mem_release_bits_payload_data;
  wire[2:0] dcache_io_mem_release_bits_payload_r_type;
  wire core_io_host_pcr_req_ready;
  wire core_io_host_pcr_rep_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_pcr;
  wire core_io_imem_req_valid;
  wire[43:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire[42:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[42:0] core_io_imem_btb_update_bits_pc;
  wire[42:0] core_io_imem_btb_update_bits_target;
  wire[42:0] core_io_imem_btb_update_bits_returnAddr;
  wire core_io_imem_btb_update_bits_taken;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isCall;
  wire core_io_imem_btb_update_bits_isReturn;
  wire core_io_imem_btb_update_bits_mispredict;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire core_io_dmem_req_bits_kill;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_phys;
  wire[43:0] core_io_dmem_req_bits_addr;
  wire[8:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[63:0] core_io_dmem_req_bits_data;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_sret;
  wire[7:0] core_io_ptw_status_ip;
  wire[7:0] core_io_ptw_status_im;
  wire[6:0] core_io_ptw_status_zero;
  wire core_io_ptw_status_er;
  wire core_io_ptw_status_vm;
  wire core_io_ptw_status_s64;
  wire core_io_ptw_status_u64;
  wire core_io_ptw_status_ef;
  wire core_io_ptw_status_pei;
  wire core_io_ptw_status_ei;
  wire core_io_ptw_status_ps;
  wire core_io_ptw_status_s;
  wire core_io_rocc_cmd_valid;
  wire[6:0] core_io_rocc_cmd_bits_inst_funct;
  wire[4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire core_io_rocc_cmd_bits_inst_xd;
  wire core_io_rocc_cmd_bits_inst_xs1;
  wire core_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] core_io_rocc_cmd_bits_inst_rd;
  wire[6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] core_io_rocc_cmd_bits_rs1;
  wire[63:0] core_io_rocc_cmd_bits_rs2;
  wire core_io_rocc_resp_ready;
  wire core_io_rocc_s;
  wire core_io_rocc_exception;
  wire core_io_temac_rx_axis_fifo_tready;
  wire[7:0] core_io_temac_tx_axis_fifo_tdata;
  wire core_io_temac_tx_axis_fifo_tvalid;
  wire core_io_temac_tx_axis_fifo_tlast;
  wire[11:0] core_io_temac_s_axi_awaddr;
  wire core_io_temac_s_axi_awvalid;
  wire[31:0] core_io_temac_s_axi_wdata;
  wire core_io_temac_s_axi_wvalid;
  wire core_io_temac_s_axi_bready;
  wire[11:0] core_io_temac_s_axi_araddr;
  wire core_io_temac_s_axi_arvalid;
  wire core_io_temac_s_axi_rready;
  wire core_io_temac_sfp_tx_disable;


  assign io_rocc_exception = core_io_rocc_exception;
  assign io_rocc_pptw_sret = ptw_io_requestor_4_sret;
  assign io_rocc_pptw_invalidate = ptw_io_requestor_4_invalidate;
  assign io_rocc_pptw_status_s = ptw_io_requestor_4_status_s;
  assign io_rocc_pptw_status_ps = ptw_io_requestor_4_status_ps;
  assign io_rocc_pptw_status_ei = ptw_io_requestor_4_status_ei;
  assign io_rocc_pptw_status_pei = ptw_io_requestor_4_status_pei;
  assign io_rocc_pptw_status_ef = ptw_io_requestor_4_status_ef;
  assign io_rocc_pptw_status_u64 = ptw_io_requestor_4_status_u64;
  assign io_rocc_pptw_status_s64 = ptw_io_requestor_4_status_s64;
  assign io_rocc_pptw_status_vm = ptw_io_requestor_4_status_vm;
  assign io_rocc_pptw_status_er = ptw_io_requestor_4_status_er;
  assign io_rocc_pptw_status_zero = ptw_io_requestor_4_status_zero;
  assign io_rocc_pptw_status_im = ptw_io_requestor_4_status_im;
  assign io_rocc_pptw_status_ip = ptw_io_requestor_4_status_ip;
  assign io_rocc_pptw_resp_bits_perm = ptw_io_requestor_4_resp_bits_perm;
  assign io_rocc_pptw_resp_bits_ppn = ptw_io_requestor_4_resp_bits_ppn;
  assign io_rocc_pptw_resp_bits_error = ptw_io_requestor_4_resp_bits_error;
  assign io_rocc_pptw_resp_valid = ptw_io_requestor_4_resp_valid;
  assign io_rocc_pptw_req_ready = ptw_io_requestor_4_req_ready;
  assign io_rocc_dptw_sret = ptw_io_requestor_3_sret;
  assign io_rocc_dptw_invalidate = ptw_io_requestor_3_invalidate;
  assign io_rocc_dptw_status_s = ptw_io_requestor_3_status_s;
  assign io_rocc_dptw_status_ps = ptw_io_requestor_3_status_ps;
  assign io_rocc_dptw_status_ei = ptw_io_requestor_3_status_ei;
  assign io_rocc_dptw_status_pei = ptw_io_requestor_3_status_pei;
  assign io_rocc_dptw_status_ef = ptw_io_requestor_3_status_ef;
  assign io_rocc_dptw_status_u64 = ptw_io_requestor_3_status_u64;
  assign io_rocc_dptw_status_s64 = ptw_io_requestor_3_status_s64;
  assign io_rocc_dptw_status_vm = ptw_io_requestor_3_status_vm;
  assign io_rocc_dptw_status_er = ptw_io_requestor_3_status_er;
  assign io_rocc_dptw_status_zero = ptw_io_requestor_3_status_zero;
  assign io_rocc_dptw_status_im = ptw_io_requestor_3_status_im;
  assign io_rocc_dptw_status_ip = ptw_io_requestor_3_status_ip;
  assign io_rocc_dptw_resp_bits_perm = ptw_io_requestor_3_resp_bits_perm;
  assign io_rocc_dptw_resp_bits_ppn = ptw_io_requestor_3_resp_bits_ppn;
  assign io_rocc_dptw_resp_bits_error = ptw_io_requestor_3_resp_bits_error;
  assign io_rocc_dptw_resp_valid = ptw_io_requestor_3_resp_valid;
  assign io_rocc_dptw_req_ready = ptw_io_requestor_3_req_ready;
  assign io_rocc_iptw_sret = ptw_io_requestor_2_sret;
  assign io_rocc_iptw_invalidate = ptw_io_requestor_2_invalidate;
  assign io_rocc_iptw_status_s = ptw_io_requestor_2_status_s;
  assign io_rocc_iptw_status_ps = ptw_io_requestor_2_status_ps;
  assign io_rocc_iptw_status_ei = ptw_io_requestor_2_status_ei;
  assign io_rocc_iptw_status_pei = ptw_io_requestor_2_status_pei;
  assign io_rocc_iptw_status_ef = ptw_io_requestor_2_status_ef;
  assign io_rocc_iptw_status_u64 = ptw_io_requestor_2_status_u64;
  assign io_rocc_iptw_status_s64 = ptw_io_requestor_2_status_s64;
  assign io_rocc_iptw_status_vm = ptw_io_requestor_2_status_vm;
  assign io_rocc_iptw_status_er = ptw_io_requestor_2_status_er;
  assign io_rocc_iptw_status_zero = ptw_io_requestor_2_status_zero;
  assign io_rocc_iptw_status_im = ptw_io_requestor_2_status_im;
  assign io_rocc_iptw_status_ip = ptw_io_requestor_2_status_ip;
  assign io_rocc_iptw_resp_bits_perm = ptw_io_requestor_2_resp_bits_perm;
  assign io_rocc_iptw_resp_bits_ppn = ptw_io_requestor_2_resp_bits_ppn;
  assign io_rocc_iptw_resp_bits_error = ptw_io_requestor_2_resp_bits_error;
  assign io_rocc_iptw_resp_valid = ptw_io_requestor_2_resp_valid;
  assign io_rocc_iptw_req_ready = ptw_io_requestor_2_req_ready;
  assign io_rocc_imem_finish_ready = memArb_io_in_2_finish_ready;
  assign io_rocc_imem_grant_bits_payload_g_type = memArb_io_in_2_grant_bits_payload_g_type;
  assign io_rocc_imem_grant_bits_payload_uncached = memArb_io_in_2_grant_bits_payload_uncached;
  assign io_rocc_imem_grant_bits_payload_master_xact_id = memArb_io_in_2_grant_bits_payload_master_xact_id;
  assign io_rocc_imem_grant_bits_payload_client_xact_id = memArb_io_in_2_grant_bits_payload_client_xact_id;
  assign io_rocc_imem_grant_bits_payload_data = memArb_io_in_2_grant_bits_payload_data;
  assign io_rocc_imem_grant_bits_header_dst = memArb_io_in_2_grant_bits_header_dst;
  assign io_rocc_imem_grant_bits_header_src = memArb_io_in_2_grant_bits_header_src;
  assign io_rocc_imem_grant_valid = memArb_io_in_2_grant_valid;
  assign io_rocc_imem_acquire_ready = memArb_io_in_2_acquire_ready;
  assign io_rocc_s = core_io_rocc_s;
  assign io_rocc_mem_resp_bits_store_data = SimpleHellaCacheIF_io_requestor_resp_bits_store_data;
  assign io_rocc_mem_resp_bits_addr = SimpleHellaCacheIF_io_requestor_resp_bits_addr;
  assign io_rocc_mem_resp_bits_cmd = SimpleHellaCacheIF_io_requestor_resp_bits_cmd;
  assign io_rocc_mem_resp_bits_tag = SimpleHellaCacheIF_io_requestor_resp_bits_tag;
  assign io_rocc_mem_resp_bits_data_subword = SimpleHellaCacheIF_io_requestor_resp_bits_data_subword;
  assign io_rocc_mem_resp_bits_has_data = SimpleHellaCacheIF_io_requestor_resp_bits_has_data;
  assign io_rocc_mem_resp_bits_typ = SimpleHellaCacheIF_io_requestor_resp_bits_typ;
  assign io_rocc_mem_resp_bits_replay = SimpleHellaCacheIF_io_requestor_resp_bits_replay;
  assign io_rocc_mem_resp_bits_nack = SimpleHellaCacheIF_io_requestor_resp_bits_nack;
  assign io_rocc_mem_resp_bits_data = SimpleHellaCacheIF_io_requestor_resp_bits_data;
  assign io_rocc_mem_resp_valid = SimpleHellaCacheIF_io_requestor_resp_valid;
  assign io_rocc_mem_req_ready = SimpleHellaCacheIF_io_requestor_req_ready;
  assign io_rocc_resp_ready = core_io_rocc_resp_ready;
  assign io_rocc_cmd_bits_rs2 = core_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = core_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = core_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = core_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = core_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = core_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = core_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = core_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = core_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = core_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = core_io_rocc_cmd_valid;
  assign io_temac_sfp_tx_disable = core_io_temac_sfp_tx_disable;
  assign io_temac_s_axi_rready = core_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = core_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = core_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = core_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = core_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = core_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = core_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = core_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = core_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = core_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = core_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = core_io_temac_rx_axis_fifo_tready;
  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_tilelink_release_bits_payload_r_type = dcache_io_mem_release_bits_payload_r_type;
  assign io_tilelink_release_bits_payload_data = dcache_io_mem_release_bits_payload_data;
  assign io_tilelink_release_bits_payload_client_xact_id = T1;
  assign T1 = T0[2'h2:1'h0];
  assign T0 = {dcache_io_mem_release_bits_payload_client_xact_id, 2'h0};
  assign io_tilelink_release_bits_payload_addr = dcache_io_mem_release_bits_payload_addr;
  assign io_tilelink_release_bits_header_dst = dcache_io_mem_release_bits_header_dst;
  assign io_tilelink_release_bits_header_src = dcache_io_mem_release_bits_header_src;
  assign io_tilelink_release_valid = dcache_io_mem_release_valid;
  assign io_tilelink_probe_ready = dcache_io_mem_probe_ready;
  assign io_tilelink_finish_bits_payload_master_xact_id = memArb_io_out_finish_bits_payload_master_xact_id;
  assign io_tilelink_finish_bits_header_dst = memArb_io_out_finish_bits_header_dst;
  assign io_tilelink_finish_bits_header_src = memArb_io_out_finish_bits_header_src;
  assign io_tilelink_finish_valid = memArb_io_out_finish_valid;
  assign io_tilelink_grant_ready = memArb_io_out_grant_ready;
  assign io_tilelink_acquire_bits_payload_subblock = memArb_io_out_acquire_bits_payload_subblock;
  assign io_tilelink_acquire_bits_payload_a_type = memArb_io_out_acquire_bits_payload_a_type;
  assign io_tilelink_acquire_bits_payload_uncached = memArb_io_out_acquire_bits_payload_uncached;
  assign io_tilelink_acquire_bits_payload_data = memArb_io_out_acquire_bits_payload_data;
  assign io_tilelink_acquire_bits_payload_client_xact_id = memArb_io_out_acquire_bits_payload_client_xact_id;
  assign io_tilelink_acquire_bits_payload_addr = memArb_io_out_acquire_bits_payload_addr;
  assign io_tilelink_acquire_bits_header_dst = memArb_io_out_acquire_bits_header_dst;
  assign io_tilelink_acquire_bits_header_src = memArb_io_out_acquire_bits_header_src;
  assign io_tilelink_acquire_valid = memArb_io_out_acquire_valid;
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_cpu_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_cpu_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_mispredict( core_io_imem_btb_update_bits_mispredict ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_cpu_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_0_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_0_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_0_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_0_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_0_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_0_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_0_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_0_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_0_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_0_sret ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_mem_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( icache_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( icache_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_1_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( memArb_io_in_1_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_1_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_cpu_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_1_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_1_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_1_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_1_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_1_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_1_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_1_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_1_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_1_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_1_sret ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_mem_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_mem_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_mem_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( dcache_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( dcache_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_0_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( memArb_io_in_0_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_0_finish_ready ),
       .io_mem_finish_valid( dcache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_tilelink_probe_valid ),
       .io_mem_probe_bits_header_src( io_tilelink_probe_bits_header_src ),
       .io_mem_probe_bits_header_dst( io_tilelink_probe_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( io_tilelink_probe_bits_payload_addr ),
       .io_mem_probe_bits_payload_p_type( io_tilelink_probe_bits_payload_p_type ),
       .io_mem_release_ready( io_tilelink_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_mem_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_mem_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_4_req_ready( ptw_io_requestor_4_req_ready ),
       .io_requestor_4_req_valid( io_rocc_pptw_req_valid ),
       .io_requestor_4_req_bits( io_rocc_pptw_req_bits ),
       .io_requestor_4_resp_valid( ptw_io_requestor_4_resp_valid ),
       .io_requestor_4_resp_bits_error( ptw_io_requestor_4_resp_bits_error ),
       .io_requestor_4_resp_bits_ppn( ptw_io_requestor_4_resp_bits_ppn ),
       .io_requestor_4_resp_bits_perm( ptw_io_requestor_4_resp_bits_perm ),
       .io_requestor_4_status_ip( ptw_io_requestor_4_status_ip ),
       .io_requestor_4_status_im( ptw_io_requestor_4_status_im ),
       .io_requestor_4_status_zero( ptw_io_requestor_4_status_zero ),
       .io_requestor_4_status_er( ptw_io_requestor_4_status_er ),
       .io_requestor_4_status_vm( ptw_io_requestor_4_status_vm ),
       .io_requestor_4_status_s64( ptw_io_requestor_4_status_s64 ),
       .io_requestor_4_status_u64( ptw_io_requestor_4_status_u64 ),
       .io_requestor_4_status_ef( ptw_io_requestor_4_status_ef ),
       .io_requestor_4_status_pei( ptw_io_requestor_4_status_pei ),
       .io_requestor_4_status_ei( ptw_io_requestor_4_status_ei ),
       .io_requestor_4_status_ps( ptw_io_requestor_4_status_ps ),
       .io_requestor_4_status_s( ptw_io_requestor_4_status_s ),
       .io_requestor_4_invalidate( ptw_io_requestor_4_invalidate ),
       .io_requestor_4_sret( ptw_io_requestor_4_sret ),
       .io_requestor_3_req_ready( ptw_io_requestor_3_req_ready ),
       .io_requestor_3_req_valid( io_rocc_dptw_req_valid ),
       .io_requestor_3_req_bits( io_rocc_dptw_req_bits ),
       .io_requestor_3_resp_valid( ptw_io_requestor_3_resp_valid ),
       .io_requestor_3_resp_bits_error( ptw_io_requestor_3_resp_bits_error ),
       .io_requestor_3_resp_bits_ppn( ptw_io_requestor_3_resp_bits_ppn ),
       .io_requestor_3_resp_bits_perm( ptw_io_requestor_3_resp_bits_perm ),
       .io_requestor_3_status_ip( ptw_io_requestor_3_status_ip ),
       .io_requestor_3_status_im( ptw_io_requestor_3_status_im ),
       .io_requestor_3_status_zero( ptw_io_requestor_3_status_zero ),
       .io_requestor_3_status_er( ptw_io_requestor_3_status_er ),
       .io_requestor_3_status_vm( ptw_io_requestor_3_status_vm ),
       .io_requestor_3_status_s64( ptw_io_requestor_3_status_s64 ),
       .io_requestor_3_status_u64( ptw_io_requestor_3_status_u64 ),
       .io_requestor_3_status_ef( ptw_io_requestor_3_status_ef ),
       .io_requestor_3_status_pei( ptw_io_requestor_3_status_pei ),
       .io_requestor_3_status_ei( ptw_io_requestor_3_status_ei ),
       .io_requestor_3_status_ps( ptw_io_requestor_3_status_ps ),
       .io_requestor_3_status_s( ptw_io_requestor_3_status_s ),
       .io_requestor_3_invalidate( ptw_io_requestor_3_invalidate ),
       .io_requestor_3_sret( ptw_io_requestor_3_sret ),
       .io_requestor_2_req_ready( ptw_io_requestor_2_req_ready ),
       .io_requestor_2_req_valid( io_rocc_iptw_req_valid ),
       .io_requestor_2_req_bits( io_rocc_iptw_req_bits ),
       .io_requestor_2_resp_valid( ptw_io_requestor_2_resp_valid ),
       .io_requestor_2_resp_bits_error( ptw_io_requestor_2_resp_bits_error ),
       .io_requestor_2_resp_bits_ppn( ptw_io_requestor_2_resp_bits_ppn ),
       .io_requestor_2_resp_bits_perm( ptw_io_requestor_2_resp_bits_perm ),
       .io_requestor_2_status_ip( ptw_io_requestor_2_status_ip ),
       .io_requestor_2_status_im( ptw_io_requestor_2_status_im ),
       .io_requestor_2_status_zero( ptw_io_requestor_2_status_zero ),
       .io_requestor_2_status_er( ptw_io_requestor_2_status_er ),
       .io_requestor_2_status_vm( ptw_io_requestor_2_status_vm ),
       .io_requestor_2_status_s64( ptw_io_requestor_2_status_s64 ),
       .io_requestor_2_status_u64( ptw_io_requestor_2_status_u64 ),
       .io_requestor_2_status_ef( ptw_io_requestor_2_status_ef ),
       .io_requestor_2_status_pei( ptw_io_requestor_2_status_pei ),
       .io_requestor_2_status_ei( ptw_io_requestor_2_status_ei ),
       .io_requestor_2_status_ps( ptw_io_requestor_2_status_ps ),
       .io_requestor_2_status_s( ptw_io_requestor_2_status_s ),
       .io_requestor_2_invalidate( ptw_io_requestor_2_invalidate ),
       .io_requestor_2_sret( ptw_io_requestor_2_sret ),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_requestor_1_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_requestor_1_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_requestor_1_status_ip( ptw_io_requestor_1_status_ip ),
       .io_requestor_1_status_im( ptw_io_requestor_1_status_im ),
       .io_requestor_1_status_zero( ptw_io_requestor_1_status_zero ),
       .io_requestor_1_status_er( ptw_io_requestor_1_status_er ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_requestor_1_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_requestor_1_status_ef( ptw_io_requestor_1_status_ef ),
       .io_requestor_1_status_pei( ptw_io_requestor_1_status_pei ),
       .io_requestor_1_status_ei( ptw_io_requestor_1_status_ei ),
       .io_requestor_1_status_ps( ptw_io_requestor_1_status_ps ),
       .io_requestor_1_status_s( ptw_io_requestor_1_status_s ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_1_sret( ptw_io_requestor_1_sret ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_requestor_0_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_requestor_0_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_requestor_0_status_ip( ptw_io_requestor_0_status_ip ),
       .io_requestor_0_status_im( ptw_io_requestor_0_status_im ),
       .io_requestor_0_status_zero( ptw_io_requestor_0_status_zero ),
       .io_requestor_0_status_er( ptw_io_requestor_0_status_er ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_requestor_0_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_requestor_0_status_ef( ptw_io_requestor_0_status_ef ),
       .io_requestor_0_status_pei( ptw_io_requestor_0_status_pei ),
       .io_requestor_0_status_ei( ptw_io_requestor_0_status_ei ),
       .io_requestor_0_status_ps( ptw_io_requestor_0_status_ps ),
       .io_requestor_0_status_s( ptw_io_requestor_0_status_s ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_requestor_0_sret( ptw_io_requestor_0_sret ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       //.io_mem_req_bits_data(  )
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       //.io_mem_ptw_req_valid(  )
       //.io_mem_ptw_req_bits(  )
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_sret( core_io_ptw_sret ),
       .io_dpath_status_ip( core_io_ptw_status_ip ),
       .io_dpath_status_im( core_io_ptw_status_im ),
       .io_dpath_status_zero( core_io_ptw_status_zero ),
       .io_dpath_status_er( core_io_ptw_status_er ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_s64( core_io_ptw_status_s64 ),
       .io_dpath_status_u64( core_io_ptw_status_u64 ),
       .io_dpath_status_ef( core_io_ptw_status_ef ),
       .io_dpath_status_pei( core_io_ptw_status_pei ),
       .io_dpath_status_ei( core_io_ptw_status_ei ),
       .io_dpath_status_ps( core_io_ptw_status_ps ),
       .io_dpath_status_s( core_io_ptw_status_s )
  );
  Core core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_imem_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_mispredict( core_io_imem_btb_update_bits_mispredict ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_imem_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       //.io_dmem_ptw_req_valid(  )
       //.io_dmem_ptw_req_bits(  )
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_sret( core_io_ptw_sret ),
       .io_ptw_status_ip( core_io_ptw_status_ip ),
       .io_ptw_status_im( core_io_ptw_status_im ),
       .io_ptw_status_zero( core_io_ptw_status_zero ),
       .io_ptw_status_er( core_io_ptw_status_er ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_s64( core_io_ptw_status_s64 ),
       .io_ptw_status_u64( core_io_ptw_status_u64 ),
       .io_ptw_status_ef( core_io_ptw_status_ef ),
       .io_ptw_status_pei( core_io_ptw_status_pei ),
       .io_ptw_status_ei( core_io_ptw_status_ei ),
       .io_ptw_status_ps( core_io_ptw_status_ps ),
       .io_ptw_status_s( core_io_ptw_status_s ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( core_io_rocc_cmd_valid ),
       .io_rocc_cmd_bits_inst_funct( core_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( core_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( core_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( core_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( core_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( core_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( core_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( core_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( core_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( core_io_rocc_cmd_bits_rs2 ),
       .io_rocc_resp_ready( core_io_rocc_resp_ready ),
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( core_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( core_io_rocc_exception ),
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( core_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( core_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( core_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( core_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( core_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( core_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( core_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( core_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( core_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( core_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( core_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( core_io_temac_s_axi_rready ),
       .io_temac_sfp_tx_disable( core_io_temac_sfp_tx_disable )
  );
  `ifndef SYNTHESIS
    assign core.io_dmem_ptw_req_valid = {1{$random}};
    assign core.io_dmem_ptw_req_bits = {1{$random}};
  `endif
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_2_req_ready( dcArb_io_requestor_2_req_ready ),
       .io_requestor_2_req_valid( SimpleHellaCacheIF_io_cache_req_valid ),
       .io_requestor_2_req_bits_kill( SimpleHellaCacheIF_io_cache_req_bits_kill ),
       .io_requestor_2_req_bits_typ( SimpleHellaCacheIF_io_cache_req_bits_typ ),
       .io_requestor_2_req_bits_phys( SimpleHellaCacheIF_io_cache_req_bits_phys ),
       .io_requestor_2_req_bits_addr( SimpleHellaCacheIF_io_cache_req_bits_addr ),
       .io_requestor_2_req_bits_tag( SimpleHellaCacheIF_io_cache_req_bits_tag ),
       .io_requestor_2_req_bits_cmd( SimpleHellaCacheIF_io_cache_req_bits_cmd ),
       .io_requestor_2_req_bits_data( SimpleHellaCacheIF_io_cache_req_bits_data ),
       .io_requestor_2_resp_valid( dcArb_io_requestor_2_resp_valid ),
       .io_requestor_2_resp_bits_data( dcArb_io_requestor_2_resp_bits_data ),
       .io_requestor_2_resp_bits_nack( dcArb_io_requestor_2_resp_bits_nack ),
       .io_requestor_2_resp_bits_replay( dcArb_io_requestor_2_resp_bits_replay ),
       .io_requestor_2_resp_bits_typ( dcArb_io_requestor_2_resp_bits_typ ),
       .io_requestor_2_resp_bits_has_data( dcArb_io_requestor_2_resp_bits_has_data ),
       .io_requestor_2_resp_bits_data_subword( dcArb_io_requestor_2_resp_bits_data_subword ),
       .io_requestor_2_resp_bits_tag( dcArb_io_requestor_2_resp_bits_tag ),
       .io_requestor_2_resp_bits_cmd( dcArb_io_requestor_2_resp_bits_cmd ),
       .io_requestor_2_resp_bits_addr( dcArb_io_requestor_2_resp_bits_addr ),
       .io_requestor_2_resp_bits_store_data( dcArb_io_requestor_2_resp_bits_store_data ),
       .io_requestor_2_replay_next_valid( dcArb_io_requestor_2_replay_next_valid ),
       .io_requestor_2_replay_next_bits( dcArb_io_requestor_2_replay_next_bits ),
       .io_requestor_2_xcpt_ma_ld( dcArb_io_requestor_2_xcpt_ma_ld ),
       .io_requestor_2_xcpt_ma_st( dcArb_io_requestor_2_xcpt_ma_st ),
       .io_requestor_2_xcpt_pf_ld( dcArb_io_requestor_2_xcpt_pf_ld ),
       .io_requestor_2_xcpt_pf_st( dcArb_io_requestor_2_xcpt_pf_st ),
       //.io_requestor_2_ptw_req_ready(  )
       //.io_requestor_2_ptw_req_valid(  )
       //.io_requestor_2_ptw_req_bits(  )
       //.io_requestor_2_ptw_resp_valid(  )
       //.io_requestor_2_ptw_resp_bits_error(  )
       //.io_requestor_2_ptw_resp_bits_ppn(  )
       //.io_requestor_2_ptw_resp_bits_perm(  )
       //.io_requestor_2_ptw_status_ip(  )
       //.io_requestor_2_ptw_status_im(  )
       //.io_requestor_2_ptw_status_zero(  )
       //.io_requestor_2_ptw_status_er(  )
       //.io_requestor_2_ptw_status_vm(  )
       //.io_requestor_2_ptw_status_s64(  )
       //.io_requestor_2_ptw_status_u64(  )
       //.io_requestor_2_ptw_status_ef(  )
       //.io_requestor_2_ptw_status_pei(  )
       //.io_requestor_2_ptw_status_ei(  )
       //.io_requestor_2_ptw_status_ps(  )
       //.io_requestor_2_ptw_status_s(  )
       //.io_requestor_2_ptw_invalidate(  )
       //.io_requestor_2_ptw_sret(  )
       .io_requestor_2_ordered( dcArb_io_requestor_2_ordered ),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_requestor_1_ptw_req_ready(  )
       //.io_requestor_1_ptw_req_valid(  )
       //.io_requestor_1_ptw_req_bits(  )
       //.io_requestor_1_ptw_resp_valid(  )
       //.io_requestor_1_ptw_resp_bits_error(  )
       //.io_requestor_1_ptw_resp_bits_ppn(  )
       //.io_requestor_1_ptw_resp_bits_perm(  )
       //.io_requestor_1_ptw_status_ip(  )
       //.io_requestor_1_ptw_status_im(  )
       //.io_requestor_1_ptw_status_zero(  )
       //.io_requestor_1_ptw_status_er(  )
       //.io_requestor_1_ptw_status_vm(  )
       //.io_requestor_1_ptw_status_s64(  )
       //.io_requestor_1_ptw_status_u64(  )
       //.io_requestor_1_ptw_status_ef(  )
       //.io_requestor_1_ptw_status_pei(  )
       //.io_requestor_1_ptw_status_ei(  )
       //.io_requestor_1_ptw_status_ps(  )
       //.io_requestor_1_ptw_status_s(  )
       //.io_requestor_1_ptw_invalidate(  )
       //.io_requestor_1_ptw_sret(  )
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       //.io_requestor_0_req_bits_data(  )
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_ptw_req_ready(  )
       //.io_requestor_0_ptw_req_valid(  )
       //.io_requestor_0_ptw_req_bits(  )
       //.io_requestor_0_ptw_resp_valid(  )
       //.io_requestor_0_ptw_resp_bits_error(  )
       //.io_requestor_0_ptw_resp_bits_ppn(  )
       //.io_requestor_0_ptw_resp_bits_perm(  )
       //.io_requestor_0_ptw_status_ip(  )
       //.io_requestor_0_ptw_status_im(  )
       //.io_requestor_0_ptw_status_zero(  )
       //.io_requestor_0_ptw_status_er(  )
       //.io_requestor_0_ptw_status_vm(  )
       //.io_requestor_0_ptw_status_s64(  )
       //.io_requestor_0_ptw_status_u64(  )
       //.io_requestor_0_ptw_status_ef(  )
       //.io_requestor_0_ptw_status_pei(  )
       //.io_requestor_0_ptw_status_ei(  )
       //.io_requestor_0_ptw_status_ps(  )
       //.io_requestor_0_ptw_status_s(  )
       //.io_requestor_0_ptw_invalidate(  )
       //.io_requestor_0_ptw_sret(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_mem_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
  `ifndef SYNTHESIS
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
    assign dcArb.io_requestor_0_req_bits_data = {2{$random}};
  `endif
  UncachedTileLinkIOArbiterThatAppendsArbiterId memArb(.clk(clk), .reset(reset),
       .io_in_2_acquire_ready( memArb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_in_2_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_in_2_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_in_2_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_in_2_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_in_2_grant_ready( io_rocc_imem_grant_ready ),
       .io_in_2_grant_valid( memArb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( memArb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( memArb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( memArb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( memArb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_master_xact_id( memArb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_in_2_grant_bits_payload_uncached( memArb_io_in_2_grant_bits_payload_uncached ),
       .io_in_2_grant_bits_payload_g_type( memArb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( memArb_io_in_2_finish_ready ),
       .io_in_2_finish_valid( io_rocc_imem_finish_valid ),
       .io_in_2_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_in_2_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_in_2_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       .io_in_1_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_in_1_acquire_bits_header_src(  )
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_uncached( icache_io_mem_acquire_bits_payload_uncached ),
       .io_in_1_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_subblock( icache_io_mem_acquire_bits_payload_subblock ),
       .io_in_1_grant_ready( icache_io_mem_grant_ready ),
       .io_in_1_grant_valid( memArb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_uncached( memArb_io_in_1_grant_bits_payload_uncached ),
       .io_in_1_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( memArb_io_in_1_finish_ready ),
       .io_in_1_finish_valid( icache_io_mem_finish_valid ),
       .io_in_1_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_in_1_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_in_1_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_in_0_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_in_0_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_uncached( dcache_io_mem_acquire_bits_payload_uncached ),
       .io_in_0_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_subblock( dcache_io_mem_acquire_bits_payload_subblock ),
       .io_in_0_grant_ready( dcache_io_mem_grant_ready ),
       .io_in_0_grant_valid( memArb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_uncached( memArb_io_in_0_grant_bits_payload_uncached ),
       .io_in_0_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( memArb_io_in_0_finish_ready ),
       .io_in_0_finish_valid( dcache_io_mem_finish_valid ),
       .io_in_0_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_in_0_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_in_0_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_acquire_ready( io_tilelink_acquire_ready ),
       .io_out_acquire_valid( memArb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( memArb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( memArb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( memArb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( memArb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( memArb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_uncached( memArb_io_out_acquire_bits_payload_uncached ),
       .io_out_acquire_bits_payload_a_type( memArb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_subblock( memArb_io_out_acquire_bits_payload_subblock ),
       .io_out_grant_ready( memArb_io_out_grant_ready ),
       .io_out_grant_valid( io_tilelink_grant_valid ),
       .io_out_grant_bits_header_src( io_tilelink_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_tilelink_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_tilelink_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_tilelink_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_tilelink_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_uncached( io_tilelink_grant_bits_payload_uncached ),
       .io_out_grant_bits_payload_g_type( io_tilelink_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_tilelink_finish_ready ),
       .io_out_finish_valid( memArb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( memArb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( memArb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( memArb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign memArb.io_in_1_acquire_bits_header_src = {1{$random}};
    assign memArb.io_in_1_acquire_bits_header_dst = {1{$random}};
  `endif
  SimpleHellaCacheIF SimpleHellaCacheIF(.clk(clk), .reset(reset),
       .io_requestor_req_ready( SimpleHellaCacheIF_io_requestor_req_ready ),
       .io_requestor_req_valid( io_rocc_mem_req_valid ),
       .io_requestor_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_requestor_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_requestor_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_requestor_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_requestor_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_requestor_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_requestor_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_requestor_resp_valid( SimpleHellaCacheIF_io_requestor_resp_valid ),
       .io_requestor_resp_bits_data( SimpleHellaCacheIF_io_requestor_resp_bits_data ),
       .io_requestor_resp_bits_nack( SimpleHellaCacheIF_io_requestor_resp_bits_nack ),
       .io_requestor_resp_bits_replay( SimpleHellaCacheIF_io_requestor_resp_bits_replay ),
       .io_requestor_resp_bits_typ( SimpleHellaCacheIF_io_requestor_resp_bits_typ ),
       .io_requestor_resp_bits_has_data( SimpleHellaCacheIF_io_requestor_resp_bits_has_data ),
       .io_requestor_resp_bits_data_subword( SimpleHellaCacheIF_io_requestor_resp_bits_data_subword ),
       .io_requestor_resp_bits_tag( SimpleHellaCacheIF_io_requestor_resp_bits_tag ),
       .io_requestor_resp_bits_cmd( SimpleHellaCacheIF_io_requestor_resp_bits_cmd ),
       .io_requestor_resp_bits_addr( SimpleHellaCacheIF_io_requestor_resp_bits_addr ),
       .io_requestor_resp_bits_store_data( SimpleHellaCacheIF_io_requestor_resp_bits_store_data ),
       //.io_requestor_replay_next_valid(  )
       //.io_requestor_replay_next_bits(  )
       //.io_requestor_xcpt_ma_ld(  )
       //.io_requestor_xcpt_ma_st(  )
       //.io_requestor_xcpt_pf_ld(  )
       //.io_requestor_xcpt_pf_st(  )
       .io_requestor_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_requestor_ptw_req_valid(  )
       //.io_requestor_ptw_req_bits(  )
       .io_requestor_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_requestor_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_requestor_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_requestor_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_requestor_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_requestor_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_requestor_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_requestor_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_requestor_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_requestor_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_requestor_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_requestor_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_requestor_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_requestor_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_requestor_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_requestor_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_requestor_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_requestor_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_requestor_ordered(  )
       .io_cache_req_ready( dcArb_io_requestor_2_req_ready ),
       .io_cache_req_valid( SimpleHellaCacheIF_io_cache_req_valid ),
       .io_cache_req_bits_kill( SimpleHellaCacheIF_io_cache_req_bits_kill ),
       .io_cache_req_bits_typ( SimpleHellaCacheIF_io_cache_req_bits_typ ),
       .io_cache_req_bits_phys( SimpleHellaCacheIF_io_cache_req_bits_phys ),
       .io_cache_req_bits_addr( SimpleHellaCacheIF_io_cache_req_bits_addr ),
       .io_cache_req_bits_tag( SimpleHellaCacheIF_io_cache_req_bits_tag ),
       .io_cache_req_bits_cmd( SimpleHellaCacheIF_io_cache_req_bits_cmd ),
       .io_cache_req_bits_data( SimpleHellaCacheIF_io_cache_req_bits_data ),
       .io_cache_resp_valid( dcArb_io_requestor_2_resp_valid ),
       .io_cache_resp_bits_data( dcArb_io_requestor_2_resp_bits_data ),
       .io_cache_resp_bits_nack( dcArb_io_requestor_2_resp_bits_nack ),
       .io_cache_resp_bits_replay( dcArb_io_requestor_2_resp_bits_replay ),
       .io_cache_resp_bits_typ( dcArb_io_requestor_2_resp_bits_typ ),
       .io_cache_resp_bits_has_data( dcArb_io_requestor_2_resp_bits_has_data ),
       .io_cache_resp_bits_data_subword( dcArb_io_requestor_2_resp_bits_data_subword ),
       .io_cache_resp_bits_tag( dcArb_io_requestor_2_resp_bits_tag ),
       .io_cache_resp_bits_cmd( dcArb_io_requestor_2_resp_bits_cmd ),
       .io_cache_resp_bits_addr( dcArb_io_requestor_2_resp_bits_addr ),
       .io_cache_resp_bits_store_data( dcArb_io_requestor_2_resp_bits_store_data ),
       .io_cache_replay_next_valid( dcArb_io_requestor_2_replay_next_valid ),
       .io_cache_replay_next_bits( dcArb_io_requestor_2_replay_next_bits ),
       .io_cache_xcpt_ma_ld( dcArb_io_requestor_2_xcpt_ma_ld ),
       .io_cache_xcpt_ma_st( dcArb_io_requestor_2_xcpt_ma_st ),
       .io_cache_xcpt_pf_ld( dcArb_io_requestor_2_xcpt_pf_ld ),
       .io_cache_xcpt_pf_st( dcArb_io_requestor_2_xcpt_pf_st ),
       //.io_cache_ptw_req_ready(  )
       //.io_cache_ptw_req_valid(  )
       //.io_cache_ptw_req_bits(  )
       //.io_cache_ptw_resp_valid(  )
       //.io_cache_ptw_resp_bits_error(  )
       //.io_cache_ptw_resp_bits_ppn(  )
       //.io_cache_ptw_resp_bits_perm(  )
       //.io_cache_ptw_status_ip(  )
       //.io_cache_ptw_status_im(  )
       //.io_cache_ptw_status_zero(  )
       //.io_cache_ptw_status_er(  )
       //.io_cache_ptw_status_vm(  )
       //.io_cache_ptw_status_s64(  )
       //.io_cache_ptw_status_u64(  )
       //.io_cache_ptw_status_ef(  )
       //.io_cache_ptw_status_pei(  )
       //.io_cache_ptw_status_ei(  )
       //.io_cache_ptw_status_ps(  )
       //.io_cache_ptw_status_s(  )
       //.io_cache_ptw_invalidate(  )
       //.io_cache_ptw_sret(  )
       .io_cache_ordered( dcArb_io_requestor_2_ordered )
  );
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [2:0] io_enq_bits_client_xact_id,
    input [511:0] io_enq_bits_data,
    input  io_enq_bits_uncached,
    input [1:0] io_enq_bits_a_type,
    input [511:0] io_enq_bits_subblock,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[2:0] io_deq_bits_client_xact_id,
    output[511:0] io_deq_bits_data,
    output io_deq_bits_uncached,
    output[1:0] io_deq_bits_a_type,
    output[511:0] io_deq_bits_subblock,
    output io_count
);

  wire T19;
  wire[1:0] T0;
  reg  full;
  wire T20;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[511:0] T3;
  wire[1055:0] T4;
  reg [1055:0] ram [0:0];
  wire[1055:0] T5;
  wire[1055:0] T6;
  wire[1055:0] T7;
  wire[514:0] T8;
  wire[513:0] T9;
  wire[540:0] T10;
  wire[514:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[511:0] T14;
  wire[2:0] T15;
  wire[25:0] T16;
  wire T17;
  wire empty;
  wire T18;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {33{$random}};
  end
`endif

  assign io_count = T19;
  assign T19 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T20 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_subblock = T3;
  assign T3 = T4[9'h1ff:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T10, T8};
  assign T8 = {io_enq_bits_uncached, T9};
  assign T9 = {io_enq_bits_a_type, io_enq_bits_subblock};
  assign T10 = {io_enq_bits_addr, T11};
  assign T11 = {io_enq_bits_client_xact_id, io_enq_bits_data};
  assign io_deq_bits_a_type = T12;
  assign T12 = T4[10'h201:10'h200];
  assign io_deq_bits_uncached = T13;
  assign T13 = T4[10'h202:10'h202];
  assign io_deq_bits_data = T14;
  assign T14 = T4[11'h402:10'h203];
  assign io_deq_bits_client_xact_id = T15;
  assign T15 = T4[11'h405:11'h403];
  assign io_deq_bits_addr = T16;
  assign T16 = T4[11'h41f:11'h406];
  assign io_deq_valid = T17;
  assign T17 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[4:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[2:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[511:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [2:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    //output[1:0] io_mem_finish_bits_header_src
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    //output[1:0] io_mem_release_bits_header_src
    //output[1:0] io_mem_release_bits_header_dst
    output[25:0] io_mem_release_bits_payload_addr,
    output[2:0] io_mem_release_bits_payload_client_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[511:0] T348;
  wire[511:0] T349;
  wire[511:0] T350;
  wire T351;
  reg [3:0] cmd;
  wire[3:0] T20;
  wire[3:0] next_cmd;
  wire[63:0] rx_shifter_in;
  wire[47:0] T30;
  reg [63:0] rx_shifter;
  wire[63:0] T31;
  wire T59;
  wire T21;
  wire T22;
  reg [14:0] rx_count;
  wire[14:0] T338;
  wire[14:0] T23;
  wire[14:0] T24;
  wire[14:0] T25;
  wire T26;
  wire T27;
  wire[12:0] T339;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T28;
  wire[11:0] T29;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire nack;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire bad_mem_packet;
  wire T44;
  wire[2:0] T45;
  reg [39:0] addr;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire T96;
  wire T97;
  reg [3:0] state;
  wire[3:0] T337;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  wire[3:0] rx_cmd;
  wire T60;
  wire[12:0] rx_word_count;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire rx_done;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire T69;
  wire[12:0] T341;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire rx_word_done;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  reg  mem_acked;
  wire T342;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire[3:0] T88;
  wire T89;
  wire T90;
  reg [8:0] pos;
  wire[8:0] T91;
  wire[8:0] T92;
  wire[8:0] T93;
  wire[8:0] T94;
  wire T95;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T112;
  wire T113;
  wire T114;
  wire[4:0] pcr_addr;
  wire T115;
  wire T116;
  wire[1:0] pcr_coreid;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T340;
  wire[14:0] T55;
  wire[14:0] T56;
  wire[14:0] T57;
  wire T58;
  wire T102;
  wire tx_done;
  wire T103;
  wire T104;
  wire T105;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T106;
  wire T107;
  wire T108;
  wire[12:0] T343;
  wire T109;
  wire T110;
  wire[1:0] tx_subword_count;
  wire T111;
  wire[1:0] T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire T355;
  wire T356;
  wire T357;
  wire[511:0] T358;
  wire[511:0] T359;
  wire[511:0] T360;
  wire[2:0] T361;
  wire[2:0] T362;
  wire[2:0] T363;
  wire[25:0] T364;
  wire[25:0] T365;
  wire[25:0] T366;
  wire[36:0] init_addr;
  wire[39:0] T367;
  wire[25:0] T368;
  wire[25:0] T369;
  wire T370;
  wire T371;
  wire T372;
  wire[63:0] pcr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  wire[63:0] T121;
  wire[63:0] T122;
  wire T123;
  wire T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire T128;
  wire[63:0] T129;
  wire[63:0] T130;
  wire T131;
  wire T132;
  wire[63:0] T133;
  wire[63:0] T134;
  wire T135;
  wire T136;
  wire[63:0] T137;
  wire[63:0] T138;
  wire T139;
  wire T140;
  wire[63:0] T141;
  wire[63:0] T142;
  wire T143;
  wire T144;
  wire[63:0] T145;
  wire[63:0] T146;
  wire T147;
  wire T148;
  wire[63:0] T149;
  wire T150;
  wire[2:0] T151;
  wire[2:0] T152;
  wire[5:0] T153;
  wire[5:0] scr_addr;
  wire T154;
  wire T155;
  reg [2:0] mem_gxid;
  wire[2:0] T156;
  reg [1:0] mem_gsrc;
  wire[1:0] T157;
  wire T158;
  reg  mem_needs_ack;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[511:0] mem_req_data;
  wire[447:0] T163;
  wire[383:0] T164;
  wire[319:0] T165;
  wire[255:0] T166;
  wire[191:0] T167;
  wire[127:0] T168;
  wire[63:0] T169;
  wire[63:0] T170;
  wire[63:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[63:0] T174;
  wire[63:0] T175;
  wire[63:0] T176;
  reg  R177;
  wire T344;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg  R187;
  wire T345;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire[15:0] T346;
  wire[63:0] T192;
  wire[5:0] T193;
  wire[1:0] T194;
  wire[63:0] tx_data;
  wire[63:0] T195;
  wire[63:0] T196;
  reg [63:0] pcrReadData;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T199;
  wire[63:0] T347;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  wire[63:0] T203;
  wire[63:0] T204;
  wire[63:0] T205;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T206;
  wire[5:0] T207;
  wire[63:0] T208;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T209;
  wire T210;
  wire[63:0] T211;
  wire[63:0] T212;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T213;
  wire[63:0] T214;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T215;
  wire T216;
  wire T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] T220;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T221;
  wire[63:0] T222;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T223;
  wire T224;
  wire[63:0] T225;
  wire[63:0] T226;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T227;
  wire[63:0] T228;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire[63:0] T233;
  wire[63:0] T234;
  wire[63:0] T235;
  wire[63:0] T236;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T237;
  wire[63:0] T238;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T239;
  wire T240;
  wire[63:0] T241;
  wire[63:0] T242;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T243;
  wire[63:0] T244;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T245;
  wire T246;
  wire T247;
  wire[63:0] T248;
  wire[63:0] T249;
  wire[63:0] T250;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T251;
  wire[63:0] T252;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T253;
  wire T254;
  wire[63:0] T255;
  wire[63:0] T256;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T257;
  wire[63:0] T258;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[63:0] T264;
  wire[63:0] T265;
  wire[63:0] T266;
  wire[63:0] T267;
  wire[63:0] T268;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T269;
  wire[63:0] T270;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T271;
  wire T272;
  wire[63:0] T273;
  wire[63:0] T274;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T275;
  wire[63:0] T276;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T277;
  wire T278;
  wire T279;
  wire[63:0] T280;
  wire[63:0] T281;
  wire[63:0] T282;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T283;
  wire[63:0] T284;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T285;
  wire T286;
  wire[63:0] T287;
  wire[63:0] T288;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T289;
  wire[63:0] T290;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire[63:0] T295;
  wire[63:0] T296;
  wire[63:0] T297;
  wire[63:0] T298;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T299;
  wire[63:0] T300;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T301;
  wire T302;
  wire[63:0] T303;
  wire[63:0] T304;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T305;
  wire[63:0] T306;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T307;
  wire T308;
  wire T309;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] T312;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T313;
  wire[63:0] T314;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T315;
  wire T316;
  wire[63:0] T317;
  wire[63:0] T318;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T319;
  wire[63:0] T320;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[63:0] tx_header;
  wire[15:0] T330;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T331;
  reg [7:0] seqno;
  wire[7:0] T332;
  wire[7:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire acq_q_io_enq_ready;
  wire acq_q_io_deq_valid;
  wire[25:0] acq_q_io_deq_bits_addr;
  wire[2:0] acq_q_io_deq_bits_client_xact_id;
  wire acq_q_io_deq_bits_uncached;
  wire[1:0] acq_q_io_deq_bits_a_type;
  wire[511:0] acq_q_io_deq_bits_subblock;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cmd = {1{$random}};
    rx_shifter = {2{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    addr = {2{$random}};
    state = {1{$random}};
    mem_acked = {1{$random}};
    pos = {1{$random}};
    tx_count = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    mem_gxid = {1{$random}};
    mem_gsrc = {1{$random}};
    mem_needs_ack = {1{$random}};
    R177 = {1{$random}};
    R187 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
`endif

  assign T348 = T351 ? T350 : T349;
  assign T349 = 512'h7;
  assign T350 = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
  assign T351 = cmd == 4'h1;
  assign T20 = T21 ? next_cmd : cmd;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign rx_shifter_in = {io_host_in_bits, T30};
  assign T30 = rx_shifter[6'h3f:5'h10];
  assign T31 = T59 ? rx_shifter_in : rx_shifter;
  assign T59 = io_host_in_valid & io_host_in_ready;
  assign T21 = T59 & T22;
  assign T22 = rx_count == 15'h3;
  assign T338 = reset ? 15'h0 : T23;
  assign T23 = T26 ? 15'h0 : T24;
  assign T24 = T59 ? T25 : rx_count;
  assign T25 = rx_count + 15'h1;
  assign T26 = T102 & T27;
  assign T27 = tx_word_count == T339;
  assign T339 = {1'h0, tx_size};
  assign tx_size = T32 ? size : 12'h0;
  assign T28 = T21 ? T29 : size;
  assign T29 = rx_shifter_in[4'hf:3'h4];
  assign T32 = T38 & T33;
  assign T33 = T35 | T34;
  assign T34 = cmd == 4'h3;
  assign T35 = T37 | T36;
  assign T36 = cmd == 4'h2;
  assign T37 = cmd == 4'h0;
  assign T38 = nack ^ 1'h1;
  assign nack = T52 ? bad_mem_packet : T39;
  assign T39 = T41 ? T40 : 1'h1;
  assign T40 = size != 12'h1;
  assign T41 = T43 | T42;
  assign T42 = cmd == 4'h3;
  assign T43 = cmd == 4'h2;
  assign bad_mem_packet = T50 | T44;
  assign T44 = T45 != 3'h0;
  assign T45 = addr[2'h2:1'h0];
  assign T46 = T96 ? T49 : T47;
  assign T47 = T21 ? T48 : addr;
  assign T48 = rx_shifter_in[6'h3f:5'h18];
  assign T49 = addr + 40'h8;
  assign T96 = T97 & io_mem_finish_ready;
  assign T97 = state == 4'h7;
  assign T337 = reset ? 4'h0 : T4;
  assign T4 = T118 ? 4'h8 : T5;
  assign T5 = io_cpu_0_pcr_rep_valid ? 4'h8 : T6;
  assign T6 = T113 ? 4'h8 : T7;
  assign T7 = T112 ? 4'h2 : T8;
  assign T8 = T102 ? T98 : T9;
  assign T9 = T96 ? T88 : T10;
  assign T10 = T87 ? 4'h7 : T11;
  assign T11 = T81 ? 4'h7 : T12;
  assign T12 = T79 ? 4'h5 : T13;
  assign T13 = T77 ? 4'h6 : T14;
  assign T14 = T64 ? T15 : state;
  assign T15 = T63 ? 4'h3 : T16;
  assign T16 = T62 ? 4'h4 : T17;
  assign T17 = T18 ? 4'h1 : 4'h8;
  assign T18 = T61 | T19;
  assign T19 = rx_cmd == 4'h3;
  assign rx_cmd = T60 ? next_cmd : cmd;
  assign T60 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T61 = rx_cmd == 4'h2;
  assign T62 = rx_cmd == 4'h1;
  assign T63 = rx_cmd == 4'h0;
  assign T64 = T76 & rx_done;
  assign rx_done = rx_word_done & T65;
  assign T65 = T73 ? T70 : T66;
  assign T66 = T69 | T67;
  assign T67 = T68 == 3'h0;
  assign T68 = rx_word_count[2'h2:1'h0];
  assign T69 = rx_word_count == T341;
  assign T341 = {1'h0, size};
  assign T70 = T72 & T71;
  assign T71 = next_cmd != 4'h3;
  assign T72 = next_cmd != 4'h1;
  assign T73 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T74;
  assign T74 = T75 == 2'h3;
  assign T75 = rx_count[1'h1:1'h0];
  assign T76 = state == 4'h0;
  assign T77 = T78 & acq_q_io_enq_ready;
  assign T78 = state == 4'h4;
  assign T79 = T80 & acq_q_io_enq_ready;
  assign T80 = state == 4'h3;
  assign T81 = T86 & mem_acked;
  assign T342 = reset ? 1'h0 : T82;
  assign T82 = T85 ? 1'h0 : T83;
  assign T83 = T81 ? 1'h0 : T84;
  assign T84 = io_mem_grant_valid ? 1'h1 : mem_acked;
  assign T85 = state == 4'h5;
  assign T86 = state == 4'h6;
  assign T87 = T85 & io_mem_grant_valid;
  assign T88 = T89 ? 4'h8 : 4'h0;
  assign T89 = T95 | T90;
  assign T90 = pos == 9'h1;
  assign T91 = T96 ? T94 : T92;
  assign T92 = T21 ? T93 : pos;
  assign T93 = rx_shifter_in[4'hf:3'h7];
  assign T94 = pos - 9'h1;
  assign T95 = cmd == 4'h0;
  assign T98 = T99 ? 4'h3 : 4'h0;
  assign T99 = T101 & T100;
  assign T100 = pos != 9'h0;
  assign T101 = cmd == 4'h0;
  assign T112 = io_cpu_0_pcr_req_valid & io_cpu_0_pcr_req_ready;
  assign T113 = T115 & T114;
  assign T114 = pcr_addr == 5'h1d;
  assign pcr_addr = addr[3'h4:1'h0];
  assign T115 = T117 & T116;
  assign T116 = pcr_coreid == 2'h0;
  assign pcr_coreid = addr[5'h15:5'h14];
  assign T117 = state == 4'h1;
  assign T118 = T120 & T119;
  assign T119 = pcr_coreid == 2'h3;
  assign T120 = state == 4'h1;
  assign T50 = T51 != 3'h0;
  assign T51 = size[2'h2:1'h0];
  assign T52 = T54 | T53;
  assign T53 = cmd == 4'h1;
  assign T54 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T340 = reset ? 15'h0 : T55;
  assign T55 = T26 ? 15'h0 : T56;
  assign T56 = T58 ? T57 : tx_count;
  assign T57 = tx_count + 15'h1;
  assign T58 = io_host_out_valid & io_host_out_ready;
  assign T102 = T111 & tx_done;
  assign tx_done = T109 & T103;
  assign T103 = T108 | T104;
  assign T104 = T107 & T105;
  assign T105 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T106 - 3'h1;
  assign T106 = tx_word_count[2'h2:1'h0];
  assign T107 = 13'h0 < tx_word_count;
  assign T108 = tx_word_count == T343;
  assign T343 = {1'h0, tx_size};
  assign T109 = io_host_out_ready & T110;
  assign T110 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T111 = state == 4'h8;
  assign T352 = T351 ? T354 : T353;
  assign T353 = 2'h0;
  assign T354 = 2'h1;
  assign T355 = T351 ? T357 : T356;
  assign T356 = 1'h1;
  assign T357 = 1'h1;
  assign T358 = T351 ? T360 : T359;
  assign T359 = 512'h0;
  assign T360 = 512'h0;
  assign T361 = T351 ? T363 : T362;
  assign T362 = 3'h0;
  assign T363 = 3'h0;
  assign T364 = T351 ? T368 : T365;
  assign T365 = T366;
  assign T366 = init_addr[5'h19:1'h0];
  assign init_addr = T367 >> 2'h3;
  assign T367 = addr;
  assign T368 = T369;
  assign T369 = init_addr[5'h19:1'h0];
  assign T370 = T372 | T371;
  assign T371 = state == 4'h4;
  assign T372 = state == 4'h3;
  assign io_scr_wdata = pcr_wdata;
  assign pcr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_payload_data[9'h1ff:9'h1c0];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 4'h5;
  assign T122 = io_mem_grant_bits_payload_data[9'h1bf:9'h180];
  assign T123 = T124 & io_mem_grant_valid;
  assign T124 = state == 4'h5;
  assign T126 = io_mem_grant_bits_payload_data[9'h17f:9'h140];
  assign T127 = T128 & io_mem_grant_valid;
  assign T128 = state == 4'h5;
  assign T130 = io_mem_grant_bits_payload_data[9'h13f:9'h100];
  assign T131 = T132 & io_mem_grant_valid;
  assign T132 = state == 4'h5;
  assign T134 = io_mem_grant_bits_payload_data[8'hff:8'hc0];
  assign T135 = T136 & io_mem_grant_valid;
  assign T136 = state == 4'h5;
  assign T138 = io_mem_grant_bits_payload_data[8'hbf:8'h80];
  assign T139 = T140 & io_mem_grant_valid;
  assign T140 = state == 4'h5;
  assign T142 = io_mem_grant_bits_payload_data[7'h7f:7'h40];
  assign T143 = T144 & io_mem_grant_valid;
  assign T144 = state == 4'h5;
  assign T146 = io_mem_grant_bits_payload_data[6'h3f:1'h0];
  assign T147 = T148 & io_mem_grant_valid;
  assign T148 = state == 4'h5;
  assign T150 = rx_word_done & io_host_in_ready;
  assign T151 = T152 - 3'h1;
  assign T152 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T153;
  assign T153 = scr_addr;
  assign scr_addr = addr[3'h5:1'h0];
  assign io_scr_wen = T154;
  assign T154 = T118 ? T155 : 1'h0;
  assign T155 = cmd == 4'h3;
  assign io_mem_release_valid = 1'h0;
  assign io_mem_probe_ready = 1'h0;
  assign io_mem_finish_bits_payload_master_xact_id = mem_gxid;
  assign T156 = io_mem_grant_valid ? io_mem_grant_bits_payload_master_xact_id : mem_gxid;
  assign io_mem_finish_bits_header_dst = mem_gsrc;
  assign T157 = io_mem_grant_valid ? io_mem_grant_bits_header_src : mem_gsrc;
  assign io_mem_finish_valid = T158;
  assign T158 = T162 & mem_needs_ack;
  assign T159 = io_mem_grant_valid ? T160 : mem_needs_ack;
  assign T160 = io_mem_grant_bits_payload_uncached | T161;
  assign T161 = io_mem_grant_bits_payload_g_type != 2'h0;
  assign T162 = state == 4'h7;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_payload_subblock = acq_q_io_deq_bits_subblock;
  assign io_mem_acquire_bits_payload_a_type = acq_q_io_deq_bits_a_type;
  assign io_mem_acquire_bits_payload_uncached = acq_q_io_deq_bits_uncached;
  assign io_mem_acquire_bits_payload_data = mem_req_data;
  assign mem_req_data = {T176, T163};
  assign T163 = {T175, T164};
  assign T164 = {T174, T165};
  assign T165 = {T173, T166};
  assign T166 = {T172, T167};
  assign T167 = {T171, T168};
  assign T168 = {T170, T169};
  assign T169 = packet_ram[3'h0];
  assign T170 = packet_ram[3'h1];
  assign T171 = packet_ram[3'h2];
  assign T172 = packet_ram[3'h3];
  assign T173 = packet_ram[3'h4];
  assign T174 = packet_ram[3'h5];
  assign T175 = packet_ram[3'h6];
  assign T176 = packet_ram[3'h7];
  assign io_mem_acquire_bits_payload_client_xact_id = acq_q_io_deq_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = acq_q_io_deq_bits_addr;
  assign io_mem_acquire_bits_header_dst = 2'h0;
  assign io_mem_acquire_bits_header_src = 2'h2;
  assign io_mem_acquire_valid = acq_q_io_deq_valid;
  assign io_cpu_0_ipi_rep_valid = R177;
  assign T344 = reset ? 1'h0 : T178;
  assign T178 = T180 ? 1'h1 : T179;
  assign T179 = io_cpu_0_ipi_rep_ready ? 1'h0 : R177;
  assign T180 = io_cpu_0_ipi_req_valid & T181;
  assign T181 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = pcr_wdata;
  assign io_cpu_0_pcr_req_bits_addr = pcr_addr;
  assign io_cpu_0_pcr_req_bits_rw = T182;
  assign T182 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T183;
  assign T183 = T185 & T184;
  assign T184 = pcr_addr != 5'h1d;
  assign T185 = T186 & T116;
  assign T186 = state == 4'h1;
  assign io_cpu_0_reset = R187;
  assign T345 = reset ? 1'h1 : T188;
  assign T188 = T190 ? T189 : R187;
  assign T189 = pcr_wdata[1'h0:1'h0];
  assign T190 = T113 & T191;
  assign T191 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T346;
  assign T346 = T192[4'hf:1'h0];
  assign T192 = tx_data >> T193;
  assign T193 = {T194, 4'h0};
  assign T194 = tx_count[1'h1:1'h0];
  assign tx_data = T334 ? tx_header : T195;
  assign T195 = T327 ? pcrReadData : T196;
  assign T196 = packet_ram[packet_ram_raddr];
  assign T197 = T118 ? T200 : T198;
  assign T198 = io_cpu_0_pcr_rep_valid ? io_cpu_0_pcr_rep_bits : T199;
  assign T199 = T113 ? T347 : pcrReadData;
  assign T347 = {63'h0, R187};
  assign T200 = T326 ? T264 : T201;
  assign T201 = T263 ? T233 : T202;
  assign T202 = T232 ? T218 : T203;
  assign T203 = T217 ? T211 : T204;
  assign T204 = T210 ? T208 : T205;
  assign T205 = T206 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T206 = T207[1'h0:1'h0];
  assign T207 = scr_addr;
  assign T208 = T209 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T209 = T207[1'h0:1'h0];
  assign T210 = T207[1'h1:1'h1];
  assign T211 = T216 ? T214 : T212;
  assign T212 = T213 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T213 = T207[1'h0:1'h0];
  assign T214 = T215 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T215 = T207[1'h0:1'h0];
  assign T216 = T207[1'h1:1'h1];
  assign T217 = T207[2'h2:2'h2];
  assign T218 = T231 ? T225 : T219;
  assign T219 = T224 ? T222 : T220;
  assign T220 = T221 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T221 = T207[1'h0:1'h0];
  assign T222 = T223 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T223 = T207[1'h0:1'h0];
  assign T224 = T207[1'h1:1'h1];
  assign T225 = T230 ? T228 : T226;
  assign T226 = T227 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T227 = T207[1'h0:1'h0];
  assign T228 = T229 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T229 = T207[1'h0:1'h0];
  assign T230 = T207[1'h1:1'h1];
  assign T231 = T207[2'h2:2'h2];
  assign T232 = T207[2'h3:2'h3];
  assign T233 = T262 ? T248 : T234;
  assign T234 = T247 ? T241 : T235;
  assign T235 = T240 ? T238 : T236;
  assign T236 = T237 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T237 = T207[1'h0:1'h0];
  assign T238 = T239 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T239 = T207[1'h0:1'h0];
  assign T240 = T207[1'h1:1'h1];
  assign T241 = T246 ? T244 : T242;
  assign T242 = T243 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T243 = T207[1'h0:1'h0];
  assign T244 = T245 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T245 = T207[1'h0:1'h0];
  assign T246 = T207[1'h1:1'h1];
  assign T247 = T207[2'h2:2'h2];
  assign T248 = T261 ? T255 : T249;
  assign T249 = T254 ? T252 : T250;
  assign T250 = T251 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T251 = T207[1'h0:1'h0];
  assign T252 = T253 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T253 = T207[1'h0:1'h0];
  assign T254 = T207[1'h1:1'h1];
  assign T255 = T260 ? T258 : T256;
  assign T256 = T257 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T257 = T207[1'h0:1'h0];
  assign T258 = T259 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T259 = T207[1'h0:1'h0];
  assign T260 = T207[1'h1:1'h1];
  assign T261 = T207[2'h2:2'h2];
  assign T262 = T207[2'h3:2'h3];
  assign T263 = T207[3'h4:3'h4];
  assign T264 = T325 ? T295 : T265;
  assign T265 = T294 ? T280 : T266;
  assign T266 = T279 ? T273 : T267;
  assign T267 = T272 ? T270 : T268;
  assign T268 = T269 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T269 = T207[1'h0:1'h0];
  assign T270 = T271 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T271 = T207[1'h0:1'h0];
  assign T272 = T207[1'h1:1'h1];
  assign T273 = T278 ? T276 : T274;
  assign T274 = T275 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T275 = T207[1'h0:1'h0];
  assign T276 = T277 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T277 = T207[1'h0:1'h0];
  assign T278 = T207[1'h1:1'h1];
  assign T279 = T207[2'h2:2'h2];
  assign T280 = T293 ? T287 : T281;
  assign T281 = T286 ? T284 : T282;
  assign T282 = T283 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T283 = T207[1'h0:1'h0];
  assign T284 = T285 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T285 = T207[1'h0:1'h0];
  assign T286 = T207[1'h1:1'h1];
  assign T287 = T292 ? T290 : T288;
  assign T288 = T289 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T289 = T207[1'h0:1'h0];
  assign T290 = T291 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T291 = T207[1'h0:1'h0];
  assign T292 = T207[1'h1:1'h1];
  assign T293 = T207[2'h2:2'h2];
  assign T294 = T207[2'h3:2'h3];
  assign T295 = T324 ? T310 : T296;
  assign T296 = T309 ? T303 : T297;
  assign T297 = T302 ? T300 : T298;
  assign T298 = T299 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T299 = T207[1'h0:1'h0];
  assign T300 = T301 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T301 = T207[1'h0:1'h0];
  assign T302 = T207[1'h1:1'h1];
  assign T303 = T308 ? T306 : T304;
  assign T304 = T305 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T305 = T207[1'h0:1'h0];
  assign T306 = T307 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T307 = T207[1'h0:1'h0];
  assign T308 = T207[1'h1:1'h1];
  assign T309 = T207[2'h2:2'h2];
  assign T310 = T323 ? T317 : T311;
  assign T311 = T316 ? T314 : T312;
  assign T312 = T313 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T313 = T207[1'h0:1'h0];
  assign T314 = T315 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T315 = T207[1'h0:1'h0];
  assign T316 = T207[1'h1:1'h1];
  assign T317 = T322 ? T320 : T318;
  assign T318 = T319 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T319 = T207[1'h0:1'h0];
  assign T320 = T321 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T321 = T207[1'h0:1'h0];
  assign T322 = T207[1'h1:1'h1];
  assign T323 = T207[2'h2:2'h2];
  assign T324 = T207[2'h3:2'h3];
  assign T325 = T207[3'h4:3'h4];
  assign T326 = T207[3'h5:3'h5];
  assign T327 = T329 | T328;
  assign T328 = cmd == 4'h3;
  assign T329 = cmd == 4'h2;
  assign tx_header = {T331, T330};
  assign T330 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T331 = {addr, seqno};
  assign T332 = T21 ? T333 : seqno;
  assign T333 = rx_shifter_in[5'h17:5'h10];
  assign T334 = tx_word_count == 13'h0;
  assign io_host_out_valid = T335;
  assign T335 = state == 4'h8;
  assign io_host_in_ready = T336;
  assign T336 = state == 4'h0;
  Queue_13 acq_q(.clk(clk), .reset(reset),
       .io_enq_ready( acq_q_io_enq_ready ),
       .io_enq_valid( T370 ),
       .io_enq_bits_addr( T364 ),
       .io_enq_bits_client_xact_id( T361 ),
       .io_enq_bits_data( T358 ),
       .io_enq_bits_uncached( T355 ),
       .io_enq_bits_a_type( T352 ),
       .io_enq_bits_subblock( T348 ),
       .io_deq_ready( io_mem_acquire_ready ),
       .io_deq_valid( acq_q_io_deq_valid ),
       .io_deq_bits_addr( acq_q_io_deq_bits_addr ),
       .io_deq_bits_client_xact_id( acq_q_io_deq_bits_client_xact_id ),
       //.io_deq_bits_data(  )
       .io_deq_bits_uncached( acq_q_io_deq_bits_uncached ),
       .io_deq_bits_a_type( acq_q_io_deq_bits_a_type ),
       .io_deq_bits_subblock( acq_q_io_deq_bits_subblock )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T21) begin
      cmd <= next_cmd;
    end
    if(T59) begin
      rx_shifter <= rx_shifter_in;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T26) begin
      rx_count <= 15'h0;
    end else if(T59) begin
      rx_count <= T25;
    end
    if(T21) begin
      size <= T29;
    end
    if(T96) begin
      addr <= T49;
    end else if(T21) begin
      addr <= T48;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T118) begin
      state <= 4'h8;
    end else if(io_cpu_0_pcr_rep_valid) begin
      state <= 4'h8;
    end else if(T113) begin
      state <= 4'h8;
    end else if(T112) begin
      state <= 4'h2;
    end else if(T102) begin
      state <= T98;
    end else if(T96) begin
      state <= T88;
    end else if(T87) begin
      state <= 4'h7;
    end else if(T81) begin
      state <= 4'h7;
    end else if(T79) begin
      state <= 4'h5;
    end else if(T77) begin
      state <= 4'h6;
    end else if(T64) begin
      state <= T15;
    end
    if(reset) begin
      mem_acked <= 1'h0;
    end else if(T85) begin
      mem_acked <= 1'h0;
    end else if(T81) begin
      mem_acked <= 1'h0;
    end else if(io_mem_grant_valid) begin
      mem_acked <= 1'h1;
    end
    if(T96) begin
      pos <= T94;
    end else if(T21) begin
      pos <= T93;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T26) begin
      tx_count <= 15'h0;
    end else if(T58) begin
      tx_count <= T57;
    end
    if (T2)
      packet_ram[3'h7] <= T1;
    if (T123)
      packet_ram[3'h6] <= T122;
    if (T127)
      packet_ram[3'h5] <= T126;
    if (T131)
      packet_ram[3'h4] <= T130;
    if (T135)
      packet_ram[3'h3] <= T134;
    if (T139)
      packet_ram[3'h2] <= T138;
    if (T143)
      packet_ram[3'h1] <= T142;
    if (T147)
      packet_ram[3'h0] <= T146;
    if (T150)
      packet_ram[T151] <= rx_shifter_in;
    if(io_mem_grant_valid) begin
      mem_gxid <= io_mem_grant_bits_payload_master_xact_id;
    end
    if(io_mem_grant_valid) begin
      mem_gsrc <= io_mem_grant_bits_header_src;
    end
    if(io_mem_grant_valid) begin
      mem_needs_ack <= T160;
    end
    if(reset) begin
      R177 <= 1'h0;
    end else if(T180) begin
      R177 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R177 <= 1'h0;
    end
    if(reset) begin
      R187 <= 1'h1;
    end else if(T190) begin
      R187 <= T189;
    end
    if(T118) begin
      pcrReadData <= T200;
    end else if(io_cpu_0_pcr_rep_valid) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T113) begin
      pcrReadData <= T347;
    end
    if(T21) begin
      seqno <= T333;
    end
  end
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [511:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [511:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [511:0] io_in_0_bits_payload_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_a_type,
    output[511:0] io_out_bits_payload_subblock,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T79;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[511:0] T10;
  wire[511:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[511:0] T23;
  wire[511:0] T24;
  wire T25;
  wire T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire T29;
  wire T30;
  wire[25:0] T31;
  wire[25:0] T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T79 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_subblock = T10;
  assign T10 = T14 ? io_in_2_bits_payload_subblock : T11;
  assign T11 = T12 ? io_in_1_bits_payload_subblock : io_in_0_bits_payload_subblock;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T15;
  assign T15 = T18 ? io_in_2_bits_payload_a_type : T16;
  assign T16 = T17 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_uncached = T19;
  assign T19 = T22 ? io_in_2_bits_payload_uncached : T20;
  assign T20 = T21 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T23;
  assign T23 = T26 ? io_in_2_bits_payload_data : T24;
  assign T24 = T25 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T27;
  assign T27 = T30 ? io_in_2_bits_payload_client_xact_id : T28;
  assign T28 = T29 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T31;
  assign T31 = T34 ? io_in_2_bits_payload_addr : T32;
  assign T32 = T33 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T35;
  assign T35 = T38 ? io_in_2_bits_header_dst : T36;
  assign T36 = T37 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T39;
  assign T39 = T42 ? io_in_2_bits_header_src : T40;
  assign T40 = T41 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T41 = T13[1'h0:1'h0];
  assign T42 = T13[1'h1:1'h1];
  assign io_out_valid = T43;
  assign T43 = T46 ? io_in_2_valid : T44;
  assign T44 = T45 ? io_in_1_valid : io_in_0_valid;
  assign T45 = T13[1'h0:1'h0];
  assign T46 = T13[1'h1:1'h1];
  assign io_in_0_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T58 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T53 | T51;
  assign T51 = io_in_2_valid & T52;
  assign T52 = last_grant < 2'h2;
  assign T53 = T56 | T54;
  assign T54 = io_in_1_valid & T55;
  assign T55 = last_grant < 2'h1;
  assign T56 = io_in_0_valid & T57;
  assign T57 = last_grant < 2'h0;
  assign T58 = last_grant < 2'h0;
  assign io_in_1_ready = T59;
  assign T59 = T60 & io_out_ready;
  assign T60 = T65 | T61;
  assign T61 = T62 ^ 1'h1;
  assign T62 = T63 | io_in_0_valid;
  assign T63 = T64 | T51;
  assign T64 = T56 | T54;
  assign T65 = T67 & T66;
  assign T66 = last_grant < 2'h1;
  assign T67 = T56 ^ 1'h1;
  assign io_in_2_ready = T68;
  assign T68 = T69 & io_out_ready;
  assign T69 = T75 | T70;
  assign T70 = T71 ^ 1'h1;
  assign T71 = T72 | io_in_1_valid;
  assign T72 = T73 | io_in_0_valid;
  assign T73 = T74 | T51;
  assign T74 = T56 | T54;
  assign T75 = T77 & T76;
  assign T76 = last_grant < 2'h2;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T56 | T54;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [511:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [511:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [511:0] io_in_0_bits_payload_subblock,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[2:0] io_out_2_bits_payload_client_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output io_out_2_bits_payload_uncached,
    output[1:0] io_out_2_bits_payload_a_type,
    output[511:0] io_out_2_bits_payload_subblock,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[2:0] io_out_1_bits_payload_client_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output io_out_1_bits_payload_uncached,
    output[1:0] io_out_1_bits_payload_a_type,
    output[511:0] io_out_1_bits_payload_subblock,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[2:0] io_out_0_bits_payload_client_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output io_out_0_bits_payload_uncached,
    output[1:0] io_out_0_bits_payload_a_type,
    output[511:0] io_out_0_bits_payload_subblock
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_0_io_in_2_ready;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire LockingRRArbiter_0_io_out_valid;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire LockingRRArbiter_0_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_subblock;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire LockingRRArbiter_1_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_subblock;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire LockingRRArbiter_2_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_subblock;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_subblock = LockingRRArbiter_0_io_out_bits_payload_subblock;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_uncached = LockingRRArbiter_0_io_out_bits_payload_uncached;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_subblock = LockingRRArbiter_1_io_out_bits_payload_subblock;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_1_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_uncached = LockingRRArbiter_1_io_out_bits_payload_uncached;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_subblock = LockingRRArbiter_2_io_out_bits_payload_subblock;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_uncached = LockingRRArbiter_2_io_out_bits_payload_uncached;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_2_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_1_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_0_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_2_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_1_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_0_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_2_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_1_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_0_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_0 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_bits_payload_subblock ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_0_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_0_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_bits_payload_subblock ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_1_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_1_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_1_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_bits_payload_subblock ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_2_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_2_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T71;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[511:0] T15;
  wire[511:0] T16;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire T21;
  wire T22;
  wire[25:0] T23;
  wire[25:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T71 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_r_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_r_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T15;
  assign T15 = T18 ? io_in_2_bits_payload_data : T16;
  assign T16 = T17 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T19;
  assign T19 = T22 ? io_in_2_bits_payload_client_xact_id : T20;
  assign T20 = T21 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T23;
  assign T23 = T26 ? io_in_2_bits_payload_addr : T24;
  assign T24 = T25 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T27;
  assign T27 = T30 ? io_in_2_bits_header_dst : T28;
  assign T28 = T29 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T31;
  assign T31 = T34 ? io_in_2_bits_header_src : T32;
  assign T32 = T33 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_valid = T35;
  assign T35 = T38 ? io_in_2_valid : T36;
  assign T36 = T37 ? io_in_1_valid : io_in_0_valid;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_in_0_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T50 | T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T45 | T43;
  assign T43 = io_in_2_valid & T44;
  assign T44 = last_grant < 2'h2;
  assign T45 = T48 | T46;
  assign T46 = io_in_1_valid & T47;
  assign T47 = last_grant < 2'h1;
  assign T48 = io_in_0_valid & T49;
  assign T49 = last_grant < 2'h0;
  assign T50 = last_grant < 2'h0;
  assign io_in_1_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T57 | T53;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T55 | io_in_0_valid;
  assign T55 = T56 | T43;
  assign T56 = T48 | T46;
  assign T57 = T59 & T58;
  assign T58 = last_grant < 2'h1;
  assign T59 = T48 ^ 1'h1;
  assign io_in_2_ready = T60;
  assign T60 = T61 & io_out_ready;
  assign T61 = T67 | T62;
  assign T62 = T63 ^ 1'h1;
  assign T63 = T64 | io_in_1_valid;
  assign T64 = T65 | io_in_0_valid;
  assign T65 = T66 | T43;
  assign T66 = T48 | T46;
  assign T67 = T69 & T68;
  assign T68 = last_grant < 2'h2;
  assign T69 = T70 ^ 1'h1;
  assign T70 = T48 | T46;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[2:0] io_out_2_bits_payload_client_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_r_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[2:0] io_out_1_bits_payload_client_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_r_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[2:0] io_out_0_bits_payload_client_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_r_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[1:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_3_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_3_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_r_type;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[1:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_4_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_4_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_r_type;
  wire LockingRRArbiter_5_io_in_2_ready;
  wire LockingRRArbiter_5_io_in_1_ready;
  wire LockingRRArbiter_5_io_in_0_ready;
  wire LockingRRArbiter_5_io_out_valid;
  wire[1:0] LockingRRArbiter_5_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_5_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_5_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_5_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_5_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_5_io_out_bits_payload_r_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_3_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_3_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_3_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_4_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_4_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_4_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_4_io_out_valid;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_5_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_5_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_5_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_5_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_5_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_5_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_5_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_5_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_4_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_3_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_5_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_4_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_3_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_5_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_4_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_3_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_1 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_3_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_3_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_3_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_3_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_4_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_4_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_4_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_4_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_5(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_5_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_5_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_5_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_5_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_5_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_5_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_5_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_5_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_5_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_5_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_p_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T63;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[25:0] T15;
  wire[25:0] T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T63 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_p_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_p_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T15;
  assign T15 = T18 ? io_in_2_bits_payload_addr : T16;
  assign T16 = T17 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T19;
  assign T19 = T22 ? io_in_2_bits_header_dst : T20;
  assign T20 = T21 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T23;
  assign T23 = T26 ? io_in_2_bits_header_src : T24;
  assign T24 = T25 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_valid = T27;
  assign T27 = T30 ? io_in_2_valid : T28;
  assign T28 = T29 ? io_in_1_valid : io_in_0_valid;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_in_0_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T42 | T33;
  assign T33 = T34 ^ 1'h1;
  assign T34 = T37 | T35;
  assign T35 = io_in_2_valid & T36;
  assign T36 = last_grant < 2'h2;
  assign T37 = T40 | T38;
  assign T38 = io_in_1_valid & T39;
  assign T39 = last_grant < 2'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = last_grant < 2'h0;
  assign T42 = last_grant < 2'h0;
  assign io_in_1_ready = T43;
  assign T43 = T44 & io_out_ready;
  assign T44 = T49 | T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 | io_in_0_valid;
  assign T47 = T48 | T35;
  assign T48 = T40 | T38;
  assign T49 = T51 & T50;
  assign T50 = last_grant < 2'h1;
  assign T51 = T40 ^ 1'h1;
  assign io_in_2_ready = T52;
  assign T52 = T53 & io_out_ready;
  assign T53 = T59 | T54;
  assign T54 = T55 ^ 1'h1;
  assign T55 = T56 | io_in_1_valid;
  assign T56 = T57 | io_in_0_valid;
  assign T57 = T58 | T35;
  assign T58 = T40 | T38;
  assign T59 = T61 & T60;
  assign T60 = last_grant < 2'h2;
  assign T61 = T62 ^ 1'h1;
  assign T62 = T40 | T38;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_6_io_in_2_ready;
  wire LockingRRArbiter_6_io_in_1_ready;
  wire LockingRRArbiter_6_io_in_0_ready;
  wire LockingRRArbiter_6_io_out_valid;
  wire[1:0] LockingRRArbiter_6_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_6_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_6_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_6_io_out_bits_payload_p_type;
  wire LockingRRArbiter_7_io_in_2_ready;
  wire LockingRRArbiter_7_io_in_1_ready;
  wire LockingRRArbiter_7_io_in_0_ready;
  wire LockingRRArbiter_7_io_out_valid;
  wire[1:0] LockingRRArbiter_7_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_7_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_7_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_7_io_out_bits_payload_p_type;
  wire LockingRRArbiter_8_io_in_2_ready;
  wire LockingRRArbiter_8_io_in_1_ready;
  wire LockingRRArbiter_8_io_in_0_ready;
  wire LockingRRArbiter_8_io_out_valid;
  wire[1:0] LockingRRArbiter_8_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_8_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_8_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_8_io_out_bits_payload_p_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_6_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_6_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_6_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_6_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_6_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_7_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_7_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_7_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_7_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_7_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_8_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_8_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_8_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_8_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_8_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_8_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_7_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_6_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_8_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_7_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_6_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_8_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_7_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_6_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_2 LockingRRArbiter_6(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_6_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_6_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_6_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_6_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_6_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_6_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_6_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( LockingRRArbiter_6_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_7(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_7_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_7_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_7_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_7_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_7_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_7_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_7_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( LockingRRArbiter_7_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_8(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_8_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_8_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_8_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_8_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_8_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_8_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_8_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( LockingRRArbiter_8_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T75;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire T25;
  wire T26;
  wire[511:0] T27;
  wire[511:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T75 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_g_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_g_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_uncached = T15;
  assign T15 = T18 ? io_in_2_bits_payload_uncached : T16;
  assign T16 = T17 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T19;
  assign T19 = T22 ? io_in_2_bits_payload_master_xact_id : T20;
  assign T20 = T21 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T23;
  assign T23 = T26 ? io_in_2_bits_payload_client_xact_id : T24;
  assign T24 = T25 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T27;
  assign T27 = T30 ? io_in_2_bits_payload_data : T28;
  assign T28 = T29 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T31;
  assign T31 = T34 ? io_in_2_bits_header_dst : T32;
  assign T32 = T33 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T35;
  assign T35 = T38 ? io_in_2_bits_header_src : T36;
  assign T36 = T37 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_out_valid = T39;
  assign T39 = T42 ? io_in_2_valid : T40;
  assign T40 = T41 ? io_in_1_valid : io_in_0_valid;
  assign T41 = T13[1'h0:1'h0];
  assign T42 = T13[1'h1:1'h1];
  assign io_in_0_ready = T43;
  assign T43 = T44 & io_out_ready;
  assign T44 = T54 | T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T49 | T47;
  assign T47 = io_in_2_valid & T48;
  assign T48 = last_grant < 2'h2;
  assign T49 = T52 | T50;
  assign T50 = io_in_1_valid & T51;
  assign T51 = last_grant < 2'h1;
  assign T52 = io_in_0_valid & T53;
  assign T53 = last_grant < 2'h0;
  assign T54 = last_grant < 2'h0;
  assign io_in_1_ready = T55;
  assign T55 = T56 & io_out_ready;
  assign T56 = T61 | T57;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T59 | io_in_0_valid;
  assign T59 = T60 | T47;
  assign T60 = T52 | T50;
  assign T61 = T63 & T62;
  assign T62 = last_grant < 2'h1;
  assign T63 = T52 ^ 1'h1;
  assign io_in_2_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T71 | T66;
  assign T66 = T67 ^ 1'h1;
  assign T67 = T68 | io_in_1_valid;
  assign T68 = T69 | io_in_0_valid;
  assign T69 = T70 | T47;
  assign T70 = T52 | T50;
  assign T71 = T73 & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T52 | T50;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output io_out_2_bits_payload_uncached,
    output[1:0] io_out_2_bits_payload_g_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output io_out_1_bits_payload_uncached,
    output[1:0] io_out_1_bits_payload_g_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output io_out_0_bits_payload_uncached,
    output[1:0] io_out_0_bits_payload_g_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_9_io_in_2_ready;
  wire LockingRRArbiter_9_io_in_1_ready;
  wire LockingRRArbiter_9_io_in_0_ready;
  wire LockingRRArbiter_9_io_out_valid;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_9_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_9_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_9_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_9_io_out_bits_payload_g_type;
  wire LockingRRArbiter_10_io_in_2_ready;
  wire LockingRRArbiter_10_io_in_1_ready;
  wire LockingRRArbiter_10_io_in_0_ready;
  wire LockingRRArbiter_10_io_out_valid;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_10_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_10_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_10_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_10_io_out_bits_payload_g_type;
  wire LockingRRArbiter_11_io_in_2_ready;
  wire LockingRRArbiter_11_io_in_1_ready;
  wire LockingRRArbiter_11_io_in_0_ready;
  wire LockingRRArbiter_11_io_out_valid;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_11_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_11_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_11_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_11_io_out_bits_payload_g_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_9_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_uncached = LockingRRArbiter_9_io_out_bits_payload_uncached;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_9_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_data = LockingRRArbiter_9_io_out_bits_payload_data;
  assign io_out_0_bits_header_dst = LockingRRArbiter_9_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_9_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_9_io_out_valid;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_10_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_uncached = LockingRRArbiter_10_io_out_bits_payload_uncached;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_10_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_data = LockingRRArbiter_10_io_out_bits_payload_data;
  assign io_out_1_bits_header_dst = LockingRRArbiter_10_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_10_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_10_io_out_valid;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_11_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_uncached = LockingRRArbiter_11_io_out_bits_payload_uncached;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_11_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_data = LockingRRArbiter_11_io_out_bits_payload_data;
  assign io_out_2_bits_header_dst = LockingRRArbiter_11_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_11_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_11_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_11_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_10_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_9_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_11_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_10_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_9_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_11_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_10_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_9_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_3 LockingRRArbiter_9(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_9_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_9_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_9_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_9_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_9_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_9_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_9_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_9_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_9_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_9_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_9_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_10(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_10_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_10_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_10_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_10_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_10_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_10_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_10_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_10_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_10_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_10_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_10_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_11(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_11_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_11_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_11_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_11_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_11_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_11_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_11_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_11_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_11_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_11_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_11_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T59;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T59 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_master_xact_id = T10;
  assign T10 = T14 ? io_in_2_bits_payload_master_xact_id : T11;
  assign T11 = T12 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T15;
  assign T15 = T18 ? io_in_2_bits_header_dst : T16;
  assign T16 = T17 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T19;
  assign T19 = T22 ? io_in_2_bits_header_src : T20;
  assign T20 = T21 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_valid = T23;
  assign T23 = T26 ? io_in_2_valid : T24;
  assign T24 = T25 ? io_in_1_valid : io_in_0_valid;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_in_0_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T38 | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T33 | T31;
  assign T31 = io_in_2_valid & T32;
  assign T32 = last_grant < 2'h2;
  assign T33 = T36 | T34;
  assign T34 = io_in_1_valid & T35;
  assign T35 = last_grant < 2'h1;
  assign T36 = io_in_0_valid & T37;
  assign T37 = last_grant < 2'h0;
  assign T38 = last_grant < 2'h0;
  assign io_in_1_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T45 | T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T43 | io_in_0_valid;
  assign T43 = T44 | T31;
  assign T44 = T36 | T34;
  assign T45 = T47 & T46;
  assign T46 = last_grant < 2'h1;
  assign T47 = T36 ^ 1'h1;
  assign io_in_2_ready = T48;
  assign T48 = T49 & io_out_ready;
  assign T49 = T55 | T50;
  assign T50 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_1_valid;
  assign T52 = T53 | io_in_0_valid;
  assign T53 = T54 | T31;
  assign T54 = T36 | T34;
  assign T55 = T57 & T56;
  assign T56 = last_grant < 2'h2;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T36 | T34;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[2:0] io_out_0_bits_payload_master_xact_id
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_12_io_in_2_ready;
  wire LockingRRArbiter_12_io_in_1_ready;
  wire LockingRRArbiter_12_io_in_0_ready;
  wire LockingRRArbiter_12_io_out_valid;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_12_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_13_io_in_2_ready;
  wire LockingRRArbiter_13_io_in_1_ready;
  wire LockingRRArbiter_13_io_in_0_ready;
  wire LockingRRArbiter_13_io_out_valid;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_13_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_14_io_in_2_ready;
  wire LockingRRArbiter_14_io_in_1_ready;
  wire LockingRRArbiter_14_io_in_0_ready;
  wire LockingRRArbiter_14_io_out_valid;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_14_io_out_bits_payload_master_xact_id;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_12_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_12_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_12_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_12_io_out_valid;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_13_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_13_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_13_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_13_io_out_valid;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_14_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_14_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_14_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_14_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_14_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_13_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_12_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_14_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_13_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_12_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_14_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_13_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_12_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_4 LockingRRArbiter_12(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_12_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_12_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_12_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_12_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_12_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_12_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_12_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_13(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_13_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_13_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_13_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_13_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_13_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_13_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_13_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_14(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_14_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_14_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_14_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_14_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_14_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_14_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_14_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketChipCrossbarNetwork(input clk, input reset,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [1:0] io_clients_1_acquire_bits_header_src,
    input [1:0] io_clients_1_acquire_bits_header_dst,
    input [25:0] io_clients_1_acquire_bits_payload_addr,
    input [2:0] io_clients_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_1_acquire_bits_payload_data,
    input  io_clients_1_acquire_bits_payload_uncached,
    input [1:0] io_clients_1_acquire_bits_payload_a_type,
    input [511:0] io_clients_1_acquire_bits_payload_subblock,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_header_src,
    output[1:0] io_clients_1_grant_bits_header_dst,
    output[511:0] io_clients_1_grant_bits_payload_data,
    output[2:0] io_clients_1_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_1_grant_bits_payload_master_xact_id,
    output io_clients_1_grant_bits_payload_uncached,
    output[1:0] io_clients_1_grant_bits_payload_g_type,
    output io_clients_1_finish_ready,
    input  io_clients_1_finish_valid,
    input [1:0] io_clients_1_finish_bits_header_src,
    input [1:0] io_clients_1_finish_bits_header_dst,
    input [2:0] io_clients_1_finish_bits_payload_master_xact_id,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[1:0] io_clients_1_probe_bits_header_src,
    output[1:0] io_clients_1_probe_bits_header_dst,
    output[25:0] io_clients_1_probe_bits_payload_addr,
    output[1:0] io_clients_1_probe_bits_payload_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_header_src,
    input [1:0] io_clients_1_release_bits_header_dst,
    input [25:0] io_clients_1_release_bits_payload_addr,
    input [2:0] io_clients_1_release_bits_payload_client_xact_id,
    input [511:0] io_clients_1_release_bits_payload_data,
    input [2:0] io_clients_1_release_bits_payload_r_type,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [1:0] io_clients_0_acquire_bits_header_src,
    input [1:0] io_clients_0_acquire_bits_header_dst,
    input [25:0] io_clients_0_acquire_bits_payload_addr,
    input [2:0] io_clients_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_0_acquire_bits_payload_data,
    input  io_clients_0_acquire_bits_payload_uncached,
    input [1:0] io_clients_0_acquire_bits_payload_a_type,
    input [511:0] io_clients_0_acquire_bits_payload_subblock,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_header_src,
    output[1:0] io_clients_0_grant_bits_header_dst,
    output[511:0] io_clients_0_grant_bits_payload_data,
    output[2:0] io_clients_0_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_0_grant_bits_payload_master_xact_id,
    output io_clients_0_grant_bits_payload_uncached,
    output[1:0] io_clients_0_grant_bits_payload_g_type,
    output io_clients_0_finish_ready,
    input  io_clients_0_finish_valid,
    input [1:0] io_clients_0_finish_bits_header_src,
    input [1:0] io_clients_0_finish_bits_header_dst,
    input [2:0] io_clients_0_finish_bits_payload_master_xact_id,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[1:0] io_clients_0_probe_bits_header_src,
    output[1:0] io_clients_0_probe_bits_header_dst,
    output[25:0] io_clients_0_probe_bits_payload_addr,
    output[1:0] io_clients_0_probe_bits_payload_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_header_src,
    input [1:0] io_clients_0_release_bits_header_dst,
    input [25:0] io_clients_0_release_bits_payload_addr,
    input [2:0] io_clients_0_release_bits_payload_client_xact_id,
    input [511:0] io_clients_0_release_bits_payload_data,
    input [2:0] io_clients_0_release_bits_payload_r_type,
    input  io_masters_0_acquire_ready,
    output io_masters_0_acquire_valid,
    output[1:0] io_masters_0_acquire_bits_header_src,
    output[1:0] io_masters_0_acquire_bits_header_dst,
    output[25:0] io_masters_0_acquire_bits_payload_addr,
    output[2:0] io_masters_0_acquire_bits_payload_client_xact_id,
    output[511:0] io_masters_0_acquire_bits_payload_data,
    output io_masters_0_acquire_bits_payload_uncached,
    output[1:0] io_masters_0_acquire_bits_payload_a_type,
    output[511:0] io_masters_0_acquire_bits_payload_subblock,
    output io_masters_0_grant_ready,
    input  io_masters_0_grant_valid,
    input [1:0] io_masters_0_grant_bits_header_src,
    input [1:0] io_masters_0_grant_bits_header_dst,
    input [511:0] io_masters_0_grant_bits_payload_data,
    input [2:0] io_masters_0_grant_bits_payload_client_xact_id,
    input [2:0] io_masters_0_grant_bits_payload_master_xact_id,
    input  io_masters_0_grant_bits_payload_uncached,
    input [1:0] io_masters_0_grant_bits_payload_g_type,
    input  io_masters_0_finish_ready,
    output io_masters_0_finish_valid,
    output[1:0] io_masters_0_finish_bits_header_src,
    output[1:0] io_masters_0_finish_bits_header_dst,
    output[2:0] io_masters_0_finish_bits_payload_master_xact_id,
    output io_masters_0_probe_ready,
    input  io_masters_0_probe_valid,
    input [1:0] io_masters_0_probe_bits_header_src,
    input [1:0] io_masters_0_probe_bits_header_dst,
    input [25:0] io_masters_0_probe_bits_payload_addr,
    input [1:0] io_masters_0_probe_bits_payload_p_type,
    input  io_masters_0_release_ready,
    output io_masters_0_release_valid,
    output[1:0] io_masters_0_release_bits_header_src,
    output[1:0] io_masters_0_release_bits_header_dst,
    output[25:0] io_masters_0_release_bits_payload_addr,
    output[2:0] io_masters_0_release_bits_payload_client_xact_id,
    output[511:0] io_masters_0_release_bits_payload_data,
    output[2:0] io_masters_0_release_bits_payload_r_type
);

  wire T61;
  wire[2:0] T62;
  wire[1:0] T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire T66;
  wire[2:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[511:0] T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire[1:0] T85;
  wire[25:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire[511:0] T93;
  wire[2:0] T94;
  wire[25:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire T99;
  wire[2:0] T100;
  wire[511:0] T101;
  wire[2:0] T102;
  wire[25:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire[511:0] T109;
  wire[1:0] T110;
  wire T111;
  wire[511:0] T112;
  wire[2:0] T113;
  wire[25:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire T118;
  wire[511:0] T119;
  wire[1:0] T120;
  wire T121;
  wire[511:0] T122;
  wire[2:0] T123;
  wire[25:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire T128;
  wire[2:0] T0;
  wire[511:0] T1;
  wire[2:0] T2;
  wire[25:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire[511:0] T15;
  wire[1:0] T16;
  wire T17;
  wire[511:0] T18;
  wire[2:0] T19;
  wire[25:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[511:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[25:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire[2:0] T53;
  wire[2:0] T54;
  wire[511:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire acqNet_io_in_2_ready;
  wire acqNet_io_in_1_ready;
  wire acqNet_io_out_0_valid;
  wire[1:0] acqNet_io_out_0_bits_header_src;
  wire[1:0] acqNet_io_out_0_bits_header_dst;
  wire[25:0] acqNet_io_out_0_bits_payload_addr;
  wire[2:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[511:0] acqNet_io_out_0_bits_payload_data;
  wire acqNet_io_out_0_bits_payload_uncached;
  wire[1:0] acqNet_io_out_0_bits_payload_a_type;
  wire[511:0] acqNet_io_out_0_bits_payload_subblock;
  wire relNet_io_in_2_ready;
  wire relNet_io_in_1_ready;
  wire relNet_io_out_0_valid;
  wire[1:0] relNet_io_out_0_bits_header_src;
  wire[1:0] relNet_io_out_0_bits_header_dst;
  wire[25:0] relNet_io_out_0_bits_payload_addr;
  wire[2:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire[511:0] relNet_io_out_0_bits_payload_data;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire prbNet_io_in_0_ready;
  wire prbNet_io_out_2_valid;
  wire[1:0] prbNet_io_out_2_bits_header_src;
  wire[1:0] prbNet_io_out_2_bits_header_dst;
  wire[25:0] prbNet_io_out_2_bits_payload_addr;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire prbNet_io_out_1_valid;
  wire[1:0] prbNet_io_out_1_bits_header_src;
  wire[1:0] prbNet_io_out_1_bits_header_dst;
  wire[25:0] prbNet_io_out_1_bits_payload_addr;
  wire[1:0] prbNet_io_out_1_bits_payload_p_type;
  wire gntNet_io_in_0_ready;
  wire gntNet_io_out_2_valid;
  wire[1:0] gntNet_io_out_2_bits_header_src;
  wire[1:0] gntNet_io_out_2_bits_header_dst;
  wire[511:0] gntNet_io_out_2_bits_payload_data;
  wire[2:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[2:0] gntNet_io_out_2_bits_payload_master_xact_id;
  wire gntNet_io_out_2_bits_payload_uncached;
  wire[1:0] gntNet_io_out_2_bits_payload_g_type;
  wire gntNet_io_out_1_valid;
  wire[1:0] gntNet_io_out_1_bits_header_src;
  wire[1:0] gntNet_io_out_1_bits_header_dst;
  wire[511:0] gntNet_io_out_1_bits_payload_data;
  wire[2:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire[2:0] gntNet_io_out_1_bits_payload_master_xact_id;
  wire gntNet_io_out_1_bits_payload_uncached;
  wire[1:0] gntNet_io_out_1_bits_payload_g_type;
  wire ackNet_io_in_2_ready;
  wire ackNet_io_in_1_ready;
  wire ackNet_io_out_0_valid;
  wire[1:0] ackNet_io_out_0_bits_header_src;
  wire[1:0] ackNet_io_out_0_bits_header_dst;
  wire[2:0] ackNet_io_out_0_bits_payload_master_xact_id;


  assign T61 = io_masters_0_finish_ready;
  assign T62 = io_clients_0_finish_bits_payload_master_xact_id;
  assign T63 = io_clients_0_finish_bits_header_dst;
  assign T64 = T65;
  assign T65 = io_clients_0_finish_bits_header_src + 2'h1;
  assign T66 = io_clients_0_finish_valid;
  assign T67 = io_clients_1_finish_bits_payload_master_xact_id;
  assign T68 = io_clients_1_finish_bits_header_dst;
  assign T69 = T70;
  assign T70 = io_clients_1_finish_bits_header_src + 2'h1;
  assign T71 = io_clients_1_finish_valid;
  assign T72 = io_clients_0_grant_ready;
  assign T73 = io_clients_1_grant_ready;
  assign T74 = io_masters_0_grant_bits_payload_g_type;
  assign T75 = io_masters_0_grant_bits_payload_uncached;
  assign T76 = io_masters_0_grant_bits_payload_master_xact_id;
  assign T77 = io_masters_0_grant_bits_payload_client_xact_id;
  assign T78 = io_masters_0_grant_bits_payload_data;
  assign T79 = T80;
  assign T80 = io_masters_0_grant_bits_header_dst + 2'h1;
  assign T81 = io_masters_0_grant_bits_header_src;
  assign T82 = io_masters_0_grant_valid;
  assign T83 = io_clients_0_probe_ready;
  assign T84 = io_clients_1_probe_ready;
  assign T85 = io_masters_0_probe_bits_payload_p_type;
  assign T86 = io_masters_0_probe_bits_payload_addr;
  assign T87 = T88;
  assign T88 = io_masters_0_probe_bits_header_dst + 2'h1;
  assign T89 = io_masters_0_probe_bits_header_src;
  assign T90 = io_masters_0_probe_valid;
  assign T91 = io_masters_0_release_ready;
  assign T92 = io_clients_0_release_bits_payload_r_type;
  assign T93 = io_clients_0_release_bits_payload_data;
  assign T94 = io_clients_0_release_bits_payload_client_xact_id;
  assign T95 = io_clients_0_release_bits_payload_addr;
  assign T96 = io_clients_0_release_bits_header_dst;
  assign T97 = T98;
  assign T98 = io_clients_0_release_bits_header_src + 2'h1;
  assign T99 = io_clients_0_release_valid;
  assign T100 = io_clients_1_release_bits_payload_r_type;
  assign T101 = io_clients_1_release_bits_payload_data;
  assign T102 = io_clients_1_release_bits_payload_client_xact_id;
  assign T103 = io_clients_1_release_bits_payload_addr;
  assign T104 = io_clients_1_release_bits_header_dst;
  assign T105 = T106;
  assign T106 = io_clients_1_release_bits_header_src + 2'h1;
  assign T107 = io_clients_1_release_valid;
  assign T108 = io_masters_0_acquire_ready;
  assign T109 = io_clients_0_acquire_bits_payload_subblock;
  assign T110 = io_clients_0_acquire_bits_payload_a_type;
  assign T111 = io_clients_0_acquire_bits_payload_uncached;
  assign T112 = io_clients_0_acquire_bits_payload_data;
  assign T113 = io_clients_0_acquire_bits_payload_client_xact_id;
  assign T114 = io_clients_0_acquire_bits_payload_addr;
  assign T115 = io_clients_0_acquire_bits_header_dst;
  assign T116 = T117;
  assign T117 = io_clients_0_acquire_bits_header_src + 2'h1;
  assign T118 = io_clients_0_acquire_valid;
  assign T119 = io_clients_1_acquire_bits_payload_subblock;
  assign T120 = io_clients_1_acquire_bits_payload_a_type;
  assign T121 = io_clients_1_acquire_bits_payload_uncached;
  assign T122 = io_clients_1_acquire_bits_payload_data;
  assign T123 = io_clients_1_acquire_bits_payload_client_xact_id;
  assign T124 = io_clients_1_acquire_bits_payload_addr;
  assign T125 = io_clients_1_acquire_bits_header_dst;
  assign T126 = T127;
  assign T127 = io_clients_1_acquire_bits_header_src + 2'h1;
  assign T128 = io_clients_1_acquire_valid;
  assign io_masters_0_release_bits_payload_r_type = T0;
  assign T0 = relNet_io_out_0_bits_payload_r_type;
  assign io_masters_0_release_bits_payload_data = T1;
  assign T1 = relNet_io_out_0_bits_payload_data;
  assign io_masters_0_release_bits_payload_client_xact_id = T2;
  assign T2 = relNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_release_bits_payload_addr = T3;
  assign T3 = relNet_io_out_0_bits_payload_addr;
  assign io_masters_0_release_bits_header_dst = T4;
  assign T4 = relNet_io_out_0_bits_header_dst;
  assign io_masters_0_release_bits_header_src = T5;
  assign T5 = T6;
  assign T6 = relNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_release_valid = T7;
  assign T7 = relNet_io_out_0_valid;
  assign io_masters_0_probe_ready = T8;
  assign T8 = prbNet_io_in_0_ready;
  assign io_masters_0_finish_bits_payload_master_xact_id = T9;
  assign T9 = ackNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_finish_bits_header_dst = T10;
  assign T10 = ackNet_io_out_0_bits_header_dst;
  assign io_masters_0_finish_bits_header_src = T11;
  assign T11 = T12;
  assign T12 = ackNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_finish_valid = T13;
  assign T13 = ackNet_io_out_0_valid;
  assign io_masters_0_grant_ready = T14;
  assign T14 = gntNet_io_in_0_ready;
  assign io_masters_0_acquire_bits_payload_subblock = T15;
  assign T15 = acqNet_io_out_0_bits_payload_subblock;
  assign io_masters_0_acquire_bits_payload_a_type = T16;
  assign T16 = acqNet_io_out_0_bits_payload_a_type;
  assign io_masters_0_acquire_bits_payload_uncached = T17;
  assign T17 = acqNet_io_out_0_bits_payload_uncached;
  assign io_masters_0_acquire_bits_payload_data = T18;
  assign T18 = acqNet_io_out_0_bits_payload_data;
  assign io_masters_0_acquire_bits_payload_client_xact_id = T19;
  assign T19 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_acquire_bits_payload_addr = T20;
  assign T20 = acqNet_io_out_0_bits_payload_addr;
  assign io_masters_0_acquire_bits_header_dst = T21;
  assign T21 = acqNet_io_out_0_bits_header_dst;
  assign io_masters_0_acquire_bits_header_src = T22;
  assign T22 = T23;
  assign T23 = acqNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_acquire_valid = T24;
  assign T24 = acqNet_io_out_0_valid;
  assign io_clients_0_release_ready = T25;
  assign T25 = relNet_io_in_1_ready;
  assign io_clients_0_probe_bits_payload_p_type = T26;
  assign T26 = prbNet_io_out_1_bits_payload_p_type;
  assign io_clients_0_probe_bits_payload_addr = T27;
  assign T27 = prbNet_io_out_1_bits_payload_addr;
  assign io_clients_0_probe_bits_header_dst = T28;
  assign T28 = T29;
  assign T29 = prbNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_probe_bits_header_src = T30;
  assign T30 = prbNet_io_out_1_bits_header_src;
  assign io_clients_0_probe_valid = T31;
  assign T31 = prbNet_io_out_1_valid;
  assign io_clients_0_finish_ready = T32;
  assign T32 = ackNet_io_in_1_ready;
  assign io_clients_0_grant_bits_payload_g_type = T33;
  assign T33 = gntNet_io_out_1_bits_payload_g_type;
  assign io_clients_0_grant_bits_payload_uncached = T34;
  assign T34 = gntNet_io_out_1_bits_payload_uncached;
  assign io_clients_0_grant_bits_payload_master_xact_id = T35;
  assign T35 = gntNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_grant_bits_payload_client_xact_id = T36;
  assign T36 = gntNet_io_out_1_bits_payload_client_xact_id;
  assign io_clients_0_grant_bits_payload_data = T37;
  assign T37 = gntNet_io_out_1_bits_payload_data;
  assign io_clients_0_grant_bits_header_dst = T38;
  assign T38 = T39;
  assign T39 = gntNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_grant_bits_header_src = T40;
  assign T40 = gntNet_io_out_1_bits_header_src;
  assign io_clients_0_grant_valid = T41;
  assign T41 = gntNet_io_out_1_valid;
  assign io_clients_0_acquire_ready = T42;
  assign T42 = acqNet_io_in_1_ready;
  assign io_clients_1_release_ready = T43;
  assign T43 = relNet_io_in_2_ready;
  assign io_clients_1_probe_bits_payload_p_type = T44;
  assign T44 = prbNet_io_out_2_bits_payload_p_type;
  assign io_clients_1_probe_bits_payload_addr = T45;
  assign T45 = prbNet_io_out_2_bits_payload_addr;
  assign io_clients_1_probe_bits_header_dst = T46;
  assign T46 = T47;
  assign T47 = prbNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_probe_bits_header_src = T48;
  assign T48 = prbNet_io_out_2_bits_header_src;
  assign io_clients_1_probe_valid = T49;
  assign T49 = prbNet_io_out_2_valid;
  assign io_clients_1_finish_ready = T50;
  assign T50 = ackNet_io_in_2_ready;
  assign io_clients_1_grant_bits_payload_g_type = T51;
  assign T51 = gntNet_io_out_2_bits_payload_g_type;
  assign io_clients_1_grant_bits_payload_uncached = T52;
  assign T52 = gntNet_io_out_2_bits_payload_uncached;
  assign io_clients_1_grant_bits_payload_master_xact_id = T53;
  assign T53 = gntNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_grant_bits_payload_client_xact_id = T54;
  assign T54 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign io_clients_1_grant_bits_payload_data = T55;
  assign T55 = gntNet_io_out_2_bits_payload_data;
  assign io_clients_1_grant_bits_header_dst = T56;
  assign T56 = T57;
  assign T57 = gntNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_grant_bits_header_src = T58;
  assign T58 = gntNet_io_out_2_bits_header_src;
  assign io_clients_1_grant_valid = T59;
  assign T59 = gntNet_io_out_2_valid;
  assign io_clients_1_acquire_ready = T60;
  assign T60 = acqNet_io_in_2_ready;
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T128 ),
       .io_in_2_bits_header_src( T126 ),
       .io_in_2_bits_header_dst( T125 ),
       .io_in_2_bits_payload_addr( T124 ),
       .io_in_2_bits_payload_client_xact_id( T123 ),
       .io_in_2_bits_payload_data( T122 ),
       .io_in_2_bits_payload_uncached( T121 ),
       .io_in_2_bits_payload_a_type( T120 ),
       .io_in_2_bits_payload_subblock( T119 ),
       .io_in_1_ready( acqNet_io_in_1_ready ),
       .io_in_1_valid( T118 ),
       .io_in_1_bits_header_src( T116 ),
       .io_in_1_bits_header_dst( T115 ),
       .io_in_1_bits_payload_addr( T114 ),
       .io_in_1_bits_payload_client_xact_id( T113 ),
       .io_in_1_bits_payload_data( T112 ),
       .io_in_1_bits_payload_uncached( T111 ),
       .io_in_1_bits_payload_a_type( T110 ),
       .io_in_1_bits_payload_subblock( T109 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_uncached(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_subblock(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_uncached(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_subblock(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_uncached(  )
       //.io_out_1_bits_payload_a_type(  )
       //.io_out_1_bits_payload_subblock(  )
       .io_out_0_ready( T108 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( acqNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_uncached( acqNet_io_out_0_bits_payload_uncached ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_subblock( acqNet_io_out_0_bits_payload_subblock )
  );
  `ifndef SYNTHESIS
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {16{$random}};
    assign acqNet.io_in_0_bits_payload_uncached = {1{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_subblock = {16{$random}};
  `endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T107 ),
       .io_in_2_bits_header_src( T105 ),
       .io_in_2_bits_header_dst( T104 ),
       .io_in_2_bits_payload_addr( T103 ),
       .io_in_2_bits_payload_client_xact_id( T102 ),
       .io_in_2_bits_payload_data( T101 ),
       .io_in_2_bits_payload_r_type( T100 ),
       .io_in_1_ready( relNet_io_in_1_ready ),
       .io_in_1_valid( T99 ),
       .io_in_1_bits_header_src( T97 ),
       .io_in_1_bits_header_dst( T96 ),
       .io_in_1_bits_payload_addr( T95 ),
       .io_in_1_bits_payload_client_xact_id( T94 ),
       .io_in_1_bits_payload_data( T93 ),
       .io_in_1_bits_payload_r_type( T92 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_r_type(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_r_type(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_r_type(  )
       .io_out_0_ready( T91 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( relNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type )
  );
  `ifndef SYNTHESIS
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {16{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
  `endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr(  )
       //.io_in_2_bits_payload_p_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr(  )
       //.io_in_1_bits_payload_p_type(  )
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T90 ),
       .io_in_0_bits_header_src( T89 ),
       .io_in_0_bits_header_dst( T87 ),
       .io_in_0_bits_payload_addr( T86 ),
       .io_in_0_bits_payload_p_type( T85 ),
       .io_out_2_ready( T84 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr( prbNet_io_out_2_bits_payload_addr ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( T83 ),
       .io_out_1_valid( prbNet_io_out_1_valid ),
       .io_out_1_bits_header_src( prbNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( prbNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr( prbNet_io_out_1_bits_payload_addr ),
       .io_out_1_bits_payload_p_type( prbNet_io_out_1_bits_payload_p_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr(  )
       //.io_out_0_bits_payload_p_type(  )
  );
  `ifndef SYNTHESIS
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_1_bits_header_src = {1{$random}};
    assign prbNet.io_in_1_bits_header_dst = {1{$random}};
    assign prbNet.io_in_1_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_1_bits_payload_p_type = {1{$random}};
  `endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_data(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_uncached(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_uncached(  )
       //.io_in_1_bits_payload_g_type(  )
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T82 ),
       .io_in_0_bits_header_src( T81 ),
       .io_in_0_bits_header_dst( T79 ),
       .io_in_0_bits_payload_data( T78 ),
       .io_in_0_bits_payload_client_xact_id( T77 ),
       .io_in_0_bits_payload_master_xact_id( T76 ),
       .io_in_0_bits_payload_uncached( T75 ),
       .io_in_0_bits_payload_g_type( T74 ),
       .io_out_2_ready( T73 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_master_xact_id( gntNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_uncached( gntNet_io_out_2_bits_payload_uncached ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_1_ready( T72 ),
       .io_out_1_valid( gntNet_io_out_1_valid ),
       .io_out_1_bits_header_src( gntNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( gntNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_data( gntNet_io_out_1_bits_payload_data ),
       .io_out_1_bits_payload_client_xact_id( gntNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_master_xact_id( gntNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_uncached( gntNet_io_out_1_bits_payload_uncached ),
       .io_out_1_bits_payload_g_type( gntNet_io_out_1_bits_payload_g_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_data(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_uncached(  )
       //.io_out_0_bits_payload_g_type(  )
  );
  `ifndef SYNTHESIS
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {16{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_uncached = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_1_bits_header_src = {1{$random}};
    assign gntNet.io_in_1_bits_header_dst = {1{$random}};
    assign gntNet.io_in_1_bits_payload_data = {16{$random}};
    assign gntNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_uncached = {1{$random}};
    assign gntNet.io_in_1_bits_payload_g_type = {1{$random}};
  `endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T71 ),
       .io_in_2_bits_header_src( T69 ),
       .io_in_2_bits_header_dst( T68 ),
       .io_in_2_bits_payload_master_xact_id( T67 ),
       .io_in_1_ready( ackNet_io_in_1_ready ),
       .io_in_1_valid( T66 ),
       .io_in_1_bits_header_src( T64 ),
       .io_in_1_bits_header_dst( T63 ),
       .io_in_1_bits_payload_master_xact_id( T62 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       .io_out_0_ready( T61 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_master_xact_id( ackNet_io_out_0_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module VoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[1:0] io_inner_probe_bits_header_src
    //output[1:0] io_inner_probe_bits_header_dst
    //output[25:0] io_inner_probe_bits_payload_addr
    //output[1:0] io_inner_probe_bits_payload_p_type
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T35;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [25:0] xact_addr;
  wire[25:0] T20;
  wire[7:0] T21;
  wire[1:0] T22;
  wire T23;
  wire[2:0] T24;
  reg [2:0] xact_data;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[1:0] T36;
  reg  init_client_id;
  wire T37;
  wire[1:0] T38;
  wire[1:0] T34;
  wire[1:0] T39;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T19 & T1;
  assign T1 = state != 2'h0;
  assign T35 = reset ? 2'h0 : T2;
  assign T2 = T17 ? 2'h0 : T3;
  assign T3 = T15 ? 2'h2 : T4;
  assign T4 = T13 ? T5 : state;
  assign T5 = T6 ? 2'h1 : 2'h2;
  assign T6 = T8 | T7;
  assign T7 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T8 = T10 | T9;
  assign T9 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T10 = T12 | T11;
  assign T11 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T12 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T13 = T14 & io_inner_release_valid;
  assign T14 = 2'h0 == state;
  assign T15 = T16 & io_outer_acquire_ready;
  assign T16 = 2'h1 == state;
  assign T17 = T18 & io_inner_grant_ready;
  assign T18 = 2'h2 == state;
  assign T19 = xact_addr == io_inner_release_bits_payload_addr;
  assign T20 = T13 ? io_inner_release_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = 1'h0;
  assign io_outer_acquire_bits_payload_subblock = T21;
  assign T21 = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T22;
  assign T22 = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T23;
  assign T23 = 1'h1;
  assign io_outer_acquire_bits_payload_data = T24;
  assign T24 = xact_data;
  assign T25 = T13 ? io_inner_release_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T26;
  assign T26 = 3'h0;
  assign io_outer_acquire_bits_payload_addr = T27;
  assign T27 = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T16;
  assign io_inner_release_ready = T13;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_grant_bits_payload_g_type = T28;
  assign T28 = 2'h0;
  assign io_inner_grant_bits_payload_uncached = T29;
  assign T29 = 1'h0;
  assign io_inner_grant_bits_payload_master_xact_id = T30;
  assign T30 = 3'h0;
  assign io_inner_grant_bits_payload_client_xact_id = T31;
  assign T31 = xact_client_xact_id;
  assign T32 = T13 ? io_inner_release_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T33;
  assign T33 = 3'h0;
  assign io_inner_grant_bits_header_dst = T36;
  assign T36 = {1'h0, init_client_id};
  assign T37 = T38[1'h0:1'h0];
  assign T38 = reset ? 2'h0 : T34;
  assign T34 = T13 ? io_inner_release_bits_header_src : T39;
  assign T39 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T18;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T17) begin
      state <= 2'h0;
    end else if(T15) begin
      state <= 2'h2;
    end else if(T13) begin
      state <= T5;
    end
    if(T13) begin
      xact_addr <= io_inner_release_bits_payload_addr;
    end
    if(T13) begin
      xact_data <= io_inner_release_bits_payload_data;
    end
    if(T13) begin
      xact_client_xact_id <= io_inner_release_bits_payload_client_xact_id;
    end
    init_client_id <= T37;
  end
endmodule

module AcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h1;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h1;
  assign outer_read_client_xact_id = 3'h1;
  assign outer_write_acq_client_xact_id = 3'h1;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h1;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h1;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module AcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h2;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h2;
  assign outer_read_client_xact_id = 3'h2;
  assign outer_write_acq_client_xact_id = 3'h2;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h2;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h2;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module AcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h3;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h3;
  assign outer_read_client_xact_id = 3'h3;
  assign outer_write_acq_client_xact_id = 3'h3;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h3;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h3;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module AcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h4;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h4;
  assign outer_read_client_xact_id = 3'h4;
  assign outer_write_acq_client_xact_id = 3'h4;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h4;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h4;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module AcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h5;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h5;
  assign outer_read_client_xact_id = 3'h5;
  assign outer_write_acq_client_xact_id = 3'h5;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h5;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h5;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module AcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h6;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h6;
  assign outer_read_client_xact_id = 3'h6;
  assign outer_write_acq_client_xact_id = 3'h6;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h6;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h6;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module AcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [2:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [7:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[2:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[2:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[7:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [2:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T142;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  wire T25;
  reg [1:0] xact_a_type;
  wire[1:0] T26;
  reg  xact_uncached;
  wire T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  release_count;
  wire T143;
  wire[1:0] T144;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T145;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T146;
  wire T39;
  wire[1:0] T147;
  wire T40;
  wire[1:0] T148;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg [25:0] xact_addr;
  wire[25:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] outer_write_rel_subblock;
  wire[7:0] outer_read_subblock;
  wire[7:0] outer_write_acq_subblock;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T87;
  wire T88;
  wire T89;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] outer_write_rel_data;
  wire[2:0] outer_read_data;
  wire[2:0] outer_write_acq_data;
  reg [2:0] xact_data;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T97;
  wire[25:0] T98;
  wire[25:0] T99;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[25:0] T113;
  wire[1:0] T149;
  wire T150;
  wire T151;
  reg [1:0] probe_flags;
  wire[1:0] T152;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  reg [2:0] xact_client_xact_id;
  wire[2:0] T135;
  wire[2:0] T136;
  wire[1:0] T153;
  reg  init_client_id;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T137;
  wire[1:0] T156;
  wire T138;
  wire T139;
  wire T140;
  wire T141;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_uncached = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T76 & T1;
  assign T1 = state != 3'h0;
  assign T142 = reset ? 3'h0 : T2;
  assign T2 = T72 ? 3'h0 : T3;
  assign T3 = T70 ? T67 : T4;
  assign T4 = T65 ? T64 : T5;
  assign T5 = T62 ? T59 : T6;
  assign T6 = T57 ? T55 : T7;
  assign T7 = T31 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T25 : 1'h1;
  assign T25 = xact_a_type != 2'h1;
  assign T26 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign T27 = T21 ? io_inner_acquire_bits_payload_uncached : xact_uncached;
  assign pending_outer_write = xact_uncached ? T28 : 1'h0;
  assign T28 = T30 | T29;
  assign T29 = 2'h2 == xact_a_type;
  assign T30 = 2'h1 == xact_a_type;
  assign T31 = T53 & T32;
  assign T32 = release_count == 1'h1;
  assign T143 = T144[1'h0:1'h0];
  assign T144 = reset ? 2'h0 : T33;
  assign T33 = T42 ? T148 : T34;
  assign T34 = T53 ? T147 : T35;
  assign T35 = T21 ? T36 : T145;
  assign T145 = {1'h0, release_count};
  assign T36 = T146 + T37;
  assign T37 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h1:1'h1];
  assign T146 = {1'h0, T39};
  assign T39 = probe_initial_flags[1'h0:1'h0];
  assign T147 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T148 = {1'h0, T41};
  assign T41 = release_count - 1'h1;
  assign T42 = T51 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T50 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T51 = T52 & io_inner_release_valid;
  assign T52 = 3'h1 == state;
  assign T53 = T54 & io_outer_acquire_ready;
  assign T54 = T51 & T44;
  assign T55 = pending_outer_write ? 3'h3 : T56;
  assign T56 = pending_outer_read ? 3'h2 : 3'h4;
  assign T57 = T42 & T58;
  assign T58 = release_count == 1'h1;
  assign T59 = T60 ? 3'h5 : 3'h0;
  assign T60 = io_inner_grant_bits_payload_uncached | T61;
  assign T61 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T62 = T63 & io_outer_acquire_ready;
  assign T63 = 3'h2 == state;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign T65 = T66 & io_outer_acquire_ready;
  assign T66 = 3'h3 == state;
  assign T67 = T68 ? 3'h5 : 3'h0;
  assign T68 = io_inner_grant_bits_payload_uncached | T69;
  assign T69 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T70 = T71 & io_inner_grant_ready;
  assign T71 = 3'h4 == state;
  assign T72 = T75 & T73;
  assign T73 = io_inner_finish_valid & T74;
  assign T74 = io_inner_finish_bits_payload_master_xact_id == 3'h7;
  assign T75 = 3'h5 == state;
  assign T76 = xact_addr == io_inner_release_bits_payload_addr;
  assign T77 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T78;
  assign T78 = T80 & T79;
  assign T79 = state != 3'h0;
  assign T80 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T81;
  assign T81 = T66 ? outer_write_acq_subblock : T82;
  assign T82 = T63 ? outer_read_subblock : T83;
  assign T83 = T54 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 8'hff;
  assign outer_read_subblock = 8'h7;
  assign outer_write_acq_subblock = 8'hff;
  assign io_outer_acquire_bits_payload_a_type = T84;
  assign T84 = T66 ? outer_write_acq_a_type : T85;
  assign T85 = T63 ? outer_read_a_type : T86;
  assign T86 = T54 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T87;
  assign T87 = T66 ? outer_write_acq_uncached : T88;
  assign T88 = T63 ? outer_read_uncached : T89;
  assign T89 = T54 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T90;
  assign T90 = T66 ? outer_write_acq_data : T91;
  assign T91 = T63 ? outer_read_data : T92;
  assign T92 = T54 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = 3'h0;
  assign outer_read_data = 3'h0;
  assign outer_write_acq_data = xact_data;
  assign T93 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T94;
  assign T94 = T66 ? outer_write_acq_client_xact_id : T95;
  assign T95 = T63 ? outer_read_client_xact_id : T96;
  assign T96 = T54 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h7;
  assign outer_read_client_xact_id = 3'h7;
  assign outer_write_acq_client_xact_id = 3'h7;
  assign io_outer_acquire_bits_payload_addr = T97;
  assign T97 = T66 ? outer_write_acq_addr : T98;
  assign T98 = T63 ? outer_read_addr : T99;
  assign T99 = T54 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T100;
  assign T100 = T66 ? 1'h1 : T101;
  assign T101 = T63 ? 1'h1 : T54;
  assign io_inner_release_ready = T102;
  assign T102 = T42 ? 1'h1 : T53;
  assign io_inner_probe_bits_payload_p_type = T103;
  assign T103 = T104;
  assign T104 = xact_uncached ? T107 : T105;
  assign T105 = T106 ? 2'h1 : 2'h0;
  assign T106 = xact_a_type == 2'h0;
  assign T107 = T112 ? 2'h2 : T108;
  assign T108 = T111 ? 2'h0 : T109;
  assign T109 = T110 ? 2'h0 : 2'h2;
  assign T110 = xact_a_type == 2'h2;
  assign T111 = xact_a_type == 2'h1;
  assign T112 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T113;
  assign T113 = xact_addr;
  assign io_inner_probe_bits_header_dst = T149;
  assign T149 = {1'h0, T150};
  assign T150 = T151 == 1'h0;
  assign T151 = probe_flags[1'h0:1'h0];
  assign T152 = reset ? 2'h0 : T114;
  assign T114 = T119 ? T116 : T115;
  assign T115 = T21 ? probe_initial_flags : probe_flags;
  assign T116 = probe_flags & T117;
  assign T117 = ~ T118;
  assign T118 = 1'h1 << T150;
  assign T119 = T52 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T120;
  assign T120 = T52 ? T121 : 1'h0;
  assign T121 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T122;
  assign T122 = T123;
  assign T123 = xact_uncached ? T126 : T124;
  assign T124 = T125 ? 2'h1 : 2'h2;
  assign T125 = xact_a_type == 2'h0;
  assign T126 = T131 ? 2'h0 : T127;
  assign T127 = T130 ? 2'h1 : T128;
  assign T128 = T129 ? 2'h2 : 2'h0;
  assign T129 = xact_a_type == 2'h2;
  assign T130 = xact_a_type == 2'h1;
  assign T131 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T132;
  assign T132 = xact_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = T133;
  assign T133 = 3'h7;
  assign io_inner_grant_bits_payload_client_xact_id = T134;
  assign T134 = xact_client_xact_id;
  assign T135 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T136;
  assign T136 = 3'h0;
  assign io_inner_grant_bits_header_dst = T153;
  assign T153 = {1'h0, init_client_id};
  assign T154 = T155[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T137;
  assign T137 = T21 ? io_inner_acquire_bits_header_src : T156;
  assign T156 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T138;
  assign T138 = T139 ? 1'h1 : T71;
  assign T139 = T75 & T140;
  assign T140 = io_outer_grant_valid & T141;
  assign T141 = io_outer_grant_bits_payload_client_xact_id == 3'h7;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T72) begin
      state <= 3'h0;
    end else if(T70) begin
      state <= T67;
    end else if(T65) begin
      state <= T64;
    end else if(T62) begin
      state <= T59;
    end else if(T57) begin
      state <= T55;
    end else if(T31) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    if(T21) begin
      xact_uncached <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T143;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T119) begin
      probe_flags <= T116;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T154;
  end
endmodule

module Arbiter_12(
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits : io_in_0_bits;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits : io_in_2_bits;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits : io_in_4_bits;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits : io_in_6_bits;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_valid = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_valid : io_in_0_valid;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_valid : io_in_4_valid;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_valid : io_in_6_valid;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T41 ^ 1'h1;
  assign T41 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T45 | io_in_2_valid;
  assign T45 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T46;
  assign T46 = T47 & io_out_ready;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T49 | io_in_3_valid;
  assign T49 = T50 | io_in_2_valid;
  assign T50 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T54 | io_in_4_valid;
  assign T54 = T55 | io_in_3_valid;
  assign T55 = T56 | io_in_2_valid;
  assign T56 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_5_valid;
  assign T60 = T61 | io_in_4_valid;
  assign T61 = T62 | io_in_3_valid;
  assign T62 = T63 | io_in_2_valid;
  assign T63 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_6_valid;
  assign T67 = T68 | io_in_5_valid;
  assign T68 = T69 | io_in_4_valid;
  assign T69 = T70 | io_in_3_valid;
  assign T70 = T71 | io_in_2_valid;
  assign T71 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_13(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [1:0] io_in_7_bits_payload_p_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [1:0] io_in_6_bits_payload_p_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [1:0] io_in_5_bits_payload_p_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[25:0] T23;
  wire[25:0] T24;
  wire[25:0] T25;
  wire T26;
  wire[25:0] T27;
  wire T28;
  wire T29;
  wire[25:0] T30;
  wire[25:0] T31;
  wire T32;
  wire[25:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_p_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_p_type : io_in_4_bits_payload_p_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_p_type : io_in_6_bits_payload_p_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_addr = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_valid = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_valid : io_in_0_valid;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_valid : io_in_2_valid;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_valid : io_in_4_valid;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_valid : io_in_6_valid;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T79;
  assign T79 = T80 & io_out_ready;
  assign T80 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T81;
  assign T81 = T82 & io_out_ready;
  assign T82 = T83 ^ 1'h1;
  assign T83 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T84;
  assign T84 = T85 & io_out_ready;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T87 | io_in_2_valid;
  assign T87 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T88;
  assign T88 = T89 & io_out_ready;
  assign T89 = T90 ^ 1'h1;
  assign T90 = T91 | io_in_3_valid;
  assign T91 = T92 | io_in_2_valid;
  assign T92 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = T95 ^ 1'h1;
  assign T95 = T96 | io_in_4_valid;
  assign T96 = T97 | io_in_3_valid;
  assign T97 = T98 | io_in_2_valid;
  assign T98 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T99;
  assign T99 = T100 & io_out_ready;
  assign T100 = T101 ^ 1'h1;
  assign T101 = T102 | io_in_5_valid;
  assign T102 = T103 | io_in_4_valid;
  assign T103 = T104 | io_in_3_valid;
  assign T104 = T105 | io_in_2_valid;
  assign T105 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T106;
  assign T106 = T107 & io_out_ready;
  assign T107 = T108 ^ 1'h1;
  assign T108 = T109 | io_in_6_valid;
  assign T109 = T110 | io_in_5_valid;
  assign T110 = T111 | io_in_4_valid;
  assign T111 = T112 | io_in_3_valid;
  assign T112 = T113 | io_in_2_valid;
  assign T113 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_14(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [511:0] io_in_7_bits_payload_data,
    input [2:0] io_in_7_bits_payload_client_xact_id,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input  io_in_7_bits_payload_uncached,
    input [1:0] io_in_7_bits_payload_g_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [511:0] io_in_6_bits_payload_data,
    input [2:0] io_in_6_bits_payload_client_xact_id,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input  io_in_6_bits_payload_uncached,
    input [1:0] io_in_6_bits_payload_g_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [511:0] io_in_5_bits_payload_data,
    input [2:0] io_in_5_bits_payload_client_xact_id,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input  io_in_5_bits_payload_uncached,
    input [1:0] io_in_5_bits_payload_g_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [511:0] io_in_4_bits_payload_data,
    input [2:0] io_in_4_bits_payload_client_xact_id,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input  io_in_4_bits_payload_uncached,
    input [1:0] io_in_4_bits_payload_g_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [511:0] io_in_3_bits_payload_data,
    input [2:0] io_in_3_bits_payload_client_xact_id,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input  io_in_3_bits_payload_uncached,
    input [1:0] io_in_3_bits_payload_g_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire[2:0] T39;
  wire T40;
  wire[2:0] T41;
  wire T42;
  wire T43;
  wire[2:0] T44;
  wire[2:0] T45;
  wire T46;
  wire[2:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire[2:0] T53;
  wire T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire T60;
  wire[2:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[511:0] T65;
  wire[511:0] T66;
  wire[511:0] T67;
  wire T68;
  wire[511:0] T69;
  wire T70;
  wire T71;
  wire[511:0] T72;
  wire[511:0] T73;
  wire T74;
  wire[511:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire[1:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire[1:0] T97;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_g_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_g_type : io_in_4_bits_payload_g_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_g_type : io_in_6_bits_payload_g_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_uncached = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_uncached : io_in_2_bits_payload_uncached;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_uncached : io_in_4_bits_payload_uncached;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_uncached : io_in_6_bits_payload_uncached;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_payload_data = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T93;
  assign T93 = T106 ? T100 : T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T96 = T12[1'h0:1'h0];
  assign T97 = T98 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T98 = T12[1'h0:1'h0];
  assign T99 = T12[1'h1:1'h1];
  assign T100 = T105 ? T103 : T101;
  assign T101 = T102 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T102 = T12[1'h0:1'h0];
  assign T103 = T104 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T104 = T12[1'h0:1'h0];
  assign T105 = T12[1'h1:1'h1];
  assign T106 = T12[2'h2:2'h2];
  assign io_out_valid = T107;
  assign T107 = T120 ? T114 : T108;
  assign T108 = T113 ? T111 : T109;
  assign T109 = T110 ? io_in_1_valid : io_in_0_valid;
  assign T110 = T12[1'h0:1'h0];
  assign T111 = T112 ? io_in_3_valid : io_in_2_valid;
  assign T112 = T12[1'h0:1'h0];
  assign T113 = T12[1'h1:1'h1];
  assign T114 = T119 ? T117 : T115;
  assign T115 = T116 ? io_in_5_valid : io_in_4_valid;
  assign T116 = T12[1'h0:1'h0];
  assign T117 = T118 ? io_in_7_valid : io_in_6_valid;
  assign T118 = T12[1'h0:1'h0];
  assign T119 = T12[1'h1:1'h1];
  assign T120 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T121;
  assign T121 = T122 & io_out_ready;
  assign T122 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T123;
  assign T123 = T124 & io_out_ready;
  assign T124 = T125 ^ 1'h1;
  assign T125 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T126;
  assign T126 = T127 & io_out_ready;
  assign T127 = T128 ^ 1'h1;
  assign T128 = T129 | io_in_2_valid;
  assign T129 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T130;
  assign T130 = T131 & io_out_ready;
  assign T131 = T132 ^ 1'h1;
  assign T132 = T133 | io_in_3_valid;
  assign T133 = T134 | io_in_2_valid;
  assign T134 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T135;
  assign T135 = T136 & io_out_ready;
  assign T136 = T137 ^ 1'h1;
  assign T137 = T138 | io_in_4_valid;
  assign T138 = T139 | io_in_3_valid;
  assign T139 = T140 | io_in_2_valid;
  assign T140 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T141;
  assign T141 = T142 & io_out_ready;
  assign T142 = T143 ^ 1'h1;
  assign T143 = T144 | io_in_5_valid;
  assign T144 = T145 | io_in_4_valid;
  assign T145 = T146 | io_in_3_valid;
  assign T146 = T147 | io_in_2_valid;
  assign T147 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T148;
  assign T148 = T149 & io_out_ready;
  assign T149 = T150 ^ 1'h1;
  assign T150 = T151 | io_in_6_valid;
  assign T151 = T152 | io_in_5_valid;
  assign T152 = T153 | io_in_4_valid;
  assign T153 = T154 | io_in_3_valid;
  assign T154 = T155 | io_in_2_valid;
  assign T155 = io_in_0_valid | io_in_1_valid;
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [2:0] io_in_7_bits_payload_client_xact_id,
    input [2:0] io_in_7_bits_payload_data,
    input  io_in_7_bits_payload_uncached,
    input [1:0] io_in_7_bits_payload_a_type,
    input [7:0] io_in_7_bits_payload_subblock,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [2:0] io_in_6_bits_payload_client_xact_id,
    input [2:0] io_in_6_bits_payload_data,
    input  io_in_6_bits_payload_uncached,
    input [1:0] io_in_6_bits_payload_a_type,
    input [7:0] io_in_6_bits_payload_subblock,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [2:0] io_in_5_bits_payload_client_xact_id,
    input [2:0] io_in_5_bits_payload_data,
    input  io_in_5_bits_payload_uncached,
    input [1:0] io_in_5_bits_payload_a_type,
    input [7:0] io_in_5_bits_payload_subblock,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [2:0] io_in_4_bits_payload_client_xact_id,
    input [2:0] io_in_4_bits_payload_data,
    input  io_in_4_bits_payload_uncached,
    input [1:0] io_in_4_bits_payload_a_type,
    input [7:0] io_in_4_bits_payload_subblock,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [2:0] io_in_3_bits_payload_client_xact_id,
    input [2:0] io_in_3_bits_payload_data,
    input  io_in_3_bits_payload_uncached,
    input [1:0] io_in_3_bits_payload_a_type,
    input [7:0] io_in_3_bits_payload_subblock,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [7:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [7:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [7:0] io_in_0_bits_payload_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_data,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_a_type,
    output[7:0] io_out_bits_payload_subblock,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T326;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire T78;
  wire[2:0] T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[2:0] T83;
  wire T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire[2:0] T90;
  wire[2:0] T91;
  wire T92;
  wire[2:0] T93;
  wire T94;
  wire T95;
  wire[2:0] T96;
  wire[2:0] T97;
  wire T98;
  wire[2:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[25:0] T103;
  wire[25:0] T104;
  wire[25:0] T105;
  wire T106;
  wire[25:0] T107;
  wire T108;
  wire T109;
  wire[25:0] T110;
  wire[25:0] T111;
  wire T112;
  wire[25:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire T120;
  wire[1:0] T121;
  wire T122;
  wire T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire T126;
  wire[1:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire T140;
  wire[1:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T30 ? 3'h1 : T2;
  assign T2 = T28 ? 3'h2 : T3;
  assign T3 = T26 ? 3'h3 : T4;
  assign T4 = T24 ? 3'h4 : T5;
  assign T5 = T22 ? 3'h5 : T6;
  assign T6 = T20 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T326 = reset ? 3'h0 : T18;
  assign T18 = T19 ? T0 : R17;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = io_in_6_valid & T21;
  assign T21 = R17 < 3'h6;
  assign T22 = io_in_5_valid & T23;
  assign T23 = R17 < 3'h5;
  assign T24 = io_in_4_valid & T25;
  assign T25 = R17 < 3'h4;
  assign T26 = io_in_3_valid & T27;
  assign T27 = R17 < 3'h3;
  assign T28 = io_in_2_valid & T29;
  assign T29 = R17 < 3'h2;
  assign T30 = io_in_1_valid & T31;
  assign T31 = R17 < 3'h1;
  assign io_out_bits_payload_subblock = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_payload_subblock : io_in_0_bits_payload_subblock;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = T0;
  assign T37 = T38 ? io_in_3_bits_payload_subblock : io_in_2_bits_payload_subblock;
  assign T38 = T36[1'h0:1'h0];
  assign T39 = T36[1'h1:1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_payload_subblock : io_in_4_bits_payload_subblock;
  assign T42 = T36[1'h0:1'h0];
  assign T43 = T44 ? io_in_7_bits_payload_subblock : io_in_6_bits_payload_subblock;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign T46 = T36[2'h2:2'h2];
  assign io_out_bits_payload_a_type = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T50 = T36[1'h0:1'h0];
  assign T51 = T52 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_payload_a_type : io_in_4_bits_payload_a_type;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T58 ? io_in_7_bits_payload_a_type : io_in_6_bits_payload_a_type;
  assign T58 = T36[1'h0:1'h0];
  assign T59 = T36[1'h1:1'h1];
  assign T60 = T36[2'h2:2'h2];
  assign io_out_bits_payload_uncached = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T66 ? io_in_3_bits_payload_uncached : io_in_2_bits_payload_uncached;
  assign T66 = T36[1'h0:1'h0];
  assign T67 = T36[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_payload_uncached : io_in_4_bits_payload_uncached;
  assign T70 = T36[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_payload_uncached : io_in_6_bits_payload_uncached;
  assign T72 = T36[1'h0:1'h0];
  assign T73 = T36[1'h1:1'h1];
  assign T74 = T36[2'h2:2'h2];
  assign io_out_bits_payload_data = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T78 = T36[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T80 = T36[1'h0:1'h0];
  assign T81 = T36[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T84 = T36[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T86 = T36[1'h0:1'h0];
  assign T87 = T36[1'h1:1'h1];
  assign T88 = T36[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T89;
  assign T89 = T102 ? T96 : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T92 = T36[1'h0:1'h0];
  assign T93 = T94 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T94 = T36[1'h0:1'h0];
  assign T95 = T36[1'h1:1'h1];
  assign T96 = T101 ? T99 : T97;
  assign T97 = T98 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T98 = T36[1'h0:1'h0];
  assign T99 = T100 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T100 = T36[1'h0:1'h0];
  assign T101 = T36[1'h1:1'h1];
  assign T102 = T36[2'h2:2'h2];
  assign io_out_bits_payload_addr = T103;
  assign T103 = T116 ? T110 : T104;
  assign T104 = T109 ? T107 : T105;
  assign T105 = T106 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T106 = T36[1'h0:1'h0];
  assign T107 = T108 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T108 = T36[1'h0:1'h0];
  assign T109 = T36[1'h1:1'h1];
  assign T110 = T115 ? T113 : T111;
  assign T111 = T112 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T112 = T36[1'h0:1'h0];
  assign T113 = T114 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T114 = T36[1'h0:1'h0];
  assign T115 = T36[1'h1:1'h1];
  assign T116 = T36[2'h2:2'h2];
  assign io_out_bits_header_dst = T117;
  assign T117 = T130 ? T124 : T118;
  assign T118 = T123 ? T121 : T119;
  assign T119 = T120 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T120 = T36[1'h0:1'h0];
  assign T121 = T122 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T122 = T36[1'h0:1'h0];
  assign T123 = T36[1'h1:1'h1];
  assign T124 = T129 ? T127 : T125;
  assign T125 = T126 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T126 = T36[1'h0:1'h0];
  assign T127 = T128 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T128 = T36[1'h0:1'h0];
  assign T129 = T36[1'h1:1'h1];
  assign T130 = T36[2'h2:2'h2];
  assign io_out_bits_header_src = T131;
  assign T131 = T144 ? T138 : T132;
  assign T132 = T137 ? T135 : T133;
  assign T133 = T134 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T134 = T36[1'h0:1'h0];
  assign T135 = T136 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T136 = T36[1'h0:1'h0];
  assign T137 = T36[1'h1:1'h1];
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T140 = T36[1'h0:1'h0];
  assign T141 = T142 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T142 = T36[1'h0:1'h0];
  assign T143 = T36[1'h1:1'h1];
  assign T144 = T36[2'h2:2'h2];
  assign io_out_valid = T145;
  assign T145 = T158 ? T152 : T146;
  assign T146 = T151 ? T149 : T147;
  assign T147 = T148 ? io_in_1_valid : io_in_0_valid;
  assign T148 = T36[1'h0:1'h0];
  assign T149 = T150 ? io_in_3_valid : io_in_2_valid;
  assign T150 = T36[1'h0:1'h0];
  assign T151 = T36[1'h1:1'h1];
  assign T152 = T157 ? T155 : T153;
  assign T153 = T154 ? io_in_5_valid : io_in_4_valid;
  assign T154 = T36[1'h0:1'h0];
  assign T155 = T156 ? io_in_7_valid : io_in_6_valid;
  assign T156 = T36[1'h0:1'h0];
  assign T157 = T36[1'h1:1'h1];
  assign T158 = T36[2'h2:2'h2];
  assign io_in_0_ready = T159;
  assign T159 = T160 & io_out_ready;
  assign T160 = T185 | T161;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T165 | T163;
  assign T163 = io_in_7_valid & T164;
  assign T164 = R17 < 3'h7;
  assign T165 = T168 | T166;
  assign T166 = io_in_6_valid & T167;
  assign T167 = R17 < 3'h6;
  assign T168 = T171 | T169;
  assign T169 = io_in_5_valid & T170;
  assign T170 = R17 < 3'h5;
  assign T171 = T174 | T172;
  assign T172 = io_in_4_valid & T173;
  assign T173 = R17 < 3'h4;
  assign T174 = T177 | T175;
  assign T175 = io_in_3_valid & T176;
  assign T176 = R17 < 3'h3;
  assign T177 = T180 | T178;
  assign T178 = io_in_2_valid & T179;
  assign T179 = R17 < 3'h2;
  assign T180 = T183 | T181;
  assign T181 = io_in_1_valid & T182;
  assign T182 = R17 < 3'h1;
  assign T183 = io_in_0_valid & T184;
  assign T184 = R17 < 3'h0;
  assign T185 = R17 < 3'h0;
  assign io_in_1_ready = T186;
  assign T186 = T187 & io_out_ready;
  assign T187 = T197 | T188;
  assign T188 = T189 ^ 1'h1;
  assign T189 = T190 | io_in_0_valid;
  assign T190 = T191 | T163;
  assign T191 = T192 | T166;
  assign T192 = T193 | T169;
  assign T193 = T194 | T172;
  assign T194 = T195 | T175;
  assign T195 = T196 | T178;
  assign T196 = T183 | T181;
  assign T197 = T199 & T198;
  assign T198 = R17 < 3'h1;
  assign T199 = T183 ^ 1'h1;
  assign io_in_2_ready = T200;
  assign T200 = T201 & io_out_ready;
  assign T201 = T212 | T202;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T204 | io_in_1_valid;
  assign T204 = T205 | io_in_0_valid;
  assign T205 = T206 | T163;
  assign T206 = T207 | T166;
  assign T207 = T208 | T169;
  assign T208 = T209 | T172;
  assign T209 = T210 | T175;
  assign T210 = T211 | T178;
  assign T211 = T183 | T181;
  assign T212 = T214 & T213;
  assign T213 = R17 < 3'h2;
  assign T214 = T215 ^ 1'h1;
  assign T215 = T183 | T181;
  assign io_in_3_ready = T216;
  assign T216 = T217 & io_out_ready;
  assign T217 = T229 | T218;
  assign T218 = T219 ^ 1'h1;
  assign T219 = T220 | io_in_2_valid;
  assign T220 = T221 | io_in_1_valid;
  assign T221 = T222 | io_in_0_valid;
  assign T222 = T223 | T163;
  assign T223 = T224 | T166;
  assign T224 = T225 | T169;
  assign T225 = T226 | T172;
  assign T226 = T227 | T175;
  assign T227 = T228 | T178;
  assign T228 = T183 | T181;
  assign T229 = T231 & T230;
  assign T230 = R17 < 3'h3;
  assign T231 = T232 ^ 1'h1;
  assign T232 = T233 | T178;
  assign T233 = T183 | T181;
  assign io_in_4_ready = T234;
  assign T234 = T235 & io_out_ready;
  assign T235 = T248 | T236;
  assign T236 = T237 ^ 1'h1;
  assign T237 = T238 | io_in_3_valid;
  assign T238 = T239 | io_in_2_valid;
  assign T239 = T240 | io_in_1_valid;
  assign T240 = T241 | io_in_0_valid;
  assign T241 = T242 | T163;
  assign T242 = T243 | T166;
  assign T243 = T244 | T169;
  assign T244 = T245 | T172;
  assign T245 = T246 | T175;
  assign T246 = T247 | T178;
  assign T247 = T183 | T181;
  assign T248 = T250 & T249;
  assign T249 = R17 < 3'h4;
  assign T250 = T251 ^ 1'h1;
  assign T251 = T252 | T175;
  assign T252 = T253 | T178;
  assign T253 = T183 | T181;
  assign io_in_5_ready = T254;
  assign T254 = T255 & io_out_ready;
  assign T255 = T269 | T256;
  assign T256 = T257 ^ 1'h1;
  assign T257 = T258 | io_in_4_valid;
  assign T258 = T259 | io_in_3_valid;
  assign T259 = T260 | io_in_2_valid;
  assign T260 = T261 | io_in_1_valid;
  assign T261 = T262 | io_in_0_valid;
  assign T262 = T263 | T163;
  assign T263 = T264 | T166;
  assign T264 = T265 | T169;
  assign T265 = T266 | T172;
  assign T266 = T267 | T175;
  assign T267 = T268 | T178;
  assign T268 = T183 | T181;
  assign T269 = T271 & T270;
  assign T270 = R17 < 3'h5;
  assign T271 = T272 ^ 1'h1;
  assign T272 = T273 | T172;
  assign T273 = T274 | T175;
  assign T274 = T275 | T178;
  assign T275 = T183 | T181;
  assign io_in_6_ready = T276;
  assign T276 = T277 & io_out_ready;
  assign T277 = T292 | T278;
  assign T278 = T279 ^ 1'h1;
  assign T279 = T280 | io_in_5_valid;
  assign T280 = T281 | io_in_4_valid;
  assign T281 = T282 | io_in_3_valid;
  assign T282 = T283 | io_in_2_valid;
  assign T283 = T284 | io_in_1_valid;
  assign T284 = T285 | io_in_0_valid;
  assign T285 = T286 | T163;
  assign T286 = T287 | T166;
  assign T287 = T288 | T169;
  assign T288 = T289 | T172;
  assign T289 = T290 | T175;
  assign T290 = T291 | T178;
  assign T291 = T183 | T181;
  assign T292 = T294 & T293;
  assign T293 = R17 < 3'h6;
  assign T294 = T295 ^ 1'h1;
  assign T295 = T296 | T169;
  assign T296 = T297 | T172;
  assign T297 = T298 | T175;
  assign T298 = T299 | T178;
  assign T299 = T183 | T181;
  assign io_in_7_ready = T300;
  assign T300 = T301 & io_out_ready;
  assign T301 = T317 | T302;
  assign T302 = T303 ^ 1'h1;
  assign T303 = T304 | io_in_6_valid;
  assign T304 = T305 | io_in_5_valid;
  assign T305 = T306 | io_in_4_valid;
  assign T306 = T307 | io_in_3_valid;
  assign T307 = T308 | io_in_2_valid;
  assign T308 = T309 | io_in_1_valid;
  assign T309 = T310 | io_in_0_valid;
  assign T310 = T311 | T163;
  assign T311 = T312 | T166;
  assign T312 = T313 | T169;
  assign T313 = T314 | T172;
  assign T314 = T315 | T175;
  assign T315 = T316 | T178;
  assign T316 = T183 | T181;
  assign T317 = T319 & T318;
  assign T318 = R17 < 3'h7;
  assign T319 = T320 ^ 1'h1;
  assign T320 = T321 | T166;
  assign T321 = T322 | T169;
  assign T322 = T323 | T172;
  assign T323 = T324 | T175;
  assign T324 = T325 | T178;
  assign T325 = T183 | T181;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T19) begin
      R17 <= T0;
    end
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input  io_in_7_bits_payload_master_xact_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input  io_in_6_bits_payload_master_xact_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input  io_in_5_bits_payload_master_xact_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input  io_in_4_bits_payload_master_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input  io_in_3_bits_payload_master_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input  io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input  io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input  io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output io_out_bits_payload_master_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T256;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[2:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire T64;
  wire[1:0] T65;
  wire T66;
  wire T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire T70;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T30 ? 3'h1 : T2;
  assign T2 = T28 ? 3'h2 : T3;
  assign T3 = T26 ? 3'h3 : T4;
  assign T4 = T24 ? 3'h4 : T5;
  assign T5 = T22 ? 3'h5 : T6;
  assign T6 = T20 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T256 = reset ? 3'h0 : T18;
  assign T18 = T19 ? T0 : R17;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = io_in_6_valid & T21;
  assign T21 = R17 < 3'h6;
  assign T22 = io_in_5_valid & T23;
  assign T23 = R17 < 3'h5;
  assign T24 = io_in_4_valid & T25;
  assign T25 = R17 < 3'h4;
  assign T26 = io_in_3_valid & T27;
  assign T27 = R17 < 3'h3;
  assign T28 = io_in_2_valid & T29;
  assign T29 = R17 < 3'h2;
  assign T30 = io_in_1_valid & T31;
  assign T31 = R17 < 3'h1;
  assign io_out_bits_payload_master_xact_id = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = T0;
  assign T37 = T38 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T38 = T36[1'h0:1'h0];
  assign T39 = T36[1'h1:1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T42 = T36[1'h0:1'h0];
  assign T43 = T44 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign T46 = T36[2'h2:2'h2];
  assign io_out_bits_header_dst = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T50 = T36[1'h0:1'h0];
  assign T51 = T52 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T58 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T58 = T36[1'h0:1'h0];
  assign T59 = T36[1'h1:1'h1];
  assign T60 = T36[2'h2:2'h2];
  assign io_out_bits_header_src = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T66 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T66 = T36[1'h0:1'h0];
  assign T67 = T36[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T70 = T36[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T72 = T36[1'h0:1'h0];
  assign T73 = T36[1'h1:1'h1];
  assign T74 = T36[2'h2:2'h2];
  assign io_out_valid = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_valid : io_in_0_valid;
  assign T78 = T36[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_valid : io_in_2_valid;
  assign T80 = T36[1'h0:1'h0];
  assign T81 = T36[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_valid : io_in_4_valid;
  assign T84 = T36[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_valid : io_in_6_valid;
  assign T86 = T36[1'h0:1'h0];
  assign T87 = T36[1'h1:1'h1];
  assign T88 = T36[2'h2:2'h2];
  assign io_in_0_ready = T89;
  assign T89 = T90 & io_out_ready;
  assign T90 = T115 | T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T95 | T93;
  assign T93 = io_in_7_valid & T94;
  assign T94 = R17 < 3'h7;
  assign T95 = T98 | T96;
  assign T96 = io_in_6_valid & T97;
  assign T97 = R17 < 3'h6;
  assign T98 = T101 | T99;
  assign T99 = io_in_5_valid & T100;
  assign T100 = R17 < 3'h5;
  assign T101 = T104 | T102;
  assign T102 = io_in_4_valid & T103;
  assign T103 = R17 < 3'h4;
  assign T104 = T107 | T105;
  assign T105 = io_in_3_valid & T106;
  assign T106 = R17 < 3'h3;
  assign T107 = T110 | T108;
  assign T108 = io_in_2_valid & T109;
  assign T109 = R17 < 3'h2;
  assign T110 = T113 | T111;
  assign T111 = io_in_1_valid & T112;
  assign T112 = R17 < 3'h1;
  assign T113 = io_in_0_valid & T114;
  assign T114 = R17 < 3'h0;
  assign T115 = R17 < 3'h0;
  assign io_in_1_ready = T116;
  assign T116 = T117 & io_out_ready;
  assign T117 = T127 | T118;
  assign T118 = T119 ^ 1'h1;
  assign T119 = T120 | io_in_0_valid;
  assign T120 = T121 | T93;
  assign T121 = T122 | T96;
  assign T122 = T123 | T99;
  assign T123 = T124 | T102;
  assign T124 = T125 | T105;
  assign T125 = T126 | T108;
  assign T126 = T113 | T111;
  assign T127 = T129 & T128;
  assign T128 = R17 < 3'h1;
  assign T129 = T113 ^ 1'h1;
  assign io_in_2_ready = T130;
  assign T130 = T131 & io_out_ready;
  assign T131 = T142 | T132;
  assign T132 = T133 ^ 1'h1;
  assign T133 = T134 | io_in_1_valid;
  assign T134 = T135 | io_in_0_valid;
  assign T135 = T136 | T93;
  assign T136 = T137 | T96;
  assign T137 = T138 | T99;
  assign T138 = T139 | T102;
  assign T139 = T140 | T105;
  assign T140 = T141 | T108;
  assign T141 = T113 | T111;
  assign T142 = T144 & T143;
  assign T143 = R17 < 3'h2;
  assign T144 = T145 ^ 1'h1;
  assign T145 = T113 | T111;
  assign io_in_3_ready = T146;
  assign T146 = T147 & io_out_ready;
  assign T147 = T159 | T148;
  assign T148 = T149 ^ 1'h1;
  assign T149 = T150 | io_in_2_valid;
  assign T150 = T151 | io_in_1_valid;
  assign T151 = T152 | io_in_0_valid;
  assign T152 = T153 | T93;
  assign T153 = T154 | T96;
  assign T154 = T155 | T99;
  assign T155 = T156 | T102;
  assign T156 = T157 | T105;
  assign T157 = T158 | T108;
  assign T158 = T113 | T111;
  assign T159 = T161 & T160;
  assign T160 = R17 < 3'h3;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T163 | T108;
  assign T163 = T113 | T111;
  assign io_in_4_ready = T164;
  assign T164 = T165 & io_out_ready;
  assign T165 = T178 | T166;
  assign T166 = T167 ^ 1'h1;
  assign T167 = T168 | io_in_3_valid;
  assign T168 = T169 | io_in_2_valid;
  assign T169 = T170 | io_in_1_valid;
  assign T170 = T171 | io_in_0_valid;
  assign T171 = T172 | T93;
  assign T172 = T173 | T96;
  assign T173 = T174 | T99;
  assign T174 = T175 | T102;
  assign T175 = T176 | T105;
  assign T176 = T177 | T108;
  assign T177 = T113 | T111;
  assign T178 = T180 & T179;
  assign T179 = R17 < 3'h4;
  assign T180 = T181 ^ 1'h1;
  assign T181 = T182 | T105;
  assign T182 = T183 | T108;
  assign T183 = T113 | T111;
  assign io_in_5_ready = T184;
  assign T184 = T185 & io_out_ready;
  assign T185 = T199 | T186;
  assign T186 = T187 ^ 1'h1;
  assign T187 = T188 | io_in_4_valid;
  assign T188 = T189 | io_in_3_valid;
  assign T189 = T190 | io_in_2_valid;
  assign T190 = T191 | io_in_1_valid;
  assign T191 = T192 | io_in_0_valid;
  assign T192 = T193 | T93;
  assign T193 = T194 | T96;
  assign T194 = T195 | T99;
  assign T195 = T196 | T102;
  assign T196 = T197 | T105;
  assign T197 = T198 | T108;
  assign T198 = T113 | T111;
  assign T199 = T201 & T200;
  assign T200 = R17 < 3'h5;
  assign T201 = T202 ^ 1'h1;
  assign T202 = T203 | T102;
  assign T203 = T204 | T105;
  assign T204 = T205 | T108;
  assign T205 = T113 | T111;
  assign io_in_6_ready = T206;
  assign T206 = T207 & io_out_ready;
  assign T207 = T222 | T208;
  assign T208 = T209 ^ 1'h1;
  assign T209 = T210 | io_in_5_valid;
  assign T210 = T211 | io_in_4_valid;
  assign T211 = T212 | io_in_3_valid;
  assign T212 = T213 | io_in_2_valid;
  assign T213 = T214 | io_in_1_valid;
  assign T214 = T215 | io_in_0_valid;
  assign T215 = T216 | T93;
  assign T216 = T217 | T96;
  assign T217 = T218 | T99;
  assign T218 = T219 | T102;
  assign T219 = T220 | T105;
  assign T220 = T221 | T108;
  assign T221 = T113 | T111;
  assign T222 = T224 & T223;
  assign T223 = R17 < 3'h6;
  assign T224 = T225 ^ 1'h1;
  assign T225 = T226 | T99;
  assign T226 = T227 | T102;
  assign T227 = T228 | T105;
  assign T228 = T229 | T108;
  assign T229 = T113 | T111;
  assign io_in_7_ready = T230;
  assign T230 = T231 & io_out_ready;
  assign T231 = T247 | T232;
  assign T232 = T233 ^ 1'h1;
  assign T233 = T234 | io_in_6_valid;
  assign T234 = T235 | io_in_5_valid;
  assign T235 = T236 | io_in_4_valid;
  assign T236 = T237 | io_in_3_valid;
  assign T237 = T238 | io_in_2_valid;
  assign T238 = T239 | io_in_1_valid;
  assign T239 = T240 | io_in_0_valid;
  assign T240 = T241 | T93;
  assign T241 = T242 | T96;
  assign T242 = T243 | T99;
  assign T243 = T244 | T102;
  assign T244 = T245 | T105;
  assign T245 = T246 | T108;
  assign T246 = T113 | T111;
  assign T247 = T249 & T248;
  assign T248 = R17 < 3'h7;
  assign T249 = T250 ^ 1'h1;
  assign T250 = T251 | T96;
  assign T251 = T252 | T99;
  assign T252 = T253 | T102;
  assign T253 = T254 | T105;
  assign T254 = T255 | T108;
  assign T255 = T113 | T111;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T19) begin
      R17 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatPassesId(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [1:0] io_in_7_acquire_bits_header_src,
    input [1:0] io_in_7_acquire_bits_header_dst,
    input [25:0] io_in_7_acquire_bits_payload_addr,
    input [2:0] io_in_7_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_7_acquire_bits_payload_data,
    input  io_in_7_acquire_bits_payload_uncached,
    input [1:0] io_in_7_acquire_bits_payload_a_type,
    input [7:0] io_in_7_acquire_bits_payload_subblock,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_header_src,
    output[1:0] io_in_7_grant_bits_header_dst,
    output[2:0] io_in_7_grant_bits_payload_data,
    output[2:0] io_in_7_grant_bits_payload_client_xact_id,
    output io_in_7_grant_bits_payload_master_xact_id,
    output io_in_7_grant_bits_payload_uncached,
    output[1:0] io_in_7_grant_bits_payload_g_type,
    output io_in_7_finish_ready,
    input  io_in_7_finish_valid,
    input [1:0] io_in_7_finish_bits_header_src,
    input [1:0] io_in_7_finish_bits_header_dst,
    input  io_in_7_finish_bits_payload_master_xact_id,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [1:0] io_in_6_acquire_bits_header_src,
    input [1:0] io_in_6_acquire_bits_header_dst,
    input [25:0] io_in_6_acquire_bits_payload_addr,
    input [2:0] io_in_6_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_6_acquire_bits_payload_data,
    input  io_in_6_acquire_bits_payload_uncached,
    input [1:0] io_in_6_acquire_bits_payload_a_type,
    input [7:0] io_in_6_acquire_bits_payload_subblock,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_header_src,
    output[1:0] io_in_6_grant_bits_header_dst,
    output[2:0] io_in_6_grant_bits_payload_data,
    output[2:0] io_in_6_grant_bits_payload_client_xact_id,
    output io_in_6_grant_bits_payload_master_xact_id,
    output io_in_6_grant_bits_payload_uncached,
    output[1:0] io_in_6_grant_bits_payload_g_type,
    output io_in_6_finish_ready,
    input  io_in_6_finish_valid,
    input [1:0] io_in_6_finish_bits_header_src,
    input [1:0] io_in_6_finish_bits_header_dst,
    input  io_in_6_finish_bits_payload_master_xact_id,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [1:0] io_in_5_acquire_bits_header_src,
    input [1:0] io_in_5_acquire_bits_header_dst,
    input [25:0] io_in_5_acquire_bits_payload_addr,
    input [2:0] io_in_5_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_5_acquire_bits_payload_data,
    input  io_in_5_acquire_bits_payload_uncached,
    input [1:0] io_in_5_acquire_bits_payload_a_type,
    input [7:0] io_in_5_acquire_bits_payload_subblock,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_header_src,
    output[1:0] io_in_5_grant_bits_header_dst,
    output[2:0] io_in_5_grant_bits_payload_data,
    output[2:0] io_in_5_grant_bits_payload_client_xact_id,
    output io_in_5_grant_bits_payload_master_xact_id,
    output io_in_5_grant_bits_payload_uncached,
    output[1:0] io_in_5_grant_bits_payload_g_type,
    output io_in_5_finish_ready,
    input  io_in_5_finish_valid,
    input [1:0] io_in_5_finish_bits_header_src,
    input [1:0] io_in_5_finish_bits_header_dst,
    input  io_in_5_finish_bits_payload_master_xact_id,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [1:0] io_in_4_acquire_bits_header_src,
    input [1:0] io_in_4_acquire_bits_header_dst,
    input [25:0] io_in_4_acquire_bits_payload_addr,
    input [2:0] io_in_4_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_4_acquire_bits_payload_data,
    input  io_in_4_acquire_bits_payload_uncached,
    input [1:0] io_in_4_acquire_bits_payload_a_type,
    input [7:0] io_in_4_acquire_bits_payload_subblock,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_header_src,
    output[1:0] io_in_4_grant_bits_header_dst,
    output[2:0] io_in_4_grant_bits_payload_data,
    output[2:0] io_in_4_grant_bits_payload_client_xact_id,
    output io_in_4_grant_bits_payload_master_xact_id,
    output io_in_4_grant_bits_payload_uncached,
    output[1:0] io_in_4_grant_bits_payload_g_type,
    output io_in_4_finish_ready,
    input  io_in_4_finish_valid,
    input [1:0] io_in_4_finish_bits_header_src,
    input [1:0] io_in_4_finish_bits_header_dst,
    input  io_in_4_finish_bits_payload_master_xact_id,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [1:0] io_in_3_acquire_bits_header_src,
    input [1:0] io_in_3_acquire_bits_header_dst,
    input [25:0] io_in_3_acquire_bits_payload_addr,
    input [2:0] io_in_3_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_3_acquire_bits_payload_data,
    input  io_in_3_acquire_bits_payload_uncached,
    input [1:0] io_in_3_acquire_bits_payload_a_type,
    input [7:0] io_in_3_acquire_bits_payload_subblock,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_header_src,
    output[1:0] io_in_3_grant_bits_header_dst,
    output[2:0] io_in_3_grant_bits_payload_data,
    output[2:0] io_in_3_grant_bits_payload_client_xact_id,
    output io_in_3_grant_bits_payload_master_xact_id,
    output io_in_3_grant_bits_payload_uncached,
    output[1:0] io_in_3_grant_bits_payload_g_type,
    output io_in_3_finish_ready,
    input  io_in_3_finish_valid,
    input [1:0] io_in_3_finish_bits_header_src,
    input [1:0] io_in_3_finish_bits_header_dst,
    input  io_in_3_finish_bits_payload_master_xact_id,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [2:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_2_acquire_bits_payload_data,
    input  io_in_2_acquire_bits_payload_uncached,
    input [1:0] io_in_2_acquire_bits_payload_a_type,
    input [7:0] io_in_2_acquire_bits_payload_subblock,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[2:0] io_in_2_grant_bits_payload_data,
    output[2:0] io_in_2_grant_bits_payload_client_xact_id,
    output io_in_2_grant_bits_payload_master_xact_id,
    output io_in_2_grant_bits_payload_uncached,
    output[1:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input  io_in_2_finish_bits_payload_master_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [2:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_1_acquire_bits_payload_data,
    input  io_in_1_acquire_bits_payload_uncached,
    input [1:0] io_in_1_acquire_bits_payload_a_type,
    input [7:0] io_in_1_acquire_bits_payload_subblock,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[2:0] io_in_1_grant_bits_payload_data,
    output[2:0] io_in_1_grant_bits_payload_client_xact_id,
    output io_in_1_grant_bits_payload_master_xact_id,
    output io_in_1_grant_bits_payload_uncached,
    output[1:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input  io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [2:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [2:0] io_in_0_acquire_bits_payload_data,
    input  io_in_0_acquire_bits_payload_uncached,
    input [1:0] io_in_0_acquire_bits_payload_a_type,
    input [7:0] io_in_0_acquire_bits_payload_subblock,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[2:0] io_in_0_grant_bits_payload_data,
    output[2:0] io_in_0_grant_bits_payload_client_xact_id,
    output io_in_0_grant_bits_payload_master_xact_id,
    output io_in_0_grant_bits_payload_uncached,
    output[1:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input  io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[2:0] io_out_acquire_bits_payload_client_xact_id,
    output[2:0] io_out_acquire_bits_payload_data,
    output io_out_acquire_bits_payload_uncached,
    output[1:0] io_out_acquire_bits_payload_a_type,
    output[7:0] io_out_acquire_bits_payload_subblock,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [2:0] io_out_grant_bits_payload_data,
    input [2:0] io_out_grant_bits_payload_client_xact_id,
    input  io_out_grant_bits_payload_master_xact_id,
    input  io_out_grant_bits_payload_uncached,
    input [1:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output io_out_finish_bits_payload_master_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire RRArbiter_2_io_in_7_ready;
  wire RRArbiter_2_io_in_6_ready;
  wire RRArbiter_2_io_in_5_ready;
  wire RRArbiter_2_io_in_4_ready;
  wire RRArbiter_2_io_in_3_ready;
  wire RRArbiter_2_io_in_2_ready;
  wire RRArbiter_2_io_in_1_ready;
  wire RRArbiter_2_io_in_0_ready;
  wire RRArbiter_2_io_out_valid;
  wire[1:0] RRArbiter_2_io_out_bits_header_src;
  wire[1:0] RRArbiter_2_io_out_bits_header_dst;
  wire[25:0] RRArbiter_2_io_out_bits_payload_addr;
  wire[2:0] RRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[2:0] RRArbiter_2_io_out_bits_payload_data;
  wire RRArbiter_2_io_out_bits_payload_uncached;
  wire[1:0] RRArbiter_2_io_out_bits_payload_a_type;
  wire[7:0] RRArbiter_2_io_out_bits_payload_subblock;
  wire RRArbiter_3_io_in_7_ready;
  wire RRArbiter_3_io_in_6_ready;
  wire RRArbiter_3_io_in_5_ready;
  wire RRArbiter_3_io_in_4_ready;
  wire RRArbiter_3_io_in_3_ready;
  wire RRArbiter_3_io_in_2_ready;
  wire RRArbiter_3_io_in_1_ready;
  wire RRArbiter_3_io_in_0_ready;
  wire RRArbiter_3_io_out_valid;
  wire[1:0] RRArbiter_3_io_out_bits_header_src;
  wire[1:0] RRArbiter_3_io_out_bits_header_dst;
  wire RRArbiter_3_io_out_bits_payload_master_xact_id;


  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_3_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_3_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_3_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_3_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T15 ? io_in_7_grant_ready : T1;
  assign T1 = T14 ? io_in_6_grant_ready : T2;
  assign T2 = T13 ? io_in_5_grant_ready : T3;
  assign T3 = T12 ? io_in_4_grant_ready : T4;
  assign T4 = T11 ? io_in_3_grant_ready : T5;
  assign T5 = T10 ? io_in_2_grant_ready : T6;
  assign T6 = T9 ? io_in_1_grant_ready : T7;
  assign T7 = T8 ? io_in_0_grant_ready : 1'h0;
  assign T8 = io_out_grant_bits_payload_client_xact_id == 3'h0;
  assign T9 = io_out_grant_bits_payload_client_xact_id == 3'h1;
  assign T10 = io_out_grant_bits_payload_client_xact_id == 3'h2;
  assign T11 = io_out_grant_bits_payload_client_xact_id == 3'h3;
  assign T12 = io_out_grant_bits_payload_client_xact_id == 3'h4;
  assign T13 = io_out_grant_bits_payload_client_xact_id == 3'h5;
  assign T14 = io_out_grant_bits_payload_client_xact_id == 3'h6;
  assign T15 = io_out_grant_bits_payload_client_xact_id == 3'h7;
  assign io_out_acquire_bits_payload_subblock = RRArbiter_2_io_out_bits_payload_subblock;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_uncached = RRArbiter_2_io_out_bits_payload_uncached;
  assign io_out_acquire_bits_payload_data = RRArbiter_2_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_2_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_2_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_2_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_2_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_3_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T16;
  assign T16 = T8 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_2_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_3_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_2_io_in_1_ready;
  assign io_in_2_finish_ready = RRArbiter_3_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_2_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T18;
  assign T18 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = RRArbiter_2_io_in_2_ready;
  assign io_in_3_finish_ready = RRArbiter_3_io_in_3_ready;
  assign io_in_3_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_3_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_3_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_3_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_3_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_3_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_3_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_3_grant_valid = T19;
  assign T19 = T11 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = RRArbiter_2_io_in_3_ready;
  assign io_in_4_finish_ready = RRArbiter_3_io_in_4_ready;
  assign io_in_4_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_4_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_4_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_4_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_4_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_4_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_4_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_4_grant_valid = T20;
  assign T20 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = RRArbiter_2_io_in_4_ready;
  assign io_in_5_finish_ready = RRArbiter_3_io_in_5_ready;
  assign io_in_5_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_5_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_5_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_5_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_5_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_5_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_5_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_5_grant_valid = T21;
  assign T21 = T13 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = RRArbiter_2_io_in_5_ready;
  assign io_in_6_finish_ready = RRArbiter_3_io_in_6_ready;
  assign io_in_6_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_6_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_6_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_6_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_6_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_6_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_6_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_6_grant_valid = T22;
  assign T22 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = RRArbiter_2_io_in_6_ready;
  assign io_in_7_finish_ready = RRArbiter_3_io_in_7_ready;
  assign io_in_7_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_7_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_7_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_7_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_7_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_7_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_7_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_7_grant_valid = T23;
  assign T23 = T15 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = RRArbiter_2_io_in_7_ready;
  RRArbiter_3 RRArbiter_2(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_2_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_header_src( io_in_7_acquire_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_acquire_bits_header_dst ),
       .io_in_7_bits_payload_addr( io_in_7_acquire_bits_payload_addr ),
       .io_in_7_bits_payload_client_xact_id( io_in_7_acquire_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_data( io_in_7_acquire_bits_payload_data ),
       .io_in_7_bits_payload_uncached( io_in_7_acquire_bits_payload_uncached ),
       .io_in_7_bits_payload_a_type( io_in_7_acquire_bits_payload_a_type ),
       .io_in_7_bits_payload_subblock( io_in_7_acquire_bits_payload_subblock ),
       .io_in_6_ready( RRArbiter_2_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_header_src( io_in_6_acquire_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_acquire_bits_header_dst ),
       .io_in_6_bits_payload_addr( io_in_6_acquire_bits_payload_addr ),
       .io_in_6_bits_payload_client_xact_id( io_in_6_acquire_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_data( io_in_6_acquire_bits_payload_data ),
       .io_in_6_bits_payload_uncached( io_in_6_acquire_bits_payload_uncached ),
       .io_in_6_bits_payload_a_type( io_in_6_acquire_bits_payload_a_type ),
       .io_in_6_bits_payload_subblock( io_in_6_acquire_bits_payload_subblock ),
       .io_in_5_ready( RRArbiter_2_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_header_src( io_in_5_acquire_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_acquire_bits_header_dst ),
       .io_in_5_bits_payload_addr( io_in_5_acquire_bits_payload_addr ),
       .io_in_5_bits_payload_client_xact_id( io_in_5_acquire_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_data( io_in_5_acquire_bits_payload_data ),
       .io_in_5_bits_payload_uncached( io_in_5_acquire_bits_payload_uncached ),
       .io_in_5_bits_payload_a_type( io_in_5_acquire_bits_payload_a_type ),
       .io_in_5_bits_payload_subblock( io_in_5_acquire_bits_payload_subblock ),
       .io_in_4_ready( RRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_header_src( io_in_4_acquire_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_acquire_bits_header_dst ),
       .io_in_4_bits_payload_addr( io_in_4_acquire_bits_payload_addr ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_acquire_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_data( io_in_4_acquire_bits_payload_data ),
       .io_in_4_bits_payload_uncached( io_in_4_acquire_bits_payload_uncached ),
       .io_in_4_bits_payload_a_type( io_in_4_acquire_bits_payload_a_type ),
       .io_in_4_bits_payload_subblock( io_in_4_acquire_bits_payload_subblock ),
       .io_in_3_ready( RRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_header_src( io_in_3_acquire_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_acquire_bits_header_dst ),
       .io_in_3_bits_payload_addr( io_in_3_acquire_bits_payload_addr ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_acquire_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_data( io_in_3_acquire_bits_payload_data ),
       .io_in_3_bits_payload_uncached( io_in_3_acquire_bits_payload_uncached ),
       .io_in_3_bits_payload_a_type( io_in_3_acquire_bits_payload_a_type ),
       .io_in_3_bits_payload_subblock( io_in_3_acquire_bits_payload_subblock ),
       .io_in_2_ready( RRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_acquire_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_acquire_bits_payload_subblock ),
       .io_in_1_ready( RRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_acquire_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_acquire_bits_payload_subblock ),
       .io_in_0_ready( RRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_acquire_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_acquire_bits_payload_subblock ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( RRArbiter_2_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( RRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( RRArbiter_2_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  RRArbiter_4 RRArbiter_3(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_3_io_in_7_ready ),
       .io_in_7_valid( io_in_7_finish_valid ),
       .io_in_7_bits_header_src( io_in_7_finish_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_finish_bits_header_dst ),
       .io_in_7_bits_payload_master_xact_id( io_in_7_finish_bits_payload_master_xact_id ),
       .io_in_6_ready( RRArbiter_3_io_in_6_ready ),
       .io_in_6_valid( io_in_6_finish_valid ),
       .io_in_6_bits_header_src( io_in_6_finish_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_finish_bits_header_dst ),
       .io_in_6_bits_payload_master_xact_id( io_in_6_finish_bits_payload_master_xact_id ),
       .io_in_5_ready( RRArbiter_3_io_in_5_ready ),
       .io_in_5_valid( io_in_5_finish_valid ),
       .io_in_5_bits_header_src( io_in_5_finish_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_finish_bits_header_dst ),
       .io_in_5_bits_payload_master_xact_id( io_in_5_finish_bits_payload_master_xact_id ),
       .io_in_4_ready( RRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( io_in_4_finish_valid ),
       .io_in_4_bits_header_src( io_in_4_finish_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_finish_bits_header_dst ),
       .io_in_4_bits_payload_master_xact_id( io_in_4_finish_bits_payload_master_xact_id ),
       .io_in_3_ready( RRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( io_in_3_finish_valid ),
       .io_in_3_bits_header_src( io_in_3_finish_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_finish_bits_header_dst ),
       .io_in_3_bits_payload_master_xact_id( io_in_3_finish_bits_payload_master_xact_id ),
       .io_in_2_ready( RRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_finish_bits_payload_master_xact_id ),
       .io_in_1_ready( RRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_3_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module L2CoherenceAgent(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [2:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [511:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[2:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [2:0] io_inner_release_bits_payload_client_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    output[1:0] io_outer_acquire_bits_header_dst,
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[511:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    output io_outer_finish_valid,
    output[1:0] io_outer_finish_bits_header_src,
    output[1:0] io_outer_finish_bits_header_dst,
    output io_outer_finish_bits_payload_master_xact_id,
    input  io_incoherent_1,
    input  io_incoherent_0
);

  wire[2:0] T85;
  wire[511:0] T86;
  wire[511:0] T87;
  wire[511:0] T88;
  wire[511:0] T89;
  wire[511:0] T90;
  wire[511:0] T91;
  wire[511:0] T92;
  wire[511:0] T93;
  wire T94;
  wire T95;
  wire any_acquire_conflict;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T96;
  wire sdq_rdy;
  wire T67;
  reg  sdq_val;
  wire T79;
  wire[3:0] T80;
  wire[3:0] T21;
  wire[3:0] T81;
  wire[3:0] T22;
  wire[3:0] T82;
  wire T23;
  wire sdq_enq;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[3:0] T83;
  wire free_sdq;
  wire is_in_sdq;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire[1:0] free_sdq_id;
  wire[3:0] T84;
  wire T37;
  wire[1:0] T97;
  wire[1:0] T98;
  wire T99;
  wire T100;
  wire[2:0] release_idx;
  wire[2:0] conflict_idx;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T77;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T78;
  wire voluntary;
  wire[7:0] T101;
  wire[2:0] T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire[7:0] T107;
  wire[2:0] T108;
  wire[1:0] T109;
  wire[1:0] T110;
  wire T111;
  wire T112;
  wire[7:0] T113;
  wire[2:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire[7:0] T119;
  wire[2:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire T124;
  wire[7:0] T125;
  wire[2:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire T129;
  wire T130;
  wire[7:0] T131;
  wire[2:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire[7:0] T137;
  wire[2:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire[7:0] T143;
  wire[2:0] T144;
  wire[1:0] T145;
  wire[511:0] T75;
  wire[511:0] T0;
  wire[511:0] T1;
  reg [511:0] vwbdq_0;
  wire[511:0] T2;
  wire T3;
  wire T4;
  wire[1:0] T5;
  wire T6;
  wire T76;
  wire T12;
  wire T13;
  wire is_in_vwbdq;
  reg [511:0] sdq_0;
  wire[511:0] T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[2:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T66;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire VoluntaryReleaseTracker_io_inner_acquire_ready;
  wire VoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_src;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_dst;
  wire[2:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_data;
  wire[2:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id;
  wire VoluntaryReleaseTracker_io_inner_grant_bits_payload_uncached;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type;
  wire VoluntaryReleaseTracker_io_inner_probe_valid;
  wire VoluntaryReleaseTracker_io_inner_release_ready;
  wire VoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_header_src;
  wire[25:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data;
  wire VoluntaryReleaseTracker_io_outer_acquire_bits_payload_uncached;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type;
  wire[7:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subblock;
  wire VoluntaryReleaseTracker_io_outer_grant_ready;
  wire VoluntaryReleaseTracker_io_has_acquire_conflict;
  wire AcquireTracker_0_io_inner_acquire_ready;
  wire AcquireTracker_0_io_inner_grant_valid;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_0_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_0_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_0_io_inner_probe_valid;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_0_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_0_io_inner_release_ready;
  wire AcquireTracker_0_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_0_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_0_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_0_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_0_io_outer_grant_ready;
  wire AcquireTracker_0_io_has_acquire_conflict;
  wire AcquireTracker_0_io_has_release_conflict;
  wire AcquireTracker_1_io_inner_acquire_ready;
  wire AcquireTracker_1_io_inner_grant_valid;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_1_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_1_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_1_io_inner_probe_valid;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_1_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_1_io_inner_release_ready;
  wire AcquireTracker_1_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_1_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_1_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_1_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_1_io_outer_grant_ready;
  wire AcquireTracker_1_io_has_acquire_conflict;
  wire AcquireTracker_1_io_has_release_conflict;
  wire AcquireTracker_2_io_inner_acquire_ready;
  wire AcquireTracker_2_io_inner_grant_valid;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_2_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_2_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_2_io_inner_probe_valid;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_2_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_2_io_inner_release_ready;
  wire AcquireTracker_2_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_2_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_2_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_2_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_2_io_outer_grant_ready;
  wire AcquireTracker_2_io_has_acquire_conflict;
  wire AcquireTracker_2_io_has_release_conflict;
  wire AcquireTracker_3_io_inner_acquire_ready;
  wire AcquireTracker_3_io_inner_grant_valid;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_3_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_3_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_3_io_inner_probe_valid;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_3_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_3_io_inner_release_ready;
  wire AcquireTracker_3_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_3_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_3_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_3_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_3_io_outer_grant_ready;
  wire AcquireTracker_3_io_has_acquire_conflict;
  wire AcquireTracker_3_io_has_release_conflict;
  wire AcquireTracker_4_io_inner_acquire_ready;
  wire AcquireTracker_4_io_inner_grant_valid;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_4_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_4_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_4_io_inner_probe_valid;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_4_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_4_io_inner_release_ready;
  wire AcquireTracker_4_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_4_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_4_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_4_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_4_io_outer_grant_ready;
  wire AcquireTracker_4_io_has_acquire_conflict;
  wire AcquireTracker_4_io_has_release_conflict;
  wire AcquireTracker_5_io_inner_acquire_ready;
  wire AcquireTracker_5_io_inner_grant_valid;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_5_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_5_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_5_io_inner_probe_valid;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_5_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_5_io_inner_release_ready;
  wire AcquireTracker_5_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_5_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_5_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_5_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_5_io_outer_grant_ready;
  wire AcquireTracker_5_io_has_acquire_conflict;
  wire AcquireTracker_5_io_has_release_conflict;
  wire AcquireTracker_6_io_inner_acquire_ready;
  wire AcquireTracker_6_io_inner_grant_valid;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_dst;
  wire[2:0] AcquireTracker_6_io_inner_grant_bits_payload_data;
  wire[2:0] AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id;
  wire AcquireTracker_6_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_6_io_inner_probe_valid;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_6_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_6_io_inner_release_ready;
  wire AcquireTracker_6_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_6_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_6_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_payload_a_type;
  wire[7:0] AcquireTracker_6_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_6_io_outer_grant_ready;
  wire AcquireTracker_6_io_has_acquire_conflict;
  wire AcquireTracker_6_io_has_release_conflict;
  wire alloc_arb_io_in_7_ready;
  wire alloc_arb_io_in_6_ready;
  wire alloc_arb_io_in_5_ready;
  wire alloc_arb_io_in_4_ready;
  wire alloc_arb_io_in_3_ready;
  wire alloc_arb_io_in_2_ready;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire probe_arb_io_in_7_ready;
  wire probe_arb_io_in_6_ready;
  wire probe_arb_io_in_5_ready;
  wire probe_arb_io_in_4_ready;
  wire probe_arb_io_in_3_ready;
  wire probe_arb_io_in_2_ready;
  wire probe_arb_io_in_1_ready;
  wire probe_arb_io_in_0_ready;
  wire probe_arb_io_out_valid;
  wire[1:0] probe_arb_io_out_bits_header_src;
  wire[1:0] probe_arb_io_out_bits_header_dst;
  wire[25:0] probe_arb_io_out_bits_payload_addr;
  wire[1:0] probe_arb_io_out_bits_payload_p_type;
  wire grant_arb_io_in_7_ready;
  wire grant_arb_io_in_6_ready;
  wire grant_arb_io_in_5_ready;
  wire grant_arb_io_in_4_ready;
  wire grant_arb_io_in_3_ready;
  wire grant_arb_io_in_2_ready;
  wire grant_arb_io_in_1_ready;
  wire grant_arb_io_in_0_ready;
  wire grant_arb_io_out_valid;
  wire[1:0] grant_arb_io_out_bits_header_src;
  wire[1:0] grant_arb_io_out_bits_header_dst;
  wire[2:0] grant_arb_io_out_bits_payload_client_xact_id;
  wire[2:0] grant_arb_io_out_bits_payload_master_xact_id;
  wire grant_arb_io_out_bits_payload_uncached;
  wire[1:0] grant_arb_io_out_bits_payload_g_type;
  wire outer_arb_io_in_7_acquire_ready;
  wire outer_arb_io_in_7_grant_valid;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_7_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_7_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_7_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_7_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_7_grant_bits_payload_g_type;
  wire outer_arb_io_in_7_finish_ready;
  wire outer_arb_io_in_6_acquire_ready;
  wire outer_arb_io_in_6_grant_valid;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_6_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_6_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_6_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_6_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_6_grant_bits_payload_g_type;
  wire outer_arb_io_in_6_finish_ready;
  wire outer_arb_io_in_5_acquire_ready;
  wire outer_arb_io_in_5_grant_valid;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_5_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_5_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_5_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_5_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_5_grant_bits_payload_g_type;
  wire outer_arb_io_in_5_finish_ready;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_4_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_4_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_4_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_4_grant_bits_payload_g_type;
  wire outer_arb_io_in_4_finish_ready;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_3_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_3_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_3_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_3_grant_bits_payload_g_type;
  wire outer_arb_io_in_3_finish_ready;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_2_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_2_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_2_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_2_grant_bits_payload_g_type;
  wire outer_arb_io_in_2_finish_ready;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_1_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_1_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_1_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_1_grant_bits_payload_g_type;
  wire outer_arb_io_in_1_finish_ready;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_dst;
  wire[2:0] outer_arb_io_in_0_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_0_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_payload_master_xact_id;
  wire outer_arb_io_in_0_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_0_grant_bits_payload_g_type;
  wire outer_arb_io_in_0_finish_ready;
  wire outer_arb_io_out_acquire_valid;
  wire[1:0] outer_arb_io_out_acquire_bits_header_src;
  wire[1:0] outer_arb_io_out_acquire_bits_header_dst;
  wire[25:0] outer_arb_io_out_acquire_bits_payload_addr;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_data;
  wire outer_arb_io_out_acquire_bits_payload_uncached;
  wire[1:0] outer_arb_io_out_acquire_bits_payload_a_type;
  wire[7:0] outer_arb_io_out_acquire_bits_payload_subblock;
  wire outer_arb_io_out_grant_ready;
  wire outer_arb_io_out_finish_valid;
  wire[1:0] outer_arb_io_out_finish_bits_header_src;
  wire[1:0] outer_arb_io_out_finish_bits_header_dst;
  wire outer_arb_io_out_finish_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    vwbdq_0 = {16{$random}};
    sdq_0 = {16{$random}};
  end
`endif

  assign T85 = io_outer_grant_bits_payload_data[2'h2:1'h0];
  assign T86 = {509'h0, VoluntaryReleaseTracker_io_inner_grant_bits_payload_data};
  assign T87 = {509'h0, AcquireTracker_0_io_inner_grant_bits_payload_data};
  assign T88 = {509'h0, AcquireTracker_1_io_inner_grant_bits_payload_data};
  assign T89 = {509'h0, AcquireTracker_2_io_inner_grant_bits_payload_data};
  assign T90 = {509'h0, AcquireTracker_3_io_inner_grant_bits_payload_data};
  assign T91 = {509'h0, AcquireTracker_4_io_inner_grant_bits_payload_data};
  assign T92 = {509'h0, AcquireTracker_5_io_inner_grant_bits_payload_data};
  assign T93 = {509'h0, AcquireTracker_6_io_inner_grant_bits_payload_data};
  assign T94 = T96 & T95;
  assign T95 = any_acquire_conflict ^ 1'h1;
  assign any_acquire_conflict = T60 | AcquireTracker_6_io_has_acquire_conflict;
  assign T60 = T61 | AcquireTracker_5_io_has_acquire_conflict;
  assign T61 = T62 | AcquireTracker_4_io_has_acquire_conflict;
  assign T62 = T63 | AcquireTracker_3_io_has_acquire_conflict;
  assign T63 = T64 | AcquireTracker_2_io_has_acquire_conflict;
  assign T64 = T65 | AcquireTracker_1_io_has_acquire_conflict;
  assign T65 = VoluntaryReleaseTracker_io_has_acquire_conflict | AcquireTracker_0_io_has_acquire_conflict;
  assign T96 = io_inner_acquire_valid & sdq_rdy;
  assign sdq_rdy = T67 ^ 1'h1;
  assign T67 = sdq_val == 1'h1;
  assign T79 = T80[1'h0:1'h0];
  assign T80 = reset ? 4'h0 : T21;
  assign T21 = T37 ? T22 : T81;
  assign T81 = {3'h0, sdq_val};
  assign T22 = T27 | T82;
  assign T82 = {3'h0, T23};
  assign T23 = T24 & sdq_enq;
  assign sdq_enq = T42 & T38;
  assign T38 = io_inner_acquire_bits_payload_uncached ? T39 : 1'h0;
  assign T39 = T41 | T40;
  assign T40 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T41 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T42 = io_inner_acquire_valid & io_inner_acquire_ready;
  assign T24 = T25;
  assign T25 = ~ T26;
  assign T26 = sdq_val;
  assign T27 = T84 & T28;
  assign T28 = ~ T29;
  assign T29 = T36 & T83;
  assign T83 = {3'h0, free_sdq};
  assign free_sdq = T30 & is_in_sdq;
  assign is_in_sdq = outer_arb_io_out_acquire_bits_payload_data[1'h0:1'h0];
  assign T30 = T35 & T31;
  assign T31 = io_outer_acquire_bits_payload_uncached ? T32 : 1'h0;
  assign T32 = T34 | T33;
  assign T33 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T34 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T35 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T36 = 1'h1 << free_sdq_id;
  assign free_sdq_id = outer_arb_io_out_acquire_bits_payload_data >> 1'h1;
  assign T84 = {3'h0, sdq_val};
  assign T37 = io_outer_acquire_valid | sdq_enq;
  assign T97 = T98;
  assign T98 = {io_incoherent_1, io_incoherent_0};
  assign T99 = io_inner_release_valid & T100;
  assign T100 = release_idx == 3'h7;
  assign release_idx = voluntary ? 3'h0 : conflict_idx;
  assign conflict_idx = AcquireTracker_6_io_has_release_conflict ? 3'h7 : T7;
  assign T7 = AcquireTracker_5_io_has_release_conflict ? 3'h6 : T8;
  assign T8 = AcquireTracker_4_io_has_release_conflict ? 3'h5 : T9;
  assign T9 = AcquireTracker_3_io_has_release_conflict ? 3'h4 : T77;
  assign T77 = {1'h0, T10};
  assign T10 = AcquireTracker_2_io_has_release_conflict ? 2'h3 : T11;
  assign T11 = AcquireTracker_1_io_has_release_conflict ? 2'h2 : T78;
  assign T78 = {1'h0, AcquireTracker_0_io_has_release_conflict};
  assign voluntary = io_inner_release_bits_payload_r_type == 3'h0;
  assign T101 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T102 = {1'h0, T103};
  assign T103 = {1'h0, 1'h1};
  assign T104 = T98;
  assign T105 = io_inner_release_valid & T106;
  assign T106 = release_idx == 3'h6;
  assign T107 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T108 = {1'h0, T109};
  assign T109 = {1'h0, 1'h1};
  assign T110 = T98;
  assign T111 = io_inner_release_valid & T112;
  assign T112 = release_idx == 3'h5;
  assign T113 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T114 = {1'h0, T115};
  assign T115 = {1'h0, 1'h1};
  assign T116 = T98;
  assign T117 = io_inner_release_valid & T118;
  assign T118 = release_idx == 3'h4;
  assign T119 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T120 = {1'h0, T121};
  assign T121 = {1'h0, 1'h1};
  assign T122 = T98;
  assign T123 = io_inner_release_valid & T124;
  assign T124 = release_idx == 3'h3;
  assign T125 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T126 = {1'h0, T127};
  assign T127 = {1'h0, 1'h1};
  assign T128 = T98;
  assign T129 = io_inner_release_valid & T130;
  assign T130 = release_idx == 3'h2;
  assign T131 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T132 = {1'h0, T133};
  assign T133 = {1'h0, 1'h1};
  assign T134 = T98;
  assign T135 = io_inner_release_valid & T136;
  assign T136 = release_idx == 3'h1;
  assign T137 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T138 = {1'h0, T139};
  assign T139 = {1'h0, 1'h1};
  assign T140 = T98;
  assign T141 = io_inner_release_valid & T142;
  assign T142 = release_idx == 3'h0;
  assign T143 = io_inner_acquire_bits_payload_subblock[3'h7:1'h0];
  assign T144 = {1'h0, T145};
  assign T145 = {1'h0, 1'h1};
  assign io_outer_finish_bits_payload_master_xact_id = outer_arb_io_out_finish_bits_payload_master_xact_id;
  assign io_outer_finish_bits_header_dst = outer_arb_io_out_finish_bits_header_dst;
  assign io_outer_finish_bits_header_src = outer_arb_io_out_finish_bits_header_src;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T75;
  assign T75 = {504'h0, outer_arb_io_out_acquire_bits_payload_subblock};
  assign io_outer_acquire_bits_payload_a_type = outer_arb_io_out_acquire_bits_payload_a_type;
  assign io_outer_acquire_bits_payload_uncached = outer_arb_io_out_acquire_bits_payload_uncached;
  assign io_outer_acquire_bits_payload_data = T0;
  assign T0 = is_in_sdq ? sdq_0 : T1;
  assign T1 = is_in_vwbdq ? vwbdq_0 : io_inner_release_bits_payload_data;
  assign T2 = T3 ? io_inner_release_bits_payload_data : vwbdq_0;
  assign T3 = T12 & T4;
  assign T4 = T5[1'h0:1'h0];
  assign T5 = 1'h1 << T6;
  assign T6 = T76;
  assign T76 = release_idx[1'h0:1'h0];
  assign T12 = voluntary & T13;
  assign T13 = io_inner_release_ready & io_inner_release_valid;
  assign is_in_vwbdq = outer_arb_io_out_acquire_bits_payload_data[1'h1:1'h1];
  assign T14 = T15 ? io_inner_acquire_bits_payload_data : sdq_0;
  assign T15 = sdq_enq & T16;
  assign T16 = T17[1'h0:1'h0];
  assign T17 = 1'h1 << T18;
  assign T18 = 1'h0;
  assign io_outer_acquire_bits_payload_client_xact_id = outer_arb_io_out_acquire_bits_payload_client_xact_id;
  assign io_outer_acquire_bits_payload_addr = outer_arb_io_out_acquire_bits_payload_addr;
  assign io_outer_acquire_bits_header_dst = outer_arb_io_out_acquire_bits_header_dst;
  assign io_outer_acquire_bits_header_src = outer_arb_io_out_acquire_bits_header_src;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T43;
  assign T43 = T57 ? T51 : T44;
  assign T44 = T50 ? T48 : T45;
  assign T45 = T46 ? AcquireTracker_0_io_inner_release_ready : VoluntaryReleaseTracker_io_inner_release_ready;
  assign T46 = T47[1'h0:1'h0];
  assign T47 = release_idx;
  assign T48 = T49 ? AcquireTracker_2_io_inner_release_ready : AcquireTracker_1_io_inner_release_ready;
  assign T49 = T47[1'h0:1'h0];
  assign T50 = T47[1'h1:1'h1];
  assign T51 = T56 ? T54 : T52;
  assign T52 = T53 ? AcquireTracker_4_io_inner_release_ready : AcquireTracker_3_io_inner_release_ready;
  assign T53 = T47[1'h0:1'h0];
  assign T54 = T55 ? AcquireTracker_6_io_inner_release_ready : AcquireTracker_5_io_inner_release_ready;
  assign T55 = T47[1'h0:1'h0];
  assign T56 = T47[1'h1:1'h1];
  assign T57 = T47[2'h2:2'h2];
  assign io_inner_probe_bits_payload_p_type = probe_arb_io_out_bits_payload_p_type;
  assign io_inner_probe_bits_payload_addr = probe_arb_io_out_bits_payload_addr;
  assign io_inner_probe_bits_header_dst = probe_arb_io_out_bits_header_dst;
  assign io_inner_probe_bits_header_src = probe_arb_io_out_bits_header_src;
  assign io_inner_probe_valid = probe_arb_io_out_valid;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_grant_bits_payload_g_type = grant_arb_io_out_bits_payload_g_type;
  assign io_inner_grant_bits_payload_uncached = grant_arb_io_out_bits_payload_uncached;
  assign io_inner_grant_bits_payload_master_xact_id = grant_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_grant_bits_payload_client_xact_id = grant_arb_io_out_bits_payload_client_xact_id;
  assign io_inner_grant_bits_payload_data = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = grant_arb_io_out_bits_header_dst;
  assign io_inner_grant_bits_header_src = grant_arb_io_out_bits_header_src;
  assign io_inner_grant_valid = grant_arb_io_out_valid;
  assign io_inner_acquire_ready = T58;
  assign T58 = T66 & T59;
  assign T59 = any_acquire_conflict ^ 1'h1;
  assign T66 = T68 & sdq_rdy;
  assign T68 = T69 | AcquireTracker_6_io_inner_acquire_ready;
  assign T69 = T70 | AcquireTracker_5_io_inner_acquire_ready;
  assign T70 = T71 | AcquireTracker_4_io_inner_acquire_ready;
  assign T71 = T72 | AcquireTracker_3_io_inner_acquire_ready;
  assign T72 = T73 | AcquireTracker_2_io_inner_acquire_ready;
  assign T73 = T74 | AcquireTracker_1_io_inner_acquire_ready;
  assign T74 = VoluntaryReleaseTracker_io_inner_acquire_ready | AcquireTracker_0_io_inner_acquire_ready;
  VoluntaryReleaseTracker VoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_0_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T144 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T143 ),
       .io_inner_grant_ready( grant_arb_io_in_0_ready ),
       .io_inner_grant_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( VoluntaryReleaseTracker_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_0_ready ),
       .io_inner_probe_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_header_src(  )
       //.io_inner_probe_bits_header_dst(  )
       //.io_inner_probe_bits_payload_addr(  )
       //.io_inner_probe_bits_payload_p_type(  )
       .io_inner_release_ready( VoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T141 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h2 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_0_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T140 ),
       .io_has_acquire_conflict( VoluntaryReleaseTracker_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_0 AcquireTracker_0(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_0_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_1_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T138 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T137 ),
       .io_inner_grant_ready( grant_arb_io_in_1_ready ),
       .io_inner_grant_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_0_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_1_ready ),
       .io_inner_probe_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_0_io_inner_release_ready ),
       .io_inner_release_valid( T135 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_0_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_0_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_1_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T134 ),
       .io_has_acquire_conflict( AcquireTracker_0_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_0_io_has_release_conflict )
  );
  AcquireTracker_1 AcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_2_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T132 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T131 ),
       .io_inner_grant_ready( grant_arb_io_in_2_ready ),
       .io_inner_grant_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_1_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_2_ready ),
       .io_inner_probe_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T129 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_1_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_1_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_2_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T128 ),
       .io_has_acquire_conflict( AcquireTracker_1_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_1_io_has_release_conflict )
  );
  AcquireTracker_2 AcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_3_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T126 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T125 ),
       .io_inner_grant_ready( grant_arb_io_in_3_ready ),
       .io_inner_grant_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_2_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_3_ready ),
       .io_inner_probe_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T123 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_2_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_2_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_3_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T122 ),
       .io_has_acquire_conflict( AcquireTracker_2_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_2_io_has_release_conflict )
  );
  AcquireTracker_3 AcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_4_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T120 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T119 ),
       .io_inner_grant_ready( grant_arb_io_in_4_ready ),
       .io_inner_grant_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_3_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_4_ready ),
       .io_inner_probe_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T117 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_3_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_3_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_4_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T116 ),
       .io_has_acquire_conflict( AcquireTracker_3_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_3_io_has_release_conflict )
  );
  AcquireTracker_4 AcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_5_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T114 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T113 ),
       .io_inner_grant_ready( grant_arb_io_in_5_ready ),
       .io_inner_grant_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_4_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_5_ready ),
       .io_inner_probe_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( T111 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_4_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_4_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_5_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T110 ),
       .io_has_acquire_conflict( AcquireTracker_4_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_4_io_has_release_conflict )
  );
  AcquireTracker_5 AcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_6_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T108 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T107 ),
       .io_inner_grant_ready( grant_arb_io_in_6_ready ),
       .io_inner_grant_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_5_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_6_ready ),
       .io_inner_probe_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( T105 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_5_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_5_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_6_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T104 ),
       .io_has_acquire_conflict( AcquireTracker_5_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_5_io_has_release_conflict )
  );
  AcquireTracker_6 AcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_7_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T102 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T101 ),
       .io_inner_grant_ready( grant_arb_io_in_7_ready ),
       .io_inner_grant_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_6_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_7_ready ),
       .io_inner_probe_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( T99 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( 3'h0 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_6_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_6_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_7_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T97 ),
       .io_has_acquire_conflict( AcquireTracker_6_io_has_acquire_conflict ),
       .io_has_release_conflict( AcquireTracker_6_io_has_release_conflict )
  );
  Arbiter_12 alloc_arb(
       .io_in_7_ready( alloc_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_acquire_ready ),
       //.io_in_7_bits(  )
       .io_in_6_ready( alloc_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_acquire_ready ),
       //.io_in_6_bits(  )
       .io_in_5_ready( alloc_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_acquire_ready ),
       //.io_in_5_bits(  )
       .io_in_4_ready( alloc_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_acquire_ready ),
       //.io_in_4_bits(  )
       .io_in_3_ready( alloc_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_acquire_ready ),
       //.io_in_3_bits(  )
       .io_in_2_ready( alloc_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_acquire_ready ),
       //.io_in_2_bits(  )
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_acquire_ready ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T94 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_7_bits = {1{$random}};
    assign alloc_arb.io_in_6_bits = {1{$random}};
    assign alloc_arb.io_in_5_bits = {1{$random}};
    assign alloc_arb.io_in_4_bits = {1{$random}};
    assign alloc_arb.io_in_3_bits = {1{$random}};
    assign alloc_arb.io_in_2_bits = {1{$random}};
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  Arbiter_13 probe_arb(
       .io_in_7_ready( probe_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_in_7_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_in_7_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_in_6_ready( probe_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_in_6_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_in_6_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_in_5_ready( probe_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_in_5_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_in_5_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_in_4_ready( probe_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_in_4_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_in_4_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_in_3_ready( probe_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_in_3_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_in_3_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_in_2_ready( probe_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_in_2_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_in_1_ready( probe_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_in_1_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_in_0_ready( probe_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_p_type(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( probe_arb_io_out_valid ),
       .io_out_bits_header_src( probe_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( probe_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( probe_arb_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( probe_arb_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign probe_arb.io_in_0_bits_header_src = {1{$random}};
    assign probe_arb.io_in_0_bits_header_dst = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_addr = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_p_type = {1{$random}};
  `endif
  Arbiter_14 grant_arb(
       .io_in_7_ready( grant_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_in_7_bits_payload_data( T93 ),
       .io_in_7_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_uncached( AcquireTracker_6_io_inner_grant_bits_payload_uncached ),
       .io_in_7_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       .io_in_6_ready( grant_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_in_6_bits_payload_data( T92 ),
       .io_in_6_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_uncached( AcquireTracker_5_io_inner_grant_bits_payload_uncached ),
       .io_in_6_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       .io_in_5_ready( grant_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_in_5_bits_payload_data( T91 ),
       .io_in_5_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_uncached( AcquireTracker_4_io_inner_grant_bits_payload_uncached ),
       .io_in_5_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       .io_in_4_ready( grant_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_in_4_bits_payload_data( T90 ),
       .io_in_4_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_uncached( AcquireTracker_3_io_inner_grant_bits_payload_uncached ),
       .io_in_4_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       .io_in_3_ready( grant_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_in_3_bits_payload_data( T89 ),
       .io_in_3_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_uncached( AcquireTracker_2_io_inner_grant_bits_payload_uncached ),
       .io_in_3_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       .io_in_2_ready( grant_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_in_2_bits_payload_data( T88 ),
       .io_in_2_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_uncached( AcquireTracker_1_io_inner_grant_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       .io_in_1_ready( grant_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_in_1_bits_payload_data( T87 ),
       .io_in_1_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_uncached( AcquireTracker_0_io_inner_grant_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       .io_in_0_ready( grant_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_in_0_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_in_0_bits_payload_data( T86 ),
       .io_in_0_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_uncached( VoluntaryReleaseTracker_io_inner_grant_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( grant_arb_io_out_valid ),
       .io_out_bits_header_src( grant_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( grant_arb_io_out_bits_header_dst ),
       //.io_out_bits_payload_data(  )
       .io_out_bits_payload_client_xact_id( grant_arb_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( grant_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_uncached( grant_arb_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( grant_arb_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  UncachedTileLinkIOArbiterThatPassesId outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_in_7_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_in_7_acquire_bits_header_dst(  )
       .io_in_7_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_in_7_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_7_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_in_7_acquire_bits_payload_uncached( AcquireTracker_6_io_outer_acquire_bits_payload_uncached ),
       .io_in_7_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_in_7_acquire_bits_payload_subblock( AcquireTracker_6_io_outer_acquire_bits_payload_subblock ),
       .io_in_7_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_in_7_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_in_7_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_in_7_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_in_7_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_in_7_grant_bits_payload_uncached( outer_arb_io_in_7_grant_bits_payload_uncached ),
       .io_in_7_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_in_7_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_in_7_finish_valid(  )
       //.io_in_7_finish_bits_header_src(  )
       //.io_in_7_finish_bits_header_dst(  )
       //.io_in_7_finish_bits_payload_master_xact_id(  )
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_in_6_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_in_6_acquire_bits_header_dst(  )
       .io_in_6_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_in_6_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_6_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_in_6_acquire_bits_payload_uncached( AcquireTracker_5_io_outer_acquire_bits_payload_uncached ),
       .io_in_6_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_in_6_acquire_bits_payload_subblock( AcquireTracker_5_io_outer_acquire_bits_payload_subblock ),
       .io_in_6_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_in_6_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_in_6_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_in_6_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_in_6_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_in_6_grant_bits_payload_uncached( outer_arb_io_in_6_grant_bits_payload_uncached ),
       .io_in_6_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_in_6_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_in_6_finish_valid(  )
       //.io_in_6_finish_bits_header_src(  )
       //.io_in_6_finish_bits_header_dst(  )
       //.io_in_6_finish_bits_payload_master_xact_id(  )
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_in_5_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_in_5_acquire_bits_header_dst(  )
       .io_in_5_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_in_5_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_5_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_in_5_acquire_bits_payload_uncached( AcquireTracker_4_io_outer_acquire_bits_payload_uncached ),
       .io_in_5_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_in_5_acquire_bits_payload_subblock( AcquireTracker_4_io_outer_acquire_bits_payload_subblock ),
       .io_in_5_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_in_5_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_in_5_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_in_5_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_in_5_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_in_5_grant_bits_payload_uncached( outer_arb_io_in_5_grant_bits_payload_uncached ),
       .io_in_5_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_in_5_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_in_5_finish_valid(  )
       //.io_in_5_finish_bits_header_src(  )
       //.io_in_5_finish_bits_header_dst(  )
       //.io_in_5_finish_bits_payload_master_xact_id(  )
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_in_4_acquire_bits_header_dst(  )
       .io_in_4_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_in_4_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_4_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_in_4_acquire_bits_payload_uncached( AcquireTracker_3_io_outer_acquire_bits_payload_uncached ),
       .io_in_4_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_in_4_acquire_bits_payload_subblock( AcquireTracker_3_io_outer_acquire_bits_payload_subblock ),
       .io_in_4_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_in_4_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_in_4_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_in_4_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_in_4_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_in_4_grant_bits_payload_uncached( outer_arb_io_in_4_grant_bits_payload_uncached ),
       .io_in_4_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_in_4_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_in_4_finish_valid(  )
       //.io_in_4_finish_bits_header_src(  )
       //.io_in_4_finish_bits_header_dst(  )
       //.io_in_4_finish_bits_payload_master_xact_id(  )
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_in_3_acquire_bits_header_dst(  )
       .io_in_3_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_in_3_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_3_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_in_3_acquire_bits_payload_uncached( AcquireTracker_2_io_outer_acquire_bits_payload_uncached ),
       .io_in_3_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_in_3_acquire_bits_payload_subblock( AcquireTracker_2_io_outer_acquire_bits_payload_subblock ),
       .io_in_3_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_in_3_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_in_3_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_in_3_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_in_3_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_in_3_grant_bits_payload_uncached( outer_arb_io_in_3_grant_bits_payload_uncached ),
       .io_in_3_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_in_3_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_in_3_finish_valid(  )
       //.io_in_3_finish_bits_header_src(  )
       //.io_in_3_finish_bits_header_dst(  )
       //.io_in_3_finish_bits_payload_master_xact_id(  )
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_in_2_acquire_bits_header_dst(  )
       .io_in_2_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_uncached( AcquireTracker_1_io_outer_acquire_bits_payload_uncached ),
       .io_in_2_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_subblock( AcquireTracker_1_io_outer_acquire_bits_payload_subblock ),
       .io_in_2_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_in_2_grant_bits_payload_uncached( outer_arb_io_in_2_grant_bits_payload_uncached ),
       .io_in_2_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_in_2_finish_valid(  )
       //.io_in_2_finish_bits_header_src(  )
       //.io_in_2_finish_bits_header_dst(  )
       //.io_in_2_finish_bits_payload_master_xact_id(  )
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_uncached( AcquireTracker_0_io_outer_acquire_bits_payload_uncached ),
       .io_in_1_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_subblock( AcquireTracker_0_io_outer_acquire_bits_payload_subblock ),
       .io_in_1_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_uncached( outer_arb_io_in_1_grant_bits_payload_uncached ),
       .io_in_1_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_in_1_finish_valid(  )
       //.io_in_1_finish_bits_header_src(  )
       //.io_in_1_finish_bits_header_dst(  )
       //.io_in_1_finish_bits_payload_master_xact_id(  )
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_in_0_acquire_bits_header_dst(  )
       .io_in_0_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_uncached( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_uncached ),
       .io_in_0_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_subblock( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subblock ),
       .io_in_0_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_uncached( outer_arb_io_in_0_grant_bits_payload_uncached ),
       .io_in_0_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_in_0_finish_valid(  )
       //.io_in_0_finish_bits_header_src(  )
       //.io_in_0_finish_bits_header_dst(  )
       //.io_in_0_finish_bits_payload_master_xact_id(  )
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( outer_arb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( outer_arb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( outer_arb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( outer_arb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( outer_arb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_uncached( outer_arb_io_out_acquire_bits_payload_uncached ),
       .io_out_acquire_bits_payload_a_type( outer_arb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_subblock( outer_arb_io_out_acquire_bits_payload_subblock ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_header_src( io_outer_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_outer_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( T85 ),
       .io_out_grant_bits_payload_client_xact_id( io_outer_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_outer_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_uncached( io_outer_grant_bits_payload_uncached ),
       .io_out_grant_bits_payload_g_type( io_outer_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_outer_finish_ready ),
       .io_out_finish_valid( outer_arb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( outer_arb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( outer_arb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( outer_arb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign outer_arb.io_in_7_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_valid = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_6_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_valid = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_5_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_valid = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_4_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_valid = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_valid = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_valid = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_valid = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_valid = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_payload_master_xact_id = {1{$random}};
  `endif

  always @(posedge clk) begin
    sdq_val <= T79;
    if(T3) begin
      vwbdq_0 <= io_inner_release_bits_payload_data;
    end
    if(T15) begin
      sdq_0 <= io_inner_acquire_bits_payload_data;
    end
  end
endmodule

module Queue_18(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[5:0] T15;
  wire[4:0] T16;
  wire[25:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_rw = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_addr, T15};
  assign T15 = {io_enq_bits_tag, io_enq_bits_rw};
  assign io_deq_bits_tag = T16;
  assign T16 = T11[3'h5:1'h1];
  assign io_deq_bits_addr = T17;
  assign T17 = T11[5'h1f:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_19(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T16;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T17;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T18;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[127:0] T11;
  reg [127:0] ram [1:0];
  wire[127:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T16 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T17 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T18 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_data;
  end
endmodule

module MemIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [2:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input  io_uncached_acquire_bits_payload_uncached,
    input [1:0] io_uncached_acquire_bits_payload_a_type,
    input [511:0] io_uncached_acquire_bits_payload_subblock,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[2:0] io_uncached_grant_bits_payload_client_xact_id,
    output io_uncached_grant_bits_payload_master_xact_id,
    output io_uncached_grant_bits_payload_uncached,
    output[1:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input  io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire[127:0] T56;
  reg [511:0] buf_out;
  wire[511:0] T57;
  wire[511:0] T58;
  wire T30;
  wire T31;
  reg  active_out;
  wire T53;
  wire T28;
  wire T29;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [2:0] cnt_out;
  wire[2:0] T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire T41;
  reg  has_data;
  wire T54;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg  cmd_sent_out;
  wire T55;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[511:0] T59;
  wire[383:0] T60;
  wire T39;
  wire T40;
  wire T61;
  wire T62;
  wire T63;
  wire[4:0] T64;
  reg [2:0] tag_out;
  wire[2:0] T65;
  reg [25:0] addr_out;
  wire[25:0] T66;
  wire T67;
  wire T68;
  wire T0;
  wire T1;
  reg [2:0] cnt_in;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  wire T5;
  reg  active_in;
  wire T51;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire[2:0] T17;
  wire[2:0] T52;
  reg [4:0] tag_in;
  wire[4:0] T18;
  wire[511:0] T19;
  reg [511:0] buf_in;
  wire[511:0] T20;
  wire[511:0] T21;
  wire[511:0] T22;
  wire[511:0] T23;
  wire[383:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire mem_cmd_q_io_enq_ready;
  wire mem_cmd_q_io_deq_valid;
  wire[25:0] mem_cmd_q_io_deq_bits_addr;
  wire[4:0] mem_cmd_q_io_deq_bits_tag;
  wire mem_cmd_q_io_deq_bits_rw;
  wire mem_data_q_io_enq_ready;
  wire mem_data_q_io_deq_valid;
  wire[127:0] mem_data_q_io_deq_bits_data;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    buf_out = {16{$random}};
    active_out = {1{$random}};
    cnt_out = {1{$random}};
    has_data = {1{$random}};
    cmd_sent_out = {1{$random}};
    tag_out = {1{$random}};
    addr_out = {1{$random}};
    cnt_in = {1{$random}};
    active_in = {1{$random}};
    tag_in = {1{$random}};
    buf_in = {16{$random}};
  end
`endif

  assign T56 = buf_out[7'h7f:1'h0];
  assign T57 = T39 ? T59 : T58;
  assign T58 = T30 ? io_uncached_acquire_bits_payload_data : buf_out;
  assign T30 = T31 & io_uncached_acquire_valid;
  assign T31 = active_out ^ 1'h1;
  assign T53 = reset ? 1'h0 : T28;
  assign T28 = T32 ? 1'h0 : T29;
  assign T29 = T30 ? 1'h1 : active_out;
  assign T32 = active_out & T33;
  assign T33 = cmd_sent_out & T34;
  assign T34 = T41 | T35;
  assign T35 = cnt_out == 3'h4;
  assign T36 = T39 ? T38 : T37;
  assign T37 = T30 ? 3'h0 : cnt_out;
  assign T38 = cnt_out + 3'h1;
  assign T41 = has_data ^ 1'h1;
  assign T54 = reset ? 1'h0 : T42;
  assign T42 = T30 ? T43 : has_data;
  assign T43 = io_uncached_acquire_bits_payload_uncached ? T44 : 1'h0;
  assign T44 = T46 | T45;
  assign T45 = 2'h2 == io_uncached_acquire_bits_payload_a_type;
  assign T46 = 2'h1 == io_uncached_acquire_bits_payload_a_type;
  assign T55 = reset ? 1'h0 : T47;
  assign T47 = T49 ? 1'h1 : T48;
  assign T48 = T30 ? 1'h0 : cmd_sent_out;
  assign T49 = active_out & T50;
  assign T50 = mem_cmd_q_io_enq_ready & T67;
  assign T59 = {128'h0, T60};
  assign T60 = buf_out >> 8'h80;
  assign T39 = active_out & T40;
  assign T40 = mem_data_q_io_enq_ready & T61;
  assign T61 = T63 & T62;
  assign T62 = cnt_out < 3'h4;
  assign T63 = active_out & has_data;
  assign T64 = {2'h0, tag_out};
  assign T65 = T30 ? io_uncached_acquire_bits_payload_client_xact_id : tag_out;
  assign T66 = T30 ? io_uncached_acquire_bits_payload_addr : addr_out;
  assign T67 = active_out & T68;
  assign T68 = cmd_sent_out ^ 1'h1;
  assign io_mem_resp_ready = T0;
  assign T0 = T13 | T1;
  assign T1 = cnt_in < 3'h4;
  assign T2 = T11 ? T10 : T3;
  assign T3 = T4 ? 3'h1 : cnt_in;
  assign T4 = T5 & io_mem_resp_valid;
  assign T5 = active_in ^ 1'h1;
  assign T51 = reset ? 1'h0 : T6;
  assign T6 = T8 ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : active_in;
  assign T8 = active_in & T9;
  assign T9 = io_uncached_grant_ready & io_uncached_grant_valid;
  assign T10 = cnt_in + 3'h1;
  assign T11 = active_in & T12;
  assign T12 = io_mem_resp_ready & io_mem_resp_valid;
  assign T13 = active_in ^ 1'h1;
  assign io_mem_req_data_bits_data = mem_data_q_io_deq_bits_data;
  assign io_mem_req_data_valid = mem_data_q_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = mem_cmd_q_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = mem_cmd_q_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = mem_cmd_q_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = mem_cmd_q_io_deq_valid;
  assign io_uncached_grant_bits_payload_g_type = T14;
  assign T14 = 2'h0;
  assign io_uncached_grant_bits_payload_uncached = T15;
  assign T15 = 1'h1;
  assign io_uncached_grant_bits_payload_master_xact_id = T16;
  assign T16 = 1'h0;
  assign io_uncached_grant_bits_payload_client_xact_id = T17;
  assign T17 = T52;
  assign T52 = tag_in[2'h2:1'h0];
  assign T18 = T4 ? io_mem_resp_bits_tag : tag_in;
  assign io_uncached_grant_bits_payload_data = T19;
  assign T19 = buf_in;
  assign T20 = T11 ? T23 : T21;
  assign T21 = T4 ? T22 : buf_in;
  assign T22 = io_mem_resp_bits_data << 9'h180;
  assign T23 = {io_mem_resp_bits_data, T24};
  assign T24 = buf_in[9'h1ff:8'h80];
  assign io_uncached_grant_valid = T25;
  assign T25 = active_in & T26;
  assign T26 = cnt_in == 3'h4;
  assign io_uncached_acquire_ready = T27;
  assign T27 = active_out ^ 1'h1;
  Queue_18 mem_cmd_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_cmd_q_io_enq_ready ),
       .io_enq_valid( T67 ),
       .io_enq_bits_addr( addr_out ),
       .io_enq_bits_tag( T64 ),
       .io_enq_bits_rw( has_data ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( mem_cmd_q_io_deq_valid ),
       .io_deq_bits_addr( mem_cmd_q_io_deq_bits_addr ),
       .io_deq_bits_tag( mem_cmd_q_io_deq_bits_tag ),
       .io_deq_bits_rw( mem_cmd_q_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_19 mem_data_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_data_q_io_enq_ready ),
       .io_enq_valid( T61 ),
       .io_enq_bits_data( T56 ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( mem_data_q_io_deq_valid ),
       .io_deq_bits_data( mem_data_q_io_deq_bits_data )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T39) begin
      buf_out <= T59;
    end else if(T30) begin
      buf_out <= io_uncached_acquire_bits_payload_data;
    end
    if(reset) begin
      active_out <= 1'h0;
    end else if(T32) begin
      active_out <= 1'h0;
    end else if(T30) begin
      active_out <= 1'h1;
    end
    if(T39) begin
      cnt_out <= T38;
    end else if(T30) begin
      cnt_out <= 3'h0;
    end
    if(reset) begin
      has_data <= 1'h0;
    end else if(T30) begin
      has_data <= T43;
    end
    if(reset) begin
      cmd_sent_out <= 1'h0;
    end else if(T49) begin
      cmd_sent_out <= 1'h1;
    end else if(T30) begin
      cmd_sent_out <= 1'h0;
    end
    if(T30) begin
      tag_out <= io_uncached_acquire_bits_payload_client_xact_id;
    end
    if(T30) begin
      addr_out <= io_uncached_acquire_bits_payload_addr;
    end
    if(T11) begin
      cnt_in <= T10;
    end else if(T4) begin
      cnt_in <= 3'h1;
    end
    if(reset) begin
      active_in <= 1'h0;
    end else if(T8) begin
      active_in <= 1'h0;
    end else if(T4) begin
      active_in <= 1'h1;
    end
    if(T4) begin
      tag_in <= io_mem_resp_bits_tag;
    end
    if(T11) begin
      buf_in <= T23;
    end else if(T4) begin
      buf_in <= T22;
    end
  end
endmodule

module HellaFlowQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[6:0] io_count
);

  wire[4:0] T0;
  wire[4:0] T1;
  wire[132:0] T2;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire atLeastTwo;
  wire T23;
  wire[5:0] T24;
  reg [5:0] deq_ptr;
  wire[5:0] T32;
  wire[5:0] T13;
  wire[5:0] T14;
  wire do_deq;
  wire T15;
  wire do_flow;
  wire T7;
  wire T16;
  reg [5:0] enq_ptr;
  wire[5:0] T33;
  wire[5:0] T9;
  wire[5:0] T10;
  wire do_enq;
  wire T6;
  wire T8;
  wire full;
  reg  maybe_full;
  wire T34;
  wire T25;
  wire T26;
  wire ptr_match;
  wire[5:0] T12;
  wire[5:0] T17;
  wire[132:0] T3;
  wire[132:0] T4;
  wire[132:0] T5;
  reg [5:0] ram_addr;
  wire[5:0] T11;
  wire empty;
  wire T27;
  wire[127:0] T28;
  wire[127:0] T29;
  wire T30;
  reg  ram_out_valid;
  wire T31;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    ram_addr = {1{$random}};
    ram_out_valid = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = empty ? io_enq_bits_tag : T1;
  assign T1 = T2[3'h4:1'h0];
  assign T18 = io_deq_ready & T19;
  assign T19 = atLeastTwo | T20;
  assign T20 = T22 & T21;
  assign T21 = empty ^ 1'h1;
  assign T22 = io_deq_valid ^ 1'h1;
  assign atLeastTwo = full | T23;
  assign T23 = 6'h2 <= T24;
  assign T24 = enq_ptr - deq_ptr;
  assign T32 = reset ? 6'h0 : T13;
  assign T13 = do_deq ? T14 : deq_ptr;
  assign T14 = deq_ptr + 6'h1;
  assign do_deq = T16 & T15;
  assign T15 = do_flow ^ 1'h1;
  assign do_flow = T7;
  assign T7 = empty & io_deq_ready;
  assign T16 = io_deq_ready & io_deq_valid;
  assign T33 = reset ? 6'h0 : T9;
  assign T9 = do_enq ? T10 : enq_ptr;
  assign T10 = enq_ptr + 6'h1;
  assign do_enq = T8 & T6;
  assign T6 = do_flow ^ 1'h1;
  assign T8 = io_enq_ready & io_enq_valid;
  assign full = ptr_match & maybe_full;
  assign T34 = reset ? 1'h0 : T25;
  assign T25 = T26 ? do_enq : maybe_full;
  assign T26 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = io_deq_valid ? T17 : deq_ptr;
  assign T17 = deq_ptr + 6'h1;
  HellaFlowQueue_ram ram (
    .CLK(clk),
    .W0A(enq_ptr),
    .W0E(do_enq),
    .W0I(T4),
    .R1A(T12),
    .R1E(T18),
    .R1O(T2)
  );
  assign T4 = T5;
  assign T5 = {io_enq_bits_data, io_enq_bits_tag};
  assign T11 = T18 ? T12 : ram_addr;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_deq_bits_data = T28;
  assign T28 = empty ? io_enq_bits_data : T29;
  assign T29 = T2[8'h84:3'h5];
  assign io_deq_valid = T30;
  assign T30 = empty ? io_enq_valid : ram_out_valid;
  assign io_enq_ready = T31;
  assign T31 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 6'h0;
    end else if(do_deq) begin
      deq_ptr <= T14;
    end
    if(reset) begin
      enq_ptr <= 6'h0;
    end else if(do_enq) begin
      enq_ptr <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T26) begin
      maybe_full <= do_enq;
    end
    if(T18) begin
      ram_addr <= T12;
    end
    ram_out_valid <= T18;
  end
endmodule

module Queue_20(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
);

  wire[4:0] T0;
  wire[132:0] T1;
  reg [132:0] ram [0:0];
  wire[132:0] T2;
  wire[132:0] T3;
  wire[132:0] T4;
  wire do_enq;
  wire[127:0] T5;
  wire T6;
  wire empty;
  reg  full;
  wire T11;
  wire T7;
  wire T8;
  wire do_deq;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {5{$random}};
    full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[3'h4:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {io_enq_bits_data, io_enq_bits_tag};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_data = T5;
  assign T5 = T1[8'h84:3'h5];
  assign io_deq_valid = T6;
  assign T6 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign T11 = reset ? 1'h0 : T7;
  assign T7 = T8 ? do_enq : full;
  assign T8 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T9;
  assign T9 = T10 | io_deq_ready;
  assign T10 = full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      full <= 1'h0;
    end else if(T8) begin
      full <= do_enq;
    end
  end
endmodule

module HellaQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[6:0] io_count
);

  wire fq_io_enq_ready;
  wire fq_io_deq_valid;
  wire[127:0] fq_io_deq_bits_data;
  wire[4:0] fq_io_deq_bits_tag;
  wire Queue_20_io_enq_ready;
  wire Queue_20_io_deq_valid;
  wire[127:0] Queue_20_io_deq_bits_data;
  wire[4:0] Queue_20_io_deq_bits_tag;


  assign io_deq_bits_tag = Queue_20_io_deq_bits_tag;
  assign io_deq_bits_data = Queue_20_io_deq_bits_data;
  assign io_deq_valid = Queue_20_io_deq_valid;
  assign io_enq_ready = fq_io_enq_ready;
  HellaFlowQueue fq(.clk(clk), .reset(reset),
       .io_enq_ready( fq_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_data( io_enq_bits_data ),
       .io_enq_bits_tag( io_enq_bits_tag ),
       .io_deq_ready( Queue_20_io_enq_ready ),
       .io_deq_valid( fq_io_deq_valid ),
       .io_deq_bits_data( fq_io_deq_bits_data ),
       .io_deq_bits_tag( fq_io_deq_bits_tag )
       //.io_count(  )
  );
  Queue_20 Queue_20(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_20_io_enq_ready ),
       .io_enq_valid( fq_io_deq_valid ),
       .io_enq_bits_data( fq_io_deq_bits_data ),
       .io_enq_bits_tag( fq_io_deq_bits_tag ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( Queue_20_io_deq_valid ),
       .io_deq_bits_data( Queue_20_io_deq_bits_data ),
       .io_deq_bits_tag( Queue_20_io_deq_bits_tag )
  );
endmodule

module MemPipeIOMemIOConverter(input clk, input reset,
    output io_cpu_req_cmd_ready,
    input  io_cpu_req_cmd_valid,
    input [25:0] io_cpu_req_cmd_bits_addr,
    input [4:0] io_cpu_req_cmd_bits_tag,
    input  io_cpu_req_cmd_bits_rw,
    output io_cpu_req_data_ready,
    input  io_cpu_req_data_valid,
    input [127:0] io_cpu_req_data_bits_data,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[127:0] io_cpu_resp_bits_data,
    output[4:0] io_cpu_resp_bits_tag,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire T0;
  wire cmdq_mask;
  wire watermark;
  reg [6:0] count;
  wire[6:0] T17;
  wire[6:0] T1;
  wire[6:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire T5;
  wire T6;
  wire dec;
  wire T7;
  wire T8;
  wire T9;
  wire inc;
  wire T10;
  wire[6:0] T11;
  wire T12;
  wire T13;
  wire[6:0] T14;
  wire T15;
  wire T16;
  wire resp_dataq_io_deq_valid;
  wire[127:0] resp_dataq_io_deq_bits_data;
  wire[4:0] resp_dataq_io_deq_bits_tag;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    count = {1{$random}};
  end
`endif

  assign io_mem_req_data_bits_data = io_cpu_req_data_bits_data;
  assign io_mem_req_data_valid = io_cpu_req_data_valid;
  assign io_mem_req_cmd_bits_rw = io_cpu_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = io_cpu_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = io_cpu_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = T0;
  assign T0 = io_cpu_req_cmd_valid & cmdq_mask;
  assign cmdq_mask = io_cpu_req_cmd_bits_rw | watermark;
  assign watermark = 7'h4 <= count;
  assign T17 = reset ? 7'h40 : T1;
  assign T1 = T15 ? T14 : T2;
  assign T2 = T12 ? T11 : T3;
  assign T3 = T5 ? T4 : count;
  assign T4 = count + 7'h1;
  assign T5 = inc & T6;
  assign T6 = dec ^ 1'h1;
  assign dec = T7;
  assign T7 = T9 & T8;
  assign T8 = io_mem_req_cmd_bits_rw ^ 1'h1;
  assign T9 = io_mem_req_cmd_ready & io_mem_req_cmd_valid;
  assign inc = T10;
  assign T10 = io_cpu_resp_ready & resp_dataq_io_deq_valid;
  assign T11 = count - 7'h4;
  assign T12 = T13 & dec;
  assign T13 = inc ^ 1'h1;
  assign T14 = count - 7'h3;
  assign T15 = inc & dec;
  assign io_cpu_resp_bits_tag = resp_dataq_io_deq_bits_tag;
  assign io_cpu_resp_bits_data = resp_dataq_io_deq_bits_data;
  assign io_cpu_resp_valid = resp_dataq_io_deq_valid;
  assign io_cpu_req_data_ready = io_mem_req_data_ready;
  assign io_cpu_req_cmd_ready = T16;
  assign T16 = io_mem_req_cmd_ready & cmdq_mask;
  HellaQueue resp_dataq(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_data( io_mem_resp_bits_data ),
       .io_enq_bits_tag( io_mem_resp_bits_tag ),
       .io_deq_ready( io_cpu_resp_ready ),
       .io_deq_valid( resp_dataq_io_deq_valid ),
       .io_deq_bits_data( resp_dataq_io_deq_bits_data ),
       .io_deq_bits_tag( resp_dataq_io_deq_bits_tag )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      count <= 7'h40;
    end else if(T15) begin
      count <= T14;
    end else if(T12) begin
      count <= T11;
    end else if(T5) begin
      count <= T4;
    end
  end
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] ram [1:0];
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[5:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[4:0] T12;
  wire[25:0] T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_rw = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_addr, T5};
  assign T5 = {io_enq_bits_tag, io_enq_bits_rw};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_tag = T12;
  assign T12 = T1[3'h5:1'h1];
  assign io_deq_bits_addr = T13;
  assign T13 = T1[5'h1f:3'h6];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_16(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
);

  wire[127:0] T0;
  wire[127:0] T1;
  reg [127:0] ram [3:0];
  wire[127:0] T2;
  wire do_enq;
  reg [1:0] R3;
  wire[1:0] T14;
  wire[1:0] T4;
  wire[1:0] T5;
  reg [1:0] R6;
  wire[1:0] T15;
  wire[1:0] T7;
  wire[1:0] T8;
  wire do_deq;
  wire T9;
  wire empty;
  wire T10;
  reg  maybe_full;
  wire T16;
  wire T11;
  wire T12;
  wire ptr_match;
  wire T13;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {4{$random}};
    R3 = {1{$random}};
    R6 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[7'h7f:1'h0];
  assign T1 = ram[R6];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T14 = reset ? 2'h0 : T4;
  assign T4 = do_enq ? T5 : R3;
  assign T5 = R3 + 2'h1;
  assign T15 = reset ? 2'h0 : T7;
  assign T7 = do_deq ? T8 : R6;
  assign T8 = R6 + 2'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T9;
  assign T9 = empty ^ 1'h1;
  assign empty = ptr_match & T10;
  assign T10 = maybe_full ^ 1'h1;
  assign T16 = reset ? 1'h0 : T11;
  assign T11 = T12 ? do_enq : maybe_full;
  assign T12 = do_enq != do_deq;
  assign ptr_match = R3 == R6;
  assign io_enq_ready = T13;
  assign T13 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R3] <= io_enq_bits_data;
    if(reset) begin
      R3 <= 2'h0;
    end else if(do_enq) begin
      R3 <= T5;
    end
    if(reset) begin
      R6 <= 2'h0;
    end else if(do_deq) begin
      R6 <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T12) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module MemPipeIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [2:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input  io_uncached_acquire_bits_payload_uncached,
    input [1:0] io_uncached_acquire_bits_payload_a_type,
    input [511:0] io_uncached_acquire_bits_payload_subblock,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[2:0] io_uncached_grant_bits_payload_client_xact_id,
    output io_uncached_grant_bits_payload_master_xact_id,
    output io_uncached_grant_bits_payload_uncached,
    output[1:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input  io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire Queue_18_io_enq_ready;
  wire Queue_18_io_deq_valid;
  wire[25:0] Queue_18_io_deq_bits_addr;
  wire[4:0] Queue_18_io_deq_bits_tag;
  wire Queue_18_io_deq_bits_rw;
  wire Queue_19_io_enq_ready;
  wire Queue_19_io_deq_valid;
  wire[127:0] Queue_19_io_deq_bits_data;
  wire a_io_uncached_acquire_ready;
  wire a_io_uncached_grant_valid;
  wire[511:0] a_io_uncached_grant_bits_payload_data;
  wire[2:0] a_io_uncached_grant_bits_payload_client_xact_id;
  wire a_io_uncached_grant_bits_payload_master_xact_id;
  wire a_io_uncached_grant_bits_payload_uncached;
  wire[1:0] a_io_uncached_grant_bits_payload_g_type;
  wire a_io_mem_req_cmd_valid;
  wire[25:0] a_io_mem_req_cmd_bits_addr;
  wire[4:0] a_io_mem_req_cmd_bits_tag;
  wire a_io_mem_req_cmd_bits_rw;
  wire a_io_mem_req_data_valid;
  wire[127:0] a_io_mem_req_data_bits_data;
  wire a_io_mem_resp_ready;
  wire b_io_cpu_req_cmd_ready;
  wire b_io_cpu_req_data_ready;
  wire b_io_cpu_resp_valid;
  wire[127:0] b_io_cpu_resp_bits_data;
  wire[4:0] b_io_cpu_resp_bits_tag;
  wire b_io_mem_req_cmd_valid;
  wire[25:0] b_io_mem_req_cmd_bits_addr;
  wire[4:0] b_io_mem_req_cmd_bits_tag;
  wire b_io_mem_req_cmd_bits_rw;
  wire b_io_mem_req_data_valid;
  wire[127:0] b_io_mem_req_data_bits_data;


  assign io_mem_req_data_bits_data = b_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = b_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = b_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = b_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = b_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = b_io_mem_req_cmd_valid;
  assign io_uncached_grant_bits_payload_g_type = a_io_uncached_grant_bits_payload_g_type;
  assign io_uncached_grant_bits_payload_uncached = a_io_uncached_grant_bits_payload_uncached;
  assign io_uncached_grant_bits_payload_master_xact_id = a_io_uncached_grant_bits_payload_master_xact_id;
  assign io_uncached_grant_bits_payload_client_xact_id = a_io_uncached_grant_bits_payload_client_xact_id;
  assign io_uncached_grant_bits_payload_data = a_io_uncached_grant_bits_payload_data;
  assign io_uncached_grant_valid = a_io_uncached_grant_valid;
  assign io_uncached_acquire_ready = a_io_uncached_acquire_ready;
  MemIOUncachedTileLinkIOConverter a(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( a_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( io_uncached_acquire_valid ),
       .io_uncached_acquire_bits_header_src( io_uncached_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( io_uncached_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( io_uncached_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( io_uncached_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( io_uncached_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_uncached( io_uncached_acquire_bits_payload_uncached ),
       .io_uncached_acquire_bits_payload_a_type( io_uncached_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_subblock( io_uncached_acquire_bits_payload_subblock ),
       .io_uncached_grant_ready( io_uncached_grant_ready ),
       .io_uncached_grant_valid( a_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( a_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( a_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( a_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_uncached( a_io_uncached_grant_bits_payload_uncached ),
       .io_uncached_grant_bits_payload_g_type( a_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( io_uncached_finish_valid ),
       .io_uncached_finish_bits_header_src( io_uncached_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( io_uncached_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( io_uncached_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( Queue_18_io_enq_ready ),
       .io_mem_req_cmd_valid( a_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( a_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( a_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( a_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( Queue_19_io_enq_ready ),
       .io_mem_req_data_valid( a_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( a_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( a_io_mem_resp_ready ),
       .io_mem_resp_valid( b_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( b_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_tag( b_io_cpu_resp_bits_tag )
  );
  MemPipeIOMemIOConverter b(.clk(clk), .reset(reset),
       .io_cpu_req_cmd_ready( b_io_cpu_req_cmd_ready ),
       .io_cpu_req_cmd_valid( Queue_18_io_deq_valid ),
       .io_cpu_req_cmd_bits_addr( Queue_18_io_deq_bits_addr ),
       .io_cpu_req_cmd_bits_tag( Queue_18_io_deq_bits_tag ),
       .io_cpu_req_cmd_bits_rw( Queue_18_io_deq_bits_rw ),
       .io_cpu_req_data_ready( b_io_cpu_req_data_ready ),
       .io_cpu_req_data_valid( Queue_19_io_deq_valid ),
       .io_cpu_req_data_bits_data( Queue_19_io_deq_bits_data ),
       .io_cpu_resp_ready( a_io_mem_resp_ready ),
       .io_cpu_resp_valid( b_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( b_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_tag( b_io_cpu_resp_bits_tag ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( b_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( b_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( b_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( b_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( b_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( b_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
  Queue_15 Queue_18(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_18_io_enq_ready ),
       .io_enq_valid( a_io_mem_req_cmd_valid ),
       .io_enq_bits_addr( a_io_mem_req_cmd_bits_addr ),
       .io_enq_bits_tag( a_io_mem_req_cmd_bits_tag ),
       .io_enq_bits_rw( a_io_mem_req_cmd_bits_rw ),
       .io_deq_ready( b_io_cpu_req_cmd_ready ),
       .io_deq_valid( Queue_18_io_deq_valid ),
       .io_deq_bits_addr( Queue_18_io_deq_bits_addr ),
       .io_deq_bits_tag( Queue_18_io_deq_bits_tag ),
       .io_deq_bits_rw( Queue_18_io_deq_bits_rw )
  );
  Queue_16 Queue_19(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_19_io_enq_ready ),
       .io_enq_valid( a_io_mem_req_data_valid ),
       .io_enq_bits_data( a_io_mem_req_data_bits_data ),
       .io_deq_ready( b_io_cpu_req_data_ready ),
       .io_deq_valid( Queue_19_io_deq_valid ),
       .io_deq_bits_data( Queue_19_io_deq_bits_data )
  );
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [2:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input  io_tiles_0_acquire_bits_payload_uncached,
    input [1:0] io_tiles_0_acquire_bits_payload_a_type,
    input [511:0] io_tiles_0_acquire_bits_payload_subblock,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[2:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output io_tiles_0_grant_bits_payload_uncached,
    output[1:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [2:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_acquire_ready,
    input  io_htif_acquire_valid,
    input [1:0] io_htif_acquire_bits_header_src,
    input [1:0] io_htif_acquire_bits_header_dst,
    input [25:0] io_htif_acquire_bits_payload_addr,
    input [2:0] io_htif_acquire_bits_payload_client_xact_id,
    input [511:0] io_htif_acquire_bits_payload_data,
    input  io_htif_acquire_bits_payload_uncached,
    input [1:0] io_htif_acquire_bits_payload_a_type,
    input [511:0] io_htif_acquire_bits_payload_subblock,
    input  io_htif_grant_ready,
    output io_htif_grant_valid,
    output[1:0] io_htif_grant_bits_header_src,
    output[1:0] io_htif_grant_bits_header_dst,
    output[511:0] io_htif_grant_bits_payload_data,
    output[2:0] io_htif_grant_bits_payload_client_xact_id,
    output[2:0] io_htif_grant_bits_payload_master_xact_id,
    output io_htif_grant_bits_payload_uncached,
    output[1:0] io_htif_grant_bits_payload_g_type,
    output io_htif_finish_ready,
    input  io_htif_finish_valid,
    input [1:0] io_htif_finish_bits_header_src,
    input [1:0] io_htif_finish_bits_header_dst,
    input [2:0] io_htif_finish_bits_payload_master_xact_id,
    input  io_htif_probe_ready,
    output io_htif_probe_valid,
    output[1:0] io_htif_probe_bits_header_src,
    output[1:0] io_htif_probe_bits_header_dst,
    output[25:0] io_htif_probe_bits_payload_addr,
    output[1:0] io_htif_probe_bits_payload_p_type,
    output io_htif_release_ready,
    input  io_htif_release_valid,
    input [1:0] io_htif_release_bits_header_src,
    input [1:0] io_htif_release_bits_header_dst,
    input [25:0] io_htif_release_bits_payload_addr,
    input [2:0] io_htif_release_bits_payload_client_xact_id,
    input [511:0] io_htif_release_bits_payload_data,
    input [2:0] io_htif_release_bits_payload_r_type,
    input  io_incoherent_1,
    input  io_incoherent_0,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire net_io_clients_1_acquire_ready;
  wire net_io_clients_1_grant_valid;
  wire[1:0] net_io_clients_1_grant_bits_header_src;
  wire[1:0] net_io_clients_1_grant_bits_header_dst;
  wire[511:0] net_io_clients_1_grant_bits_payload_data;
  wire[2:0] net_io_clients_1_grant_bits_payload_client_xact_id;
  wire[2:0] net_io_clients_1_grant_bits_payload_master_xact_id;
  wire net_io_clients_1_grant_bits_payload_uncached;
  wire[1:0] net_io_clients_1_grant_bits_payload_g_type;
  wire net_io_clients_1_finish_ready;
  wire net_io_clients_1_probe_valid;
  wire[1:0] net_io_clients_1_probe_bits_header_src;
  wire[1:0] net_io_clients_1_probe_bits_header_dst;
  wire[25:0] net_io_clients_1_probe_bits_payload_addr;
  wire[1:0] net_io_clients_1_probe_bits_payload_p_type;
  wire net_io_clients_1_release_ready;
  wire net_io_clients_0_acquire_ready;
  wire net_io_clients_0_grant_valid;
  wire[1:0] net_io_clients_0_grant_bits_header_src;
  wire[1:0] net_io_clients_0_grant_bits_header_dst;
  wire[511:0] net_io_clients_0_grant_bits_payload_data;
  wire[2:0] net_io_clients_0_grant_bits_payload_client_xact_id;
  wire[2:0] net_io_clients_0_grant_bits_payload_master_xact_id;
  wire net_io_clients_0_grant_bits_payload_uncached;
  wire[1:0] net_io_clients_0_grant_bits_payload_g_type;
  wire net_io_clients_0_finish_ready;
  wire net_io_clients_0_probe_valid;
  wire[1:0] net_io_clients_0_probe_bits_header_src;
  wire[1:0] net_io_clients_0_probe_bits_header_dst;
  wire[25:0] net_io_clients_0_probe_bits_payload_addr;
  wire[1:0] net_io_clients_0_probe_bits_payload_p_type;
  wire net_io_clients_0_release_ready;
  wire net_io_masters_0_acquire_valid;
  wire[1:0] net_io_masters_0_acquire_bits_header_src;
  wire[1:0] net_io_masters_0_acquire_bits_header_dst;
  wire[25:0] net_io_masters_0_acquire_bits_payload_addr;
  wire[2:0] net_io_masters_0_acquire_bits_payload_client_xact_id;
  wire[511:0] net_io_masters_0_acquire_bits_payload_data;
  wire net_io_masters_0_acquire_bits_payload_uncached;
  wire[1:0] net_io_masters_0_acquire_bits_payload_a_type;
  wire[511:0] net_io_masters_0_acquire_bits_payload_subblock;
  wire net_io_masters_0_grant_ready;
  wire net_io_masters_0_finish_valid;
  wire[1:0] net_io_masters_0_finish_bits_header_src;
  wire[1:0] net_io_masters_0_finish_bits_header_dst;
  wire[2:0] net_io_masters_0_finish_bits_payload_master_xact_id;
  wire net_io_masters_0_probe_ready;
  wire net_io_masters_0_release_valid;
  wire[1:0] net_io_masters_0_release_bits_header_src;
  wire[1:0] net_io_masters_0_release_bits_header_dst;
  wire[25:0] net_io_masters_0_release_bits_payload_addr;
  wire[2:0] net_io_masters_0_release_bits_payload_client_xact_id;
  wire[511:0] net_io_masters_0_release_bits_payload_data;
  wire[2:0] net_io_masters_0_release_bits_payload_r_type;
  wire L2CoherenceAgent_io_inner_acquire_ready;
  wire L2CoherenceAgent_io_inner_grant_valid;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_dst;
  wire[511:0] L2CoherenceAgent_io_inner_grant_bits_payload_data;
  wire[2:0] L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id;
  wire L2CoherenceAgent_io_inner_grant_bits_payload_uncached;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_payload_g_type;
  wire L2CoherenceAgent_io_inner_finish_ready;
  wire L2CoherenceAgent_io_inner_probe_valid;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_dst;
  wire[25:0] L2CoherenceAgent_io_inner_probe_bits_payload_addr;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_payload_p_type;
  wire L2CoherenceAgent_io_inner_release_ready;
  wire L2CoherenceAgent_io_outer_acquire_valid;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_dst;
  wire[25:0] L2CoherenceAgent_io_outer_acquire_bits_payload_addr;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] L2CoherenceAgent_io_outer_acquire_bits_payload_data;
  wire L2CoherenceAgent_io_outer_acquire_bits_payload_uncached;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_payload_a_type;
  wire[511:0] L2CoherenceAgent_io_outer_acquire_bits_payload_subblock;
  wire L2CoherenceAgent_io_outer_grant_ready;
  wire L2CoherenceAgent_io_outer_finish_valid;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_dst;
  wire L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id;
  wire conv_io_uncached_acquire_ready;
  wire conv_io_uncached_grant_valid;
  wire[511:0] conv_io_uncached_grant_bits_payload_data;
  wire[2:0] conv_io_uncached_grant_bits_payload_client_xact_id;
  wire conv_io_uncached_grant_bits_payload_master_xact_id;
  wire conv_io_uncached_grant_bits_payload_uncached;
  wire[1:0] conv_io_uncached_grant_bits_payload_g_type;
  wire conv_io_mem_req_cmd_valid;
  wire[25:0] conv_io_mem_req_cmd_bits_addr;
  wire[4:0] conv_io_mem_req_cmd_bits_tag;
  wire conv_io_mem_req_cmd_bits_rw;
  wire conv_io_mem_req_data_valid;
  wire[127:0] conv_io_mem_req_data_bits_data;


  assign io_mem_req_data_bits_data = conv_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = conv_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = conv_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = conv_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = conv_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = conv_io_mem_req_cmd_valid;
  assign io_htif_release_ready = net_io_clients_1_release_ready;
  assign io_htif_probe_bits_payload_p_type = net_io_clients_1_probe_bits_payload_p_type;
  assign io_htif_probe_bits_payload_addr = net_io_clients_1_probe_bits_payload_addr;
  assign io_htif_probe_bits_header_dst = net_io_clients_1_probe_bits_header_dst;
  assign io_htif_probe_bits_header_src = net_io_clients_1_probe_bits_header_src;
  assign io_htif_probe_valid = net_io_clients_1_probe_valid;
  assign io_htif_finish_ready = net_io_clients_1_finish_ready;
  assign io_htif_grant_bits_payload_g_type = net_io_clients_1_grant_bits_payload_g_type;
  assign io_htif_grant_bits_payload_uncached = net_io_clients_1_grant_bits_payload_uncached;
  assign io_htif_grant_bits_payload_master_xact_id = net_io_clients_1_grant_bits_payload_master_xact_id;
  assign io_htif_grant_bits_payload_client_xact_id = net_io_clients_1_grant_bits_payload_client_xact_id;
  assign io_htif_grant_bits_payload_data = net_io_clients_1_grant_bits_payload_data;
  assign io_htif_grant_bits_header_dst = net_io_clients_1_grant_bits_header_dst;
  assign io_htif_grant_bits_header_src = net_io_clients_1_grant_bits_header_src;
  assign io_htif_grant_valid = net_io_clients_1_grant_valid;
  assign io_htif_acquire_ready = net_io_clients_1_acquire_ready;
  assign io_tiles_0_release_ready = net_io_clients_0_release_ready;
  assign io_tiles_0_probe_bits_payload_p_type = net_io_clients_0_probe_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_addr = net_io_clients_0_probe_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = net_io_clients_0_probe_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = net_io_clients_0_probe_bits_header_src;
  assign io_tiles_0_probe_valid = net_io_clients_0_probe_valid;
  assign io_tiles_0_finish_ready = net_io_clients_0_finish_ready;
  assign io_tiles_0_grant_bits_payload_g_type = net_io_clients_0_grant_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_uncached = net_io_clients_0_grant_bits_payload_uncached;
  assign io_tiles_0_grant_bits_payload_master_xact_id = net_io_clients_0_grant_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = net_io_clients_0_grant_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = net_io_clients_0_grant_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = net_io_clients_0_grant_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = net_io_clients_0_grant_bits_header_src;
  assign io_tiles_0_grant_valid = net_io_clients_0_grant_valid;
  assign io_tiles_0_acquire_ready = net_io_clients_0_acquire_ready;
  RocketChipCrossbarNetwork net(.clk(clk), .reset(reset),
       .io_clients_1_acquire_ready( net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( io_htif_acquire_valid ),
       .io_clients_1_acquire_bits_header_src( io_htif_acquire_bits_header_src ),
       .io_clients_1_acquire_bits_header_dst( io_htif_acquire_bits_header_dst ),
       .io_clients_1_acquire_bits_payload_addr( io_htif_acquire_bits_payload_addr ),
       .io_clients_1_acquire_bits_payload_client_xact_id( io_htif_acquire_bits_payload_client_xact_id ),
       .io_clients_1_acquire_bits_payload_data( io_htif_acquire_bits_payload_data ),
       .io_clients_1_acquire_bits_payload_uncached( io_htif_acquire_bits_payload_uncached ),
       .io_clients_1_acquire_bits_payload_a_type( io_htif_acquire_bits_payload_a_type ),
       .io_clients_1_acquire_bits_payload_subblock( io_htif_acquire_bits_payload_subblock ),
       .io_clients_1_grant_ready( io_htif_grant_ready ),
       .io_clients_1_grant_valid( net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_header_src( net_io_clients_1_grant_bits_header_src ),
       .io_clients_1_grant_bits_header_dst( net_io_clients_1_grant_bits_header_dst ),
       .io_clients_1_grant_bits_payload_data( net_io_clients_1_grant_bits_payload_data ),
       .io_clients_1_grant_bits_payload_client_xact_id( net_io_clients_1_grant_bits_payload_client_xact_id ),
       .io_clients_1_grant_bits_payload_master_xact_id( net_io_clients_1_grant_bits_payload_master_xact_id ),
       .io_clients_1_grant_bits_payload_uncached( net_io_clients_1_grant_bits_payload_uncached ),
       .io_clients_1_grant_bits_payload_g_type( net_io_clients_1_grant_bits_payload_g_type ),
       .io_clients_1_finish_ready( net_io_clients_1_finish_ready ),
       .io_clients_1_finish_valid( io_htif_finish_valid ),
       .io_clients_1_finish_bits_header_src( io_htif_finish_bits_header_src ),
       .io_clients_1_finish_bits_header_dst( io_htif_finish_bits_header_dst ),
       .io_clients_1_finish_bits_payload_master_xact_id( io_htif_finish_bits_payload_master_xact_id ),
       .io_clients_1_probe_ready( io_htif_probe_ready ),
       .io_clients_1_probe_valid( net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_header_src( net_io_clients_1_probe_bits_header_src ),
       .io_clients_1_probe_bits_header_dst( net_io_clients_1_probe_bits_header_dst ),
       .io_clients_1_probe_bits_payload_addr( net_io_clients_1_probe_bits_payload_addr ),
       .io_clients_1_probe_bits_payload_p_type( net_io_clients_1_probe_bits_payload_p_type ),
       .io_clients_1_release_ready( net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( io_htif_release_valid ),
       .io_clients_1_release_bits_header_src( io_htif_release_bits_header_src ),
       .io_clients_1_release_bits_header_dst( io_htif_release_bits_header_dst ),
       .io_clients_1_release_bits_payload_addr( io_htif_release_bits_payload_addr ),
       .io_clients_1_release_bits_payload_client_xact_id( io_htif_release_bits_payload_client_xact_id ),
       .io_clients_1_release_bits_payload_data( io_htif_release_bits_payload_data ),
       .io_clients_1_release_bits_payload_r_type( io_htif_release_bits_payload_r_type ),
       .io_clients_0_acquire_ready( net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_0_acquire_valid ),
       .io_clients_0_acquire_bits_header_src( io_tiles_0_acquire_bits_header_src ),
       .io_clients_0_acquire_bits_header_dst( io_tiles_0_acquire_bits_header_dst ),
       .io_clients_0_acquire_bits_payload_addr( io_tiles_0_acquire_bits_payload_addr ),
       .io_clients_0_acquire_bits_payload_client_xact_id( io_tiles_0_acquire_bits_payload_client_xact_id ),
       .io_clients_0_acquire_bits_payload_data( io_tiles_0_acquire_bits_payload_data ),
       .io_clients_0_acquire_bits_payload_uncached( io_tiles_0_acquire_bits_payload_uncached ),
       .io_clients_0_acquire_bits_payload_a_type( io_tiles_0_acquire_bits_payload_a_type ),
       .io_clients_0_acquire_bits_payload_subblock( io_tiles_0_acquire_bits_payload_subblock ),
       .io_clients_0_grant_ready( io_tiles_0_grant_ready ),
       .io_clients_0_grant_valid( net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_header_src( net_io_clients_0_grant_bits_header_src ),
       .io_clients_0_grant_bits_header_dst( net_io_clients_0_grant_bits_header_dst ),
       .io_clients_0_grant_bits_payload_data( net_io_clients_0_grant_bits_payload_data ),
       .io_clients_0_grant_bits_payload_client_xact_id( net_io_clients_0_grant_bits_payload_client_xact_id ),
       .io_clients_0_grant_bits_payload_master_xact_id( net_io_clients_0_grant_bits_payload_master_xact_id ),
       .io_clients_0_grant_bits_payload_uncached( net_io_clients_0_grant_bits_payload_uncached ),
       .io_clients_0_grant_bits_payload_g_type( net_io_clients_0_grant_bits_payload_g_type ),
       .io_clients_0_finish_ready( net_io_clients_0_finish_ready ),
       .io_clients_0_finish_valid( io_tiles_0_finish_valid ),
       .io_clients_0_finish_bits_header_src( io_tiles_0_finish_bits_header_src ),
       .io_clients_0_finish_bits_header_dst( io_tiles_0_finish_bits_header_dst ),
       .io_clients_0_finish_bits_payload_master_xact_id( io_tiles_0_finish_bits_payload_master_xact_id ),
       .io_clients_0_probe_ready( io_tiles_0_probe_ready ),
       .io_clients_0_probe_valid( net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_header_src( net_io_clients_0_probe_bits_header_src ),
       .io_clients_0_probe_bits_header_dst( net_io_clients_0_probe_bits_header_dst ),
       .io_clients_0_probe_bits_payload_addr( net_io_clients_0_probe_bits_payload_addr ),
       .io_clients_0_probe_bits_payload_p_type( net_io_clients_0_probe_bits_payload_p_type ),
       .io_clients_0_release_ready( net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_0_release_valid ),
       .io_clients_0_release_bits_header_src( io_tiles_0_release_bits_header_src ),
       .io_clients_0_release_bits_header_dst( io_tiles_0_release_bits_header_dst ),
       .io_clients_0_release_bits_payload_addr( io_tiles_0_release_bits_payload_addr ),
       .io_clients_0_release_bits_payload_client_xact_id( io_tiles_0_release_bits_payload_client_xact_id ),
       .io_clients_0_release_bits_payload_data( io_tiles_0_release_bits_payload_data ),
       .io_clients_0_release_bits_payload_r_type( io_tiles_0_release_bits_payload_r_type ),
       .io_masters_0_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_masters_0_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_masters_0_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_masters_0_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_masters_0_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_masters_0_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_masters_0_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_masters_0_acquire_bits_payload_uncached( net_io_masters_0_acquire_bits_payload_uncached ),
       .io_masters_0_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_masters_0_acquire_bits_payload_subblock( net_io_masters_0_acquire_bits_payload_subblock ),
       .io_masters_0_grant_ready( net_io_masters_0_grant_ready ),
       .io_masters_0_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_masters_0_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_masters_0_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_masters_0_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_masters_0_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_masters_0_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_masters_0_grant_bits_payload_uncached( L2CoherenceAgent_io_inner_grant_bits_payload_uncached ),
       .io_masters_0_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_masters_0_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_masters_0_finish_valid( net_io_masters_0_finish_valid ),
       .io_masters_0_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_masters_0_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_masters_0_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_masters_0_probe_ready( net_io_masters_0_probe_ready ),
       .io_masters_0_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_masters_0_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_masters_0_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_masters_0_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_masters_0_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_masters_0_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_masters_0_release_valid( net_io_masters_0_release_valid ),
       .io_masters_0_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_masters_0_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_masters_0_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_masters_0_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_masters_0_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_masters_0_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type )
  );
  L2CoherenceAgent L2CoherenceAgent(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_inner_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_inner_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_uncached( net_io_masters_0_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( net_io_masters_0_acquire_bits_payload_subblock ),
       .io_inner_grant_ready( net_io_masters_0_grant_ready ),
       .io_inner_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_uncached( L2CoherenceAgent_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_inner_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_inner_finish_valid( net_io_masters_0_finish_valid ),
       .io_inner_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( net_io_masters_0_probe_ready ),
       .io_inner_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_inner_release_valid( net_io_masters_0_release_valid ),
       .io_inner_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_inner_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type ),
       .io_outer_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_outer_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_outer_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_outer_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( L2CoherenceAgent_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( L2CoherenceAgent_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_outer_grant_valid( conv_io_uncached_grant_valid ),
       //.io_outer_grant_bits_header_src(  )
       //.io_outer_grant_bits_header_dst(  )
       .io_outer_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_uncached( conv_io_uncached_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_outer_finish_ready(  )
       .io_outer_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_outer_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_outer_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_outer_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_incoherent_1( io_incoherent_1 ),
       .io_incoherent_0( io_incoherent_0 )
  );
  `ifndef SYNTHESIS
    assign L2CoherenceAgent.io_outer_grant_bits_header_src = {1{$random}};
    assign L2CoherenceAgent.io_outer_grant_bits_header_dst = {1{$random}};
    assign L2CoherenceAgent.io_outer_finish_ready = {1{$random}};
  `endif
  MemPipeIOUncachedTileLinkIOConverter conv(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_uncached_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_uncached( L2CoherenceAgent_io_outer_acquire_bits_payload_uncached ),
       .io_uncached_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_subblock( L2CoherenceAgent_io_outer_acquire_bits_payload_subblock ),
       .io_uncached_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_uncached_grant_valid( conv_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_uncached( conv_io_uncached_grant_bits_payload_uncached ),
       .io_uncached_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_uncached_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( conv_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( conv_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( conv_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [2:0] io_enq_bits_payload_client_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input  io_enq_bits_payload_uncached,
    input [1:0] io_enq_bits_payload_a_type,
    input [511:0] io_enq_bits_payload_subblock,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[2:0] io_deq_bits_payload_client_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output io_deq_bits_payload_uncached,
    output[1:0] io_deq_bits_payload_a_type,
    output[511:0] io_deq_bits_payload_subblock
);

  wire[511:0] T0;
  wire[1059:0] T1;
  reg [1059:0] ram [1:0];
  wire[1059:0] T2;
  wire[1059:0] T3;
  wire[1059:0] T4;
  wire[1026:0] T5;
  wire[513:0] T6;
  wire[512:0] T7;
  wire[32:0] T8;
  wire[28:0] T9;
  wire[3:0] T10;
  wire do_enq;
  reg  R11;
  wire T29;
  wire T12;
  wire T13;
  reg  R14;
  wire T30;
  wire T15;
  wire T16;
  wire do_deq;
  wire[1:0] T17;
  wire T18;
  wire[511:0] T19;
  wire[2:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire empty;
  wire T25;
  reg  maybe_full;
  wire T31;
  wire T26;
  wire T27;
  wire ptr_match;
  wire T28;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {34{$random}};
    R11 = {1{$random}};
    R14 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_subblock = T0;
  assign T0 = T1[9'h1ff:1'h0];
  assign T1 = ram[R14];
  assign T3 = T4;
  assign T4 = {T8, T5};
  assign T5 = {T7, T6};
  assign T6 = {io_enq_bits_payload_a_type, io_enq_bits_payload_subblock};
  assign T7 = {io_enq_bits_payload_data, io_enq_bits_payload_uncached};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T10 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T29 = reset ? 1'h0 : T12;
  assign T12 = do_enq ? T13 : R11;
  assign T13 = R11 + 1'h1;
  assign T30 = reset ? 1'h0 : T15;
  assign T15 = do_deq ? T16 : R14;
  assign T16 = R14 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_a_type = T17;
  assign T17 = T1[10'h201:10'h200];
  assign io_deq_bits_payload_uncached = T18;
  assign T18 = T1[10'h202:10'h202];
  assign io_deq_bits_payload_data = T19;
  assign T19 = T1[11'h402:10'h203];
  assign io_deq_bits_payload_client_xact_id = T20;
  assign T20 = T1[11'h405:11'h403];
  assign io_deq_bits_payload_addr = T21;
  assign T21 = T1[11'h41f:11'h406];
  assign io_deq_bits_header_dst = T22;
  assign T22 = T1[11'h421:11'h420];
  assign io_deq_bits_header_src = T23;
  assign T23 = T1[11'h423:11'h422];
  assign io_deq_valid = T24;
  assign T24 = empty ^ 1'h1;
  assign empty = ptr_match & T25;
  assign T25 = maybe_full ^ 1'h1;
  assign T31 = reset ? 1'h0 : T26;
  assign T26 = T27 ? do_enq : maybe_full;
  assign T27 = do_enq != do_deq;
  assign ptr_match = R11 == R14;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R11] <= T3;
    if(reset) begin
      R11 <= 1'h0;
    end else if(do_enq) begin
      R11 <= T13;
    end
    if(reset) begin
      R14 <= 1'h0;
    end else if(do_deq) begin
      R14 <= T16;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T27) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [2:0] io_enq_bits_payload_client_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[2:0] io_deq_bits_payload_client_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type
);

  wire[2:0] T0;
  wire[547:0] T1;
  reg [547:0] ram [1:0];
  wire[547:0] T2;
  wire[547:0] T3;
  wire[547:0] T4;
  wire[517:0] T5;
  wire[514:0] T6;
  wire[29:0] T7;
  wire[27:0] T8;
  wire do_enq;
  reg  R9;
  wire T25;
  wire T10;
  wire T11;
  reg  R12;
  wire T26;
  wire T13;
  wire T14;
  wire do_deq;
  wire[511:0] T15;
  wire[2:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire empty;
  wire T21;
  reg  maybe_full;
  wire T27;
  wire T22;
  wire T23;
  wire ptr_match;
  wire T24;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R9 = {1{$random}};
    R12 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_r_type = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R12];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_client_xact_id, T6};
  assign T6 = {io_enq_bits_payload_data, io_enq_bits_payload_r_type};
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_addr};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T25 = reset ? 1'h0 : T10;
  assign T10 = do_enq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign T26 = reset ? 1'h0 : T13;
  assign T13 = do_deq ? T14 : R12;
  assign T14 = R12 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T15;
  assign T15 = T1[10'h202:2'h3];
  assign io_deq_bits_payload_client_xact_id = T16;
  assign T16 = T1[10'h205:10'h203];
  assign io_deq_bits_payload_addr = T17;
  assign T17 = T1[10'h21f:10'h206];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T1[10'h221:10'h220];
  assign io_deq_bits_header_src = T19;
  assign T19 = T1[10'h223:10'h222];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign T27 = reset ? 1'h0 : T22;
  assign T22 = T23 ? do_enq : maybe_full;
  assign T23 = do_enq != do_deq;
  assign ptr_match = R9 == R12;
  assign io_enq_ready = T24;
  assign T24 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R9] <= T3;
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_enq) begin
      R9 <= T11;
    end
    if(reset) begin
      R12 <= 1'h0;
    end else if(do_deq) begin
      R12 <= T14;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T23) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id
);

  wire[2:0] T0;
  wire[6:0] T1;
  reg [6:0] ram [1:0];
  wire[6:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire[4:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_master_xact_id = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_header_src, T5};
  assign T5 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_header_dst = T12;
  assign T12 = T1[3'h4:2'h3];
  assign io_deq_bits_header_src = T13;
  assign T13 = T1[3'h6:3'h5];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_enq_bits_payload_uncached,
    input [1:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output io_deq_bits_payload_uncached,
    output[1:0] io_deq_bits_payload_g_type
);

  wire[1:0] T0;
  wire[524:0] T1;
  reg [524:0] ram [0:0];
  wire[524:0] T2;
  wire[524:0] T3;
  wire[524:0] T4;
  wire[8:0] T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[515:0] T8;
  wire[513:0] T9;
  wire do_enq;
  wire T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[511:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire empty;
  reg  full;
  wire T21;
  wire T17;
  wire T18;
  wire do_deq;
  wire T19;
  wire T20;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {17{$random}};
    full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_g_type = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {T8, T5};
  assign T5 = {T7, T6};
  assign T6 = {io_enq_bits_payload_uncached, io_enq_bits_payload_g_type};
  assign T7 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_master_xact_id};
  assign T8 = {io_enq_bits_header_src, T9};
  assign T9 = {io_enq_bits_header_dst, io_enq_bits_payload_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_payload_uncached = T10;
  assign T10 = T1[2'h2:2'h2];
  assign io_deq_bits_payload_master_xact_id = T11;
  assign T11 = T1[3'h5:2'h3];
  assign io_deq_bits_payload_client_xact_id = T12;
  assign T12 = T1[4'h8:3'h6];
  assign io_deq_bits_payload_data = T13;
  assign T13 = T1[10'h208:4'h9];
  assign io_deq_bits_header_dst = T14;
  assign T14 = T1[10'h20a:10'h209];
  assign io_deq_bits_header_src = T15;
  assign T15 = T1[10'h20c:10'h20b];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T17;
  assign T17 = T18 ? do_enq : full;
  assign T18 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T19;
  assign T19 = T20 | io_deq_ready;
  assign T20 = full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      full <= 1'h0;
    end else if(T18) begin
      full <= do_enq;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_p_type
);

  wire[1:0] T0;
  wire[31:0] T1;
  reg [31:0] ram [1:0];
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[27:0] T5;
  wire[3:0] T6;
  wire do_enq;
  reg  R7;
  wire T21;
  wire T8;
  wire T9;
  reg  R10;
  wire T22;
  wire T11;
  wire T12;
  wire do_deq;
  wire[25:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire empty;
  wire T17;
  reg  maybe_full;
  wire T23;
  wire T18;
  wire T19;
  wire ptr_match;
  wire T20;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R7 = {1{$random}};
    R10 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_p_type = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = ram[R10];
  assign T3 = T4;
  assign T4 = {T6, T5};
  assign T5 = {io_enq_bits_payload_addr, io_enq_bits_payload_p_type};
  assign T6 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = do_enq ? T9 : R7;
  assign T9 = R7 + 1'h1;
  assign T22 = reset ? 1'h0 : T11;
  assign T11 = do_deq ? T12 : R10;
  assign T12 = R10 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_addr = T13;
  assign T13 = T1[5'h1b:2'h2];
  assign io_deq_bits_header_dst = T14;
  assign T14 = T1[5'h1d:5'h1c];
  assign io_deq_bits_header_src = T15;
  assign T15 = T1[5'h1f:5'h1e];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign T23 = reset ? 1'h0 : T18;
  assign T18 = T19 ? do_enq : maybe_full;
  assign T19 = do_enq != do_deq;
  assign ptr_match = R7 == R10;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R7] <= T3;
    if(reset) begin
      R7 <= 1'h0;
    end else if(do_enq) begin
      R7 <= T9;
    end
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_deq) begin
      R10 <= T12;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T19) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [2:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input  io_tiles_0_acquire_bits_payload_uncached,
    input [1:0] io_tiles_0_acquire_bits_payload_a_type,
    input [511:0] io_tiles_0_acquire_bits_payload_subblock,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[2:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output io_tiles_0_grant_bits_payload_uncached,
    output[1:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [2:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[4:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr,
    input  io_incoherent_0
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire[2:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[511:0] T8;
  wire[2:0] T9;
  wire[25:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[511:0] T14;
  wire[1:0] T15;
  wire T16;
  wire[511:0] T17;
  wire[2:0] T18;
  wire[25:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[2:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire[2:0] T27;
  wire[511:0] T28;
  wire[2:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire[511:0] T34;
  wire[1:0] T35;
  wire T36;
  wire[511:0] T37;
  wire[2:0] T38;
  wire[25:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T0;
  wire T1;
  wire T2;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[25:0] Queue_4_io_deq_bits_payload_addr;
  wire[2:0] Queue_4_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_4_io_deq_bits_payload_data;
  wire Queue_4_io_deq_bits_payload_uncached;
  wire[1:0] Queue_4_io_deq_bits_payload_a_type;
  wire[511:0] Queue_4_io_deq_bits_payload_subblock;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[1:0] Queue_5_io_deq_bits_header_src;
  wire[1:0] Queue_5_io_deq_bits_header_dst;
  wire[25:0] Queue_5_io_deq_bits_payload_addr;
  wire[2:0] Queue_5_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_5_io_deq_bits_payload_data;
  wire[2:0] Queue_5_io_deq_bits_payload_r_type;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[1:0] Queue_6_io_deq_bits_header_src;
  wire[1:0] Queue_6_io_deq_bits_header_dst;
  wire[2:0] Queue_6_io_deq_bits_payload_master_xact_id;
  wire Queue_7_io_enq_ready;
  wire Queue_7_io_deq_valid;
  wire[1:0] Queue_7_io_deq_bits_header_src;
  wire[1:0] Queue_7_io_deq_bits_header_dst;
  wire[511:0] Queue_7_io_deq_bits_payload_data;
  wire[2:0] Queue_7_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_7_io_deq_bits_payload_master_xact_id;
  wire Queue_7_io_deq_bits_payload_uncached;
  wire[1:0] Queue_7_io_deq_bits_payload_g_type;
  wire Queue_8_io_enq_ready;
  wire Queue_8_io_deq_valid;
  wire[1:0] Queue_8_io_deq_bits_header_src;
  wire[1:0] Queue_8_io_deq_bits_header_dst;
  wire[25:0] Queue_8_io_deq_bits_payload_addr;
  wire[1:0] Queue_8_io_deq_bits_payload_p_type;
  wire Queue_9_io_enq_ready;
  wire Queue_9_io_deq_valid;
  wire[1:0] Queue_9_io_deq_bits_header_src;
  wire[1:0] Queue_9_io_deq_bits_header_dst;
  wire[25:0] Queue_9_io_deq_bits_payload_addr;
  wire[2:0] Queue_9_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_9_io_deq_bits_payload_data;
  wire Queue_9_io_deq_bits_payload_uncached;
  wire[1:0] Queue_9_io_deq_bits_payload_a_type;
  wire[511:0] Queue_9_io_deq_bits_payload_subblock;
  wire Queue_10_io_enq_ready;
  wire Queue_10_io_deq_valid;
  wire[1:0] Queue_10_io_deq_bits_header_src;
  wire[1:0] Queue_10_io_deq_bits_header_dst;
  wire[25:0] Queue_10_io_deq_bits_payload_addr;
  wire[2:0] Queue_10_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_10_io_deq_bits_payload_data;
  wire[2:0] Queue_10_io_deq_bits_payload_r_type;
  wire Queue_11_io_enq_ready;
  wire Queue_11_io_deq_valid;
  wire[1:0] Queue_11_io_deq_bits_header_src;
  wire[1:0] Queue_11_io_deq_bits_header_dst;
  wire[2:0] Queue_11_io_deq_bits_payload_master_xact_id;
  wire Queue_12_io_enq_ready;
  wire Queue_12_io_deq_valid;
  wire[1:0] Queue_12_io_deq_bits_header_src;
  wire[1:0] Queue_12_io_deq_bits_header_dst;
  wire[511:0] Queue_12_io_deq_bits_payload_data;
  wire[2:0] Queue_12_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_12_io_deq_bits_payload_master_xact_id;
  wire Queue_12_io_deq_bits_payload_uncached;
  wire[1:0] Queue_12_io_deq_bits_payload_g_type;
  wire Queue_13_io_enq_ready;
  wire Queue_13_io_deq_valid;
  wire[1:0] Queue_13_io_deq_bits_header_src;
  wire[1:0] Queue_13_io_deq_bits_header_dst;
  wire[25:0] Queue_13_io_deq_bits_payload_addr;
  wire[1:0] Queue_13_io_deq_bits_payload_p_type;
  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_pcr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire[4:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_payload_addr;
  wire[2:0] htif_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] htif_io_mem_acquire_bits_payload_data;
  wire htif_io_mem_acquire_bits_payload_uncached;
  wire[1:0] htif_io_mem_acquire_bits_payload_a_type;
  wire[511:0] htif_io_mem_acquire_bits_payload_subblock;
  wire htif_io_mem_grant_ready;
  wire htif_io_mem_finish_valid;
  wire[1:0] htif_io_mem_finish_bits_header_dst;
  wire[2:0] htif_io_mem_finish_bits_payload_master_xact_id;
  wire htif_io_mem_probe_ready;
  wire htif_io_mem_release_valid;
  wire[25:0] htif_io_mem_release_bits_payload_addr;
  wire[2:0] htif_io_mem_release_bits_payload_client_xact_id;
  wire[511:0] htif_io_mem_release_bits_payload_data;
  wire[2:0] htif_io_mem_release_bits_payload_r_type;
  wire outmemsys_io_tiles_0_acquire_ready;
  wire outmemsys_io_tiles_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_dst;
  wire[511:0] outmemsys_io_tiles_0_grant_bits_payload_data;
  wire[2:0] outmemsys_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[2:0] outmemsys_io_tiles_0_grant_bits_payload_master_xact_id;
  wire outmemsys_io_tiles_0_grant_bits_payload_uncached;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_payload_g_type;
  wire outmemsys_io_tiles_0_finish_ready;
  wire outmemsys_io_tiles_0_probe_valid;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_dst;
  wire[25:0] outmemsys_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_payload_p_type;
  wire outmemsys_io_tiles_0_release_ready;
  wire outmemsys_io_htif_acquire_ready;
  wire outmemsys_io_htif_grant_valid;
  wire[1:0] outmemsys_io_htif_grant_bits_header_src;
  wire[1:0] outmemsys_io_htif_grant_bits_header_dst;
  wire[511:0] outmemsys_io_htif_grant_bits_payload_data;
  wire[2:0] outmemsys_io_htif_grant_bits_payload_client_xact_id;
  wire[2:0] outmemsys_io_htif_grant_bits_payload_master_xact_id;
  wire outmemsys_io_htif_grant_bits_payload_uncached;
  wire[1:0] outmemsys_io_htif_grant_bits_payload_g_type;
  wire outmemsys_io_htif_finish_ready;
  wire outmemsys_io_htif_probe_valid;
  wire[1:0] outmemsys_io_htif_probe_bits_header_src;
  wire[1:0] outmemsys_io_htif_probe_bits_header_dst;
  wire[25:0] outmemsys_io_htif_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_htif_probe_bits_payload_p_type;
  wire outmemsys_io_htif_release_ready;
  wire outmemsys_io_mem_req_cmd_valid;
  wire[25:0] outmemsys_io_mem_req_cmd_bits_addr;
  wire[4:0] outmemsys_io_mem_req_cmd_bits_tag;
  wire outmemsys_io_mem_req_cmd_bits_rw;
  wire outmemsys_io_mem_req_data_valid;
  wire[127:0] outmemsys_io_mem_req_data_bits_data;


  assign T3 = htif_io_mem_finish_bits_payload_master_xact_id;
  assign T4 = htif_io_mem_finish_bits_header_dst;
  assign T5 = 2'h1;
  assign T6 = htif_io_mem_finish_valid;
  assign T7 = htif_io_mem_release_bits_payload_r_type;
  assign T8 = htif_io_mem_release_bits_payload_data;
  assign T9 = htif_io_mem_release_bits_payload_client_xact_id;
  assign T10 = htif_io_mem_release_bits_payload_addr;
  assign T11 = 2'h0;
  assign T12 = 2'h1;
  assign T13 = htif_io_mem_release_valid;
  assign T14 = htif_io_mem_acquire_bits_payload_subblock;
  assign T15 = htif_io_mem_acquire_bits_payload_a_type;
  assign T16 = htif_io_mem_acquire_bits_payload_uncached;
  assign T17 = htif_io_mem_acquire_bits_payload_data;
  assign T18 = htif_io_mem_acquire_bits_payload_client_xact_id;
  assign T19 = htif_io_mem_acquire_bits_payload_addr;
  assign T20 = 2'h0;
  assign T21 = 2'h1;
  assign T22 = htif_io_mem_acquire_valid;
  assign T23 = io_tiles_0_finish_bits_payload_master_xact_id;
  assign T24 = io_tiles_0_finish_bits_header_dst;
  assign T25 = 2'h0;
  assign T26 = io_tiles_0_finish_valid;
  assign T27 = io_tiles_0_release_bits_payload_r_type;
  assign T28 = io_tiles_0_release_bits_payload_data;
  assign T29 = io_tiles_0_release_bits_payload_client_xact_id;
  assign T30 = io_tiles_0_release_bits_payload_addr;
  assign T31 = 2'h0;
  assign T32 = 2'h0;
  assign T33 = io_tiles_0_release_valid;
  assign T34 = io_tiles_0_acquire_bits_payload_subblock;
  assign T35 = io_tiles_0_acquire_bits_payload_a_type;
  assign T36 = io_tiles_0_acquire_bits_payload_uncached;
  assign T37 = io_tiles_0_acquire_bits_payload_data;
  assign T38 = io_tiles_0_acquire_bits_payload_client_xact_id;
  assign T39 = io_tiles_0_acquire_bits_payload_addr;
  assign T40 = 2'h0;
  assign T41 = 2'h0;
  assign T42 = io_tiles_0_acquire_valid;
  assign T43 = Queue_10_io_enq_ready;
  assign T44 = Queue_11_io_enq_ready;
  assign T45 = Queue_9_io_enq_ready;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_tiles_0_release_ready = T0;
  assign T0 = Queue_5_io_enq_ready;
  assign io_tiles_0_probe_bits_payload_p_type = Queue_8_io_deq_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_addr = Queue_8_io_deq_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = Queue_8_io_deq_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = Queue_8_io_deq_bits_header_src;
  assign io_tiles_0_probe_valid = Queue_8_io_deq_valid;
  assign io_tiles_0_finish_ready = T1;
  assign T1 = Queue_6_io_enq_ready;
  assign io_tiles_0_grant_bits_payload_g_type = Queue_7_io_deq_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_uncached = Queue_7_io_deq_bits_payload_uncached;
  assign io_tiles_0_grant_bits_payload_master_xact_id = Queue_7_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = Queue_7_io_deq_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = Queue_7_io_deq_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = Queue_7_io_deq_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = Queue_7_io_deq_bits_header_src;
  assign io_tiles_0_grant_valid = Queue_7_io_deq_valid;
  assign io_tiles_0_acquire_ready = T2;
  assign T2 = Queue_4_io_enq_ready;
  assign io_mem_req_data_bits_data = outmemsys_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = outmemsys_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = outmemsys_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = outmemsys_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = outmemsys_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = outmemsys_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = htif_io_host_debug_stats_pcr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_pcr( htif_io_host_debug_stats_pcr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( T45 ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( htif_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( htif_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( htif_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( htif_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( htif_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( htif_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( Queue_12_io_deq_valid ),
       .io_mem_grant_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_mem_grant_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_mem_grant_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( Queue_12_io_deq_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_uncached( Queue_12_io_deq_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type ),
       .io_mem_finish_ready( T44 ),
       .io_mem_finish_valid( htif_io_mem_finish_valid ),
       //.io_mem_finish_bits_header_src(  )
       .io_mem_finish_bits_header_dst( htif_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( htif_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( htif_io_mem_probe_ready ),
       .io_mem_probe_valid( Queue_13_io_deq_valid ),
       .io_mem_probe_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_mem_probe_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_mem_probe_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type ),
       .io_mem_release_ready( T43 ),
       .io_mem_release_valid( htif_io_mem_release_valid ),
       //.io_mem_release_bits_header_src(  )
       //.io_mem_release_bits_header_dst(  )
       .io_mem_release_bits_payload_addr( htif_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( htif_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_data( htif_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( htif_io_mem_release_bits_payload_r_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
  `ifndef SYNTHESIS
    assign htif.io_mem_release_bits_payload_addr = {1{$random}};
    assign htif.io_mem_release_bits_payload_client_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_data = {16{$random}};
    assign htif.io_mem_release_bits_payload_r_type = {1{$random}};
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
  `endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_0_acquire_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Queue_4_io_deq_valid ),
       .io_tiles_0_acquire_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_uncached( Queue_4_io_deq_bits_payload_uncached ),
       .io_tiles_0_acquire_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_subblock( Queue_4_io_deq_bits_payload_subblock ),
       .io_tiles_0_grant_ready( Queue_7_io_enq_ready ),
       .io_tiles_0_grant_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_uncached( outmemsys_io_tiles_0_grant_bits_payload_uncached ),
       .io_tiles_0_grant_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Queue_6_io_deq_valid ),
       .io_tiles_0_finish_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Queue_8_io_enq_ready ),
       .io_tiles_0_probe_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( outmemsys_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Queue_5_io_deq_valid ),
       .io_tiles_0_release_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type ),
       .io_htif_acquire_ready( outmemsys_io_htif_acquire_ready ),
       .io_htif_acquire_valid( Queue_9_io_deq_valid ),
       .io_htif_acquire_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_htif_acquire_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_htif_acquire_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_htif_acquire_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_htif_acquire_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_htif_acquire_bits_payload_uncached( Queue_9_io_deq_bits_payload_uncached ),
       .io_htif_acquire_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_htif_acquire_bits_payload_subblock( Queue_9_io_deq_bits_payload_subblock ),
       .io_htif_grant_ready( Queue_12_io_enq_ready ),
       .io_htif_grant_valid( outmemsys_io_htif_grant_valid ),
       .io_htif_grant_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_htif_grant_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_htif_grant_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_htif_grant_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_htif_grant_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_htif_grant_bits_payload_uncached( outmemsys_io_htif_grant_bits_payload_uncached ),
       .io_htif_grant_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_htif_finish_ready( outmemsys_io_htif_finish_ready ),
       .io_htif_finish_valid( Queue_11_io_deq_valid ),
       .io_htif_finish_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_htif_finish_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_htif_finish_bits_payload_master_xact_id( Queue_11_io_deq_bits_payload_master_xact_id ),
       .io_htif_probe_ready( Queue_13_io_enq_ready ),
       .io_htif_probe_valid( outmemsys_io_htif_probe_valid ),
       .io_htif_probe_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_htif_probe_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_htif_probe_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_htif_probe_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_htif_release_ready( outmemsys_io_htif_release_ready ),
       .io_htif_release_valid( Queue_10_io_deq_valid ),
       .io_htif_release_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_htif_release_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_htif_release_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_htif_release_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_htif_release_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_htif_release_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type ),
       .io_incoherent_1( 1'h1 ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( outmemsys_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( outmemsys_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( outmemsys_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( outmemsys_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( outmemsys_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( outmemsys_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( T42 ),
       .io_enq_bits_header_src( T41 ),
       .io_enq_bits_header_dst( T40 ),
       .io_enq_bits_payload_addr( T39 ),
       .io_enq_bits_payload_client_xact_id( T38 ),
       .io_enq_bits_payload_data( T37 ),
       .io_enq_bits_payload_uncached( T36 ),
       .io_enq_bits_payload_a_type( T35 ),
       .io_enq_bits_payload_subblock( T34 ),
       .io_deq_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_deq_bits_payload_uncached( Queue_4_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_subblock( Queue_4_io_deq_bits_payload_subblock )
  );
  Queue_4 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( T33 ),
       .io_enq_bits_header_src( T32 ),
       .io_enq_bits_header_dst( T31 ),
       .io_enq_bits_payload_addr( T30 ),
       .io_enq_bits_payload_client_xact_id( T29 ),
       .io_enq_bits_payload_data( T28 ),
       .io_enq_bits_payload_r_type( T27 ),
       .io_deq_ready( outmemsys_io_tiles_0_release_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type )
  );
  Queue_5 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( T26 ),
       .io_enq_bits_header_src( T25 ),
       .io_enq_bits_header_dst( T24 ),
       .io_enq_bits_payload_master_xact_id( T23 ),
       .io_deq_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id )
  );
  Queue_6 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_uncached( outmemsys_io_tiles_0_grant_bits_payload_uncached ),
       .io_enq_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_deq_ready( io_tiles_0_grant_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_7_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_7_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_uncached( Queue_7_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_g_type( Queue_7_io_deq_bits_payload_g_type )
  );
  Queue_7 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_enq_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_deq_ready( io_tiles_0_probe_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_8_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_p_type( Queue_8_io_deq_bits_payload_p_type )
  );
  Queue_3 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( T22 ),
       .io_enq_bits_header_src( T21 ),
       .io_enq_bits_header_dst( T20 ),
       .io_enq_bits_payload_addr( T19 ),
       .io_enq_bits_payload_client_xact_id( T18 ),
       .io_enq_bits_payload_data( T17 ),
       .io_enq_bits_payload_uncached( T16 ),
       .io_enq_bits_payload_a_type( T15 ),
       .io_enq_bits_payload_subblock( T14 ),
       .io_deq_ready( outmemsys_io_htif_acquire_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_deq_bits_payload_uncached( Queue_9_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_subblock( Queue_9_io_deq_bits_payload_subblock )
  );
  Queue_4 Queue_10(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_10_io_enq_ready ),
       .io_enq_valid( T13 ),
       .io_enq_bits_header_src( T12 ),
       .io_enq_bits_header_dst( T11 ),
       .io_enq_bits_payload_addr( T10 ),
       .io_enq_bits_payload_client_xact_id( T9 ),
       .io_enq_bits_payload_data( T8 ),
       .io_enq_bits_payload_r_type( T7 ),
       .io_deq_ready( outmemsys_io_htif_release_ready ),
       .io_deq_valid( Queue_10_io_deq_valid ),
       .io_deq_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type )
  );
  Queue_5 Queue_11(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_11_io_enq_ready ),
       .io_enq_valid( T6 ),
       .io_enq_bits_header_src( T5 ),
       .io_enq_bits_header_dst( T4 ),
       .io_enq_bits_payload_master_xact_id( T3 ),
       .io_deq_ready( outmemsys_io_htif_finish_ready ),
       .io_deq_valid( Queue_11_io_deq_valid ),
       .io_deq_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_11_io_deq_bits_payload_master_xact_id )
  );
  Queue_6 Queue_12(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_12_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_uncached( outmemsys_io_htif_grant_bits_payload_uncached ),
       .io_enq_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_deq_ready( htif_io_mem_grant_ready ),
       .io_deq_valid( Queue_12_io_deq_valid ),
       .io_deq_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_12_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_uncached( Queue_12_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type )
  );
  Queue_7 Queue_13(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_13_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_enq_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_deq_ready( htif_io_mem_probe_ready ),
       .io_deq_valid( Queue_13_io_deq_valid ),
       .io_deq_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type )
  );
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [4:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[4:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data
);

  wire[63:0] T0;
  wire[69:0] T1;
  reg [69:0] ram [1:0];
  wire[69:0] T2;
  wire[69:0] T3;
  wire[69:0] T4;
  wire[68:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[4:0] T12;
  wire T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_rw, T5};
  assign T5 = {io_enq_bits_addr, io_enq_bits_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_addr = T12;
  assign T12 = T1[7'h44:7'h40];
  assign io_deq_bits_rw = T13;
  assign T13 = T1[7'h45:7'h45];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits
);

  wire[63:0] T0;
  reg [63:0] ram [1:0];
  wire[63:0] T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits
);

  wire T0;
  reg [0:0] ram [1:0];
  wire T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module PearsonHasher(input clk, input reset,
    input  io_keyData_valid,
    input [7:0] io_keyData_bits,
    input [5:0] io_keyLen,
    output[7:0] io_romAddr_1,
    output[7:0] io_romAddr_0,
    input [7:0] io_romData_1,
    input [7:0] io_romData_0,
    output io_result_valid,
    output[15:0] io_result_bits,
    input  io_restart
);

  wire[15:0] T0;
  reg [7:0] h_0;
  wire[7:0] T1;
  wire[7:0] T2;
  wire T3;
  wire T4;
  wire T5;
  reg [5:0] index;
  wire[5:0] T21;
  wire[5:0] T6;
  wire[5:0] T7;
  wire[5:0] T8;
  wire T9;
  reg [7:0] h_1;
  wire[7:0] T10;
  wire[7:0] T11;
  wire T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[7:0] T15;
  wire T16;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire T20;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    h_0 = {1{$random}};
    index = {1{$random}};
    h_1 = {1{$random}};
  end
`endif

  assign io_result_bits = T0;
  assign T0 = {h_1, h_0};
  assign T1 = T3 ? io_romData_0 : T2;
  assign T2 = io_restart ? 8'h0 : h_0;
  assign T3 = T9 & T4;
  assign T4 = T5 & io_keyData_valid;
  assign T5 = index != io_keyLen;
  assign T21 = reset ? 6'h0 : T6;
  assign T6 = T3 ? T8 : T7;
  assign T7 = io_restart ? 6'h0 : index;
  assign T8 = index + 6'h1;
  assign T9 = io_restart ^ 1'h1;
  assign T10 = T3 ? io_romData_1 : T11;
  assign T11 = io_restart ? 8'h0 : h_1;
  assign io_result_valid = T12;
  assign T12 = index == io_keyLen;
  assign io_romAddr_0 = T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = h_0 ^ io_keyData_bits;
  assign T15 = io_keyData_bits + 8'h0;
  assign T16 = index == 6'h0;
  assign io_romAddr_1 = T17;
  assign T17 = T20 ? T19 : T18;
  assign T18 = h_1 ^ io_keyData_bits;
  assign T19 = io_keyData_bits + 8'h1;
  assign T20 = index == 6'h0;

  always @(posedge clk) begin
    if(T3) begin
      h_0 <= io_romData_0;
    end else if(io_restart) begin
      h_0 <= 8'h0;
    end
    if(reset) begin
      index <= 6'h0;
    end else if(T3) begin
      index <= T8;
    end else if(io_restart) begin
      index <= 6'h0;
    end
    if(T3) begin
      h_1 <= io_romData_1;
    end else if(io_restart) begin
      h_1 <= 8'h0;
    end
  end
endmodule

module HasherWriter(input clk, input reset,
    output[5:0] io_keyWriteAddr,
    output[31:0] io_keyWriteData,
    output io_keyWrite,
    output io_keyData_ready,
    input  io_keyData_valid,
    input [7:0] io_keyData_bits,
    output io_keyInfo_ready,
    input  io_keyInfo_valid,
    input [7:0] io_keyInfo_bits_len,
    input [3:0] io_keyInfo_bits_tag,
    input  io_hashOut_ready,
    output io_hashOut_valid,
    output[9:0] io_hashOut_bits_hash1,
    output[9:0] io_hashOut_bits_hash2,
    output[7:0] io_hashOut_bits_len,
    output[3:0] io_hashOut_bits_tag,
    input  io_lock,
    output io_halted
);

  reg  restart;
  wire T57;
  wire T58;
  wire T59;
  wire T8;
  reg [1:0] state;
  wire[1:0] T46;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T9;
  wire T10;
  wire[7:0] T11;
  reg [7:0] keyLen;
  wire[7:0] T12;
  reg [7:0] index;
  wire[7:0] T47;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[7:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [7:0] T60;
  reg [7:0] T61;
  wire[5:0] T62;
  wire hashInputValid;
  wire T63;
  reg [7:0] T64;
  reg [7:0] T65;
  wire[5:0] T66;
  wire T0;
  wire T1;
  reg [3:0] keyTag;
  wire[3:0] T20;
  wire[9:0] T48;
  wire[9:0] T49;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  reg  keyWrite;
  wire T50;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] byteOff;
  wire T33;
  reg [31:0] keyWriteData;
  wire[31:0] T51;
  wire[38:0] T52;
  wire[38:0] T34;
  wire[38:0] T53;
  wire[31:0] T35;
  wire[31:0] T54;
  wire T36;
  wire T37;
  wire[38:0] T38;
  wire[38:0] T39;
  wire[4:0] inputShift;
  wire[38:0] T55;
  wire T40;
  wire T41;
  reg [5:0] keyWriteAddr;
  wire[5:0] T56;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[7:0] PearsonHasher_0_io_romAddr_1;
  wire[7:0] PearsonHasher_0_io_romAddr_0;
  wire[15:0] PearsonHasher_0_io_result_bits;
  wire[7:0] PearsonHasher_1_io_romAddr_1;
  wire[7:0] PearsonHasher_1_io_romAddr_0;
  wire[15:0] PearsonHasher_1_io_result_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    restart = {1{$random}};
    state = {1{$random}};
    keyLen = {1{$random}};
    index = {1{$random}};
    keyTag = {1{$random}};
    keyWrite = {1{$random}};
    keyWriteData = {1{$random}};
    keyWriteAddr = {1{$random}};
  end
`endif

  assign T57 = reset ? 1'h0 : T58;
  assign T58 = T18 ? 1'h1 : T59;
  assign T59 = T8 ? 1'h0 : restart;
  assign T8 = 2'h0 == state;
  assign T46 = reset ? 2'h0 : T2;
  assign T2 = T18 ? 2'h0 : T3;
  assign T3 = T9 ? 2'h2 : T4;
  assign T4 = T5 ? 2'h1 : state;
  assign T5 = T8 & T6;
  assign T6 = io_keyInfo_valid & T7;
  assign T7 = io_lock ^ 1'h1;
  assign T9 = T16 & T10;
  assign T10 = index == T11;
  assign T11 = keyLen - 8'h1;
  assign T12 = T5 ? io_keyInfo_bits_len : keyLen;
  assign T47 = reset ? 8'h0 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = T5 ? 8'h0 : index;
  assign T15 = index + 8'h1;
  assign T16 = T17 & io_keyData_valid;
  assign T17 = 2'h1 == state;
  assign T18 = T19 & io_hashOut_ready;
  assign T19 = 2'h2 == state;
  always @(*) case (PearsonHasher_1_io_romAddr_0)
    0: T60 = 8'h17;
    1: T60 = 8'h7d;
    2: T60 = 8'h39;
    3: T60 = 8'h10;
    4: T60 = 8'h6;
    5: T60 = 8'h16;
    6: T60 = 8'hae;
    7: T60 = 8'haf;
    8: T60 = 8'h7b;
    9: T60 = 8'hc9;
    10: T60 = 8'hce;
    11: T60 = 8'he8;
    12: T60 = 8'h77;
    13: T60 = 8'hcf;
    14: T60 = 8'h29;
    15: T60 = 8'h89;
    16: T60 = 8'hb6;
    17: T60 = 8'h64;
    18: T60 = 8'h3c;
    19: T60 = 8'hf6;
    20: T60 = 8'h3b;
    21: T60 = 8'h0;
    22: T60 = 8'h84;
    23: T60 = 8'hda;
    24: T60 = 8'hc1;
    25: T60 = 8'h3e;
    26: T60 = 8'h75;
    27: T60 = 8'ha0;
    28: T60 = 8'he6;
    29: T60 = 8'h25;
    30: T60 = 8'h4b;
    31: T60 = 8'hb0;
    32: T60 = 8'h6b;
    33: T60 = 8'hf7;
    34: T60 = 8'h79;
    35: T60 = 8'h1f;
    36: T60 = 8'hb2;
    37: T60 = 8'h5;
    38: T60 = 8'hc7;
    39: T60 = 8'h47;
    40: T60 = 8'h55;
    41: T60 = 8'h72;
    42: T60 = 8'ha6;
    43: T60 = 8'h68;
    44: T60 = 8'hd5;
    45: T60 = 8'hac;
    46: T60 = 8'h8e;
    47: T60 = 8'h9e;
    48: T60 = 8'h18;
    49: T60 = 8'h82;
    50: T60 = 8'h96;
    51: T60 = 8'h8;
    52: T60 = 8'h93;
    53: T60 = 8'hd6;
    54: T60 = 8'h50;
    55: T60 = 8'he0;
    56: T60 = 8'h2e;
    57: T60 = 8'h9;
    58: T60 = 8'h53;
    59: T60 = 8'h7;
    60: T60 = 8'hb4;
    61: T60 = 8'had;
    62: T60 = 8'h22;
    63: T60 = 8'h66;
    64: T60 = 8'hb1;
    65: T60 = 8'h1a;
    66: T60 = 8'he5;
    67: T60 = 8'hbe;
    68: T60 = 8'h38;
    69: T60 = 8'h4e;
    70: T60 = 8'he;
    71: T60 = 8'h86;
    72: T60 = 8'h8a;
    73: T60 = 8'hb5;
    74: T60 = 8'h5a;
    75: T60 = 8'hde;
    76: T60 = 8'h9c;
    77: T60 = 8'h58;
    78: T60 = 8'hfa;
    79: T60 = 8'h7c;
    80: T60 = 8'h28;
    81: T60 = 8'h6f;
    82: T60 = 8'h51;
    83: T60 = 8'h1d;
    84: T60 = 8'he4;
    85: T60 = 8'h11;
    86: T60 = 8'h65;
    87: T60 = 8'h30;
    88: T60 = 8'hb;
    89: T60 = 8'h52;
    90: T60 = 8'h4c;
    91: T60 = 8'h4f;
    92: T60 = 8'h73;
    93: T60 = 8'h5f;
    94: T60 = 8'hb3;
    95: T60 = 8'hdc;
    96: T60 = 8'h95;
    97: T60 = 8'h3;
    98: T60 = 8'h87;
    99: T60 = 8'h56;
    100: T60 = 8'hc0;
    101: T60 = 8'hdf;
    102: T60 = 8'h14;
    103: T60 = 8'h91;
    104: T60 = 8'h19;
    105: T60 = 8'h7f;
    106: T60 = 8'hd7;
    107: T60 = 8'hc6;
    108: T60 = 8'hf8;
    109: T60 = 8'hea;
    110: T60 = 8'h61;
    111: T60 = 8'h85;
    112: T60 = 8'h97;
    113: T60 = 8'hd8;
    114: T60 = 8'h8b;
    115: T60 = 8'he9;
    116: T60 = 8'hd0;
    117: T60 = 8'hd2;
    118: T60 = 8'h2a;
    119: T60 = 8'h43;
    120: T60 = 8'h31;
    121: T60 = 8'hfc;
    122: T60 = 8'hd;
    123: T60 = 8'h6a;
    124: T60 = 8'ha5;
    125: T60 = 8'hf2;
    126: T60 = 8'hf4;
    127: T60 = 8'h12;
    128: T60 = 8'hbd;
    129: T60 = 8'h35;
    130: T60 = 8'h90;
    131: T60 = 8'hed;
    132: T60 = 8'heb;
    133: T60 = 8'haa;
    134: T60 = 8'h32;
    135: T60 = 8'h7e;
    136: T60 = 8'h76;
    137: T60 = 8'h37;
    138: T60 = 8'h24;
    139: T60 = 8'h9d;
    140: T60 = 8'h9f;
    141: T60 = 8'hb7;
    142: T60 = 8'h5e;
    143: T60 = 8'h5d;
    144: T60 = 8'hec;
    145: T60 = 8'h3a;
    146: T60 = 8'h69;
    147: T60 = 8'h49;
    148: T60 = 8'h94;
    149: T60 = 8'h57;
    150: T60 = 8'h8c;
    151: T60 = 8'h62;
    152: T60 = 8'hc8;
    153: T60 = 8'h23;
    154: T60 = 8'h70;
    155: T60 = 8'hc4;
    156: T60 = 8'h59;
    157: T60 = 8'h2b;
    158: T60 = 8'h81;
    159: T60 = 8'h5b;
    160: T60 = 8'hf5;
    161: T60 = 8'h13;
    162: T60 = 8'h20;
    163: T60 = 8'h34;
    164: T60 = 8'hba;
    165: T60 = 8'h80;
    166: T60 = 8'h46;
    167: T60 = 8'hf3;
    168: T60 = 8'h6d;
    169: T60 = 8'hbb;
    170: T60 = 8'hf1;
    171: T60 = 8'h1;
    172: T60 = 8'hee;
    173: T60 = 8'h2;
    174: T60 = 8'hfd;
    175: T60 = 8'hb9;
    176: T60 = 8'hb8;
    177: T60 = 8'hbf;
    178: T60 = 8'he3;
    179: T60 = 8'h44;
    180: T60 = 8'h83;
    181: T60 = 8'h1c;
    182: T60 = 8'h45;
    183: T60 = 8'hd1;
    184: T60 = 8'ha2;
    185: T60 = 8'ha;
    186: T60 = 8'he1;
    187: T60 = 8'hfe;
    188: T60 = 8'ha1;
    189: T60 = 8'h54;
    190: T60 = 8'h63;
    191: T60 = 8'hc2;
    192: T60 = 8'h2f;
    193: T60 = 8'h15;
    194: T60 = 8'hcc;
    195: T60 = 8'h36;
    196: T60 = 8'h33;
    197: T60 = 8'he2;
    198: T60 = 8'ha3;
    199: T60 = 8'h74;
    200: T60 = 8'h99;
    201: T60 = 8'h8d;
    202: T60 = 8'hd3;
    203: T60 = 8'hbc;
    204: T60 = 8'hca;
    205: T60 = 8'hd4;
    206: T60 = 8'ha9;
    207: T60 = 8'h1e;
    208: T60 = 8'h67;
    209: T60 = 8'h6c;
    210: T60 = 8'h9b;
    211: T60 = 8'hff;
    212: T60 = 8'h21;
    213: T60 = 8'h5c;
    214: T60 = 8'hc3;
    215: T60 = 8'hc;
    216: T60 = 8'h40;
    217: T60 = 8'h78;
    218: T60 = 8'h3d;
    219: T60 = 8'hf0;
    220: T60 = 8'h3f;
    221: T60 = 8'hfb;
    222: T60 = 8'h27;
    223: T60 = 8'h41;
    224: T60 = 8'h92;
    225: T60 = 8'h71;
    226: T60 = 8'h4d;
    227: T60 = 8'h8f;
    228: T60 = 8'h4;
    229: T60 = 8'hc5;
    230: T60 = 8'hf;
    231: T60 = 8'h2d;
    232: T60 = 8'h7a;
    233: T60 = 8'he7;
    234: T60 = 8'h26;
    235: T60 = 8'h2c;
    236: T60 = 8'h88;
    237: T60 = 8'hd9;
    238: T60 = 8'ha7;
    239: T60 = 8'hcd;
    240: T60 = 8'h98;
    241: T60 = 8'hcb;
    242: T60 = 8'h42;
    243: T60 = 8'hf9;
    244: T60 = 8'h1b;
    245: T60 = 8'hab;
    246: T60 = 8'ha4;
    247: T60 = 8'h48;
    248: T60 = 8'hdb;
    249: T60 = 8'hdd;
    250: T60 = 8'h6e;
    251: T60 = 8'ha8;
    252: T60 = 8'h4a;
    253: T60 = 8'hef;
    254: T60 = 8'h9a;
    255: T60 = 8'h60;
`ifndef SYNTHESIS
    default: T60 = {1{$random}};
`else
    default: T60 = 8'bx;
`endif
  endcase
  always @(*) case (PearsonHasher_1_io_romAddr_1)
    0: T61 = 8'h17;
    1: T61 = 8'h7d;
    2: T61 = 8'h39;
    3: T61 = 8'h10;
    4: T61 = 8'h6;
    5: T61 = 8'h16;
    6: T61 = 8'hae;
    7: T61 = 8'haf;
    8: T61 = 8'h7b;
    9: T61 = 8'hc9;
    10: T61 = 8'hce;
    11: T61 = 8'he8;
    12: T61 = 8'h77;
    13: T61 = 8'hcf;
    14: T61 = 8'h29;
    15: T61 = 8'h89;
    16: T61 = 8'hb6;
    17: T61 = 8'h64;
    18: T61 = 8'h3c;
    19: T61 = 8'hf6;
    20: T61 = 8'h3b;
    21: T61 = 8'h0;
    22: T61 = 8'h84;
    23: T61 = 8'hda;
    24: T61 = 8'hc1;
    25: T61 = 8'h3e;
    26: T61 = 8'h75;
    27: T61 = 8'ha0;
    28: T61 = 8'he6;
    29: T61 = 8'h25;
    30: T61 = 8'h4b;
    31: T61 = 8'hb0;
    32: T61 = 8'h6b;
    33: T61 = 8'hf7;
    34: T61 = 8'h79;
    35: T61 = 8'h1f;
    36: T61 = 8'hb2;
    37: T61 = 8'h5;
    38: T61 = 8'hc7;
    39: T61 = 8'h47;
    40: T61 = 8'h55;
    41: T61 = 8'h72;
    42: T61 = 8'ha6;
    43: T61 = 8'h68;
    44: T61 = 8'hd5;
    45: T61 = 8'hac;
    46: T61 = 8'h8e;
    47: T61 = 8'h9e;
    48: T61 = 8'h18;
    49: T61 = 8'h82;
    50: T61 = 8'h96;
    51: T61 = 8'h8;
    52: T61 = 8'h93;
    53: T61 = 8'hd6;
    54: T61 = 8'h50;
    55: T61 = 8'he0;
    56: T61 = 8'h2e;
    57: T61 = 8'h9;
    58: T61 = 8'h53;
    59: T61 = 8'h7;
    60: T61 = 8'hb4;
    61: T61 = 8'had;
    62: T61 = 8'h22;
    63: T61 = 8'h66;
    64: T61 = 8'hb1;
    65: T61 = 8'h1a;
    66: T61 = 8'he5;
    67: T61 = 8'hbe;
    68: T61 = 8'h38;
    69: T61 = 8'h4e;
    70: T61 = 8'he;
    71: T61 = 8'h86;
    72: T61 = 8'h8a;
    73: T61 = 8'hb5;
    74: T61 = 8'h5a;
    75: T61 = 8'hde;
    76: T61 = 8'h9c;
    77: T61 = 8'h58;
    78: T61 = 8'hfa;
    79: T61 = 8'h7c;
    80: T61 = 8'h28;
    81: T61 = 8'h6f;
    82: T61 = 8'h51;
    83: T61 = 8'h1d;
    84: T61 = 8'he4;
    85: T61 = 8'h11;
    86: T61 = 8'h65;
    87: T61 = 8'h30;
    88: T61 = 8'hb;
    89: T61 = 8'h52;
    90: T61 = 8'h4c;
    91: T61 = 8'h4f;
    92: T61 = 8'h73;
    93: T61 = 8'h5f;
    94: T61 = 8'hb3;
    95: T61 = 8'hdc;
    96: T61 = 8'h95;
    97: T61 = 8'h3;
    98: T61 = 8'h87;
    99: T61 = 8'h56;
    100: T61 = 8'hc0;
    101: T61 = 8'hdf;
    102: T61 = 8'h14;
    103: T61 = 8'h91;
    104: T61 = 8'h19;
    105: T61 = 8'h7f;
    106: T61 = 8'hd7;
    107: T61 = 8'hc6;
    108: T61 = 8'hf8;
    109: T61 = 8'hea;
    110: T61 = 8'h61;
    111: T61 = 8'h85;
    112: T61 = 8'h97;
    113: T61 = 8'hd8;
    114: T61 = 8'h8b;
    115: T61 = 8'he9;
    116: T61 = 8'hd0;
    117: T61 = 8'hd2;
    118: T61 = 8'h2a;
    119: T61 = 8'h43;
    120: T61 = 8'h31;
    121: T61 = 8'hfc;
    122: T61 = 8'hd;
    123: T61 = 8'h6a;
    124: T61 = 8'ha5;
    125: T61 = 8'hf2;
    126: T61 = 8'hf4;
    127: T61 = 8'h12;
    128: T61 = 8'hbd;
    129: T61 = 8'h35;
    130: T61 = 8'h90;
    131: T61 = 8'hed;
    132: T61 = 8'heb;
    133: T61 = 8'haa;
    134: T61 = 8'h32;
    135: T61 = 8'h7e;
    136: T61 = 8'h76;
    137: T61 = 8'h37;
    138: T61 = 8'h24;
    139: T61 = 8'h9d;
    140: T61 = 8'h9f;
    141: T61 = 8'hb7;
    142: T61 = 8'h5e;
    143: T61 = 8'h5d;
    144: T61 = 8'hec;
    145: T61 = 8'h3a;
    146: T61 = 8'h69;
    147: T61 = 8'h49;
    148: T61 = 8'h94;
    149: T61 = 8'h57;
    150: T61 = 8'h8c;
    151: T61 = 8'h62;
    152: T61 = 8'hc8;
    153: T61 = 8'h23;
    154: T61 = 8'h70;
    155: T61 = 8'hc4;
    156: T61 = 8'h59;
    157: T61 = 8'h2b;
    158: T61 = 8'h81;
    159: T61 = 8'h5b;
    160: T61 = 8'hf5;
    161: T61 = 8'h13;
    162: T61 = 8'h20;
    163: T61 = 8'h34;
    164: T61 = 8'hba;
    165: T61 = 8'h80;
    166: T61 = 8'h46;
    167: T61 = 8'hf3;
    168: T61 = 8'h6d;
    169: T61 = 8'hbb;
    170: T61 = 8'hf1;
    171: T61 = 8'h1;
    172: T61 = 8'hee;
    173: T61 = 8'h2;
    174: T61 = 8'hfd;
    175: T61 = 8'hb9;
    176: T61 = 8'hb8;
    177: T61 = 8'hbf;
    178: T61 = 8'he3;
    179: T61 = 8'h44;
    180: T61 = 8'h83;
    181: T61 = 8'h1c;
    182: T61 = 8'h45;
    183: T61 = 8'hd1;
    184: T61 = 8'ha2;
    185: T61 = 8'ha;
    186: T61 = 8'he1;
    187: T61 = 8'hfe;
    188: T61 = 8'ha1;
    189: T61 = 8'h54;
    190: T61 = 8'h63;
    191: T61 = 8'hc2;
    192: T61 = 8'h2f;
    193: T61 = 8'h15;
    194: T61 = 8'hcc;
    195: T61 = 8'h36;
    196: T61 = 8'h33;
    197: T61 = 8'he2;
    198: T61 = 8'ha3;
    199: T61 = 8'h74;
    200: T61 = 8'h99;
    201: T61 = 8'h8d;
    202: T61 = 8'hd3;
    203: T61 = 8'hbc;
    204: T61 = 8'hca;
    205: T61 = 8'hd4;
    206: T61 = 8'ha9;
    207: T61 = 8'h1e;
    208: T61 = 8'h67;
    209: T61 = 8'h6c;
    210: T61 = 8'h9b;
    211: T61 = 8'hff;
    212: T61 = 8'h21;
    213: T61 = 8'h5c;
    214: T61 = 8'hc3;
    215: T61 = 8'hc;
    216: T61 = 8'h40;
    217: T61 = 8'h78;
    218: T61 = 8'h3d;
    219: T61 = 8'hf0;
    220: T61 = 8'h3f;
    221: T61 = 8'hfb;
    222: T61 = 8'h27;
    223: T61 = 8'h41;
    224: T61 = 8'h92;
    225: T61 = 8'h71;
    226: T61 = 8'h4d;
    227: T61 = 8'h8f;
    228: T61 = 8'h4;
    229: T61 = 8'hc5;
    230: T61 = 8'hf;
    231: T61 = 8'h2d;
    232: T61 = 8'h7a;
    233: T61 = 8'he7;
    234: T61 = 8'h26;
    235: T61 = 8'h2c;
    236: T61 = 8'h88;
    237: T61 = 8'hd9;
    238: T61 = 8'ha7;
    239: T61 = 8'hcd;
    240: T61 = 8'h98;
    241: T61 = 8'hcb;
    242: T61 = 8'h42;
    243: T61 = 8'hf9;
    244: T61 = 8'h1b;
    245: T61 = 8'hab;
    246: T61 = 8'ha4;
    247: T61 = 8'h48;
    248: T61 = 8'hdb;
    249: T61 = 8'hdd;
    250: T61 = 8'h6e;
    251: T61 = 8'ha8;
    252: T61 = 8'h4a;
    253: T61 = 8'hef;
    254: T61 = 8'h9a;
    255: T61 = 8'h60;
`ifndef SYNTHESIS
    default: T61 = {1{$random}};
`else
    default: T61 = 8'bx;
`endif
  endcase
  assign T62 = keyLen[3'h5:1'h0];
  assign hashInputValid = io_keyData_valid & T63;
  assign T63 = state == 2'h1;
  always @(*) case (PearsonHasher_0_io_romAddr_0)
    0: T64 = 8'h62;
    1: T64 = 8'h6;
    2: T64 = 8'h55;
    3: T64 = 8'h96;
    4: T64 = 8'h24;
    5: T64 = 8'h17;
    6: T64 = 8'h70;
    7: T64 = 8'ha4;
    8: T64 = 8'h87;
    9: T64 = 8'hcf;
    10: T64 = 8'ha9;
    11: T64 = 8'h5;
    12: T64 = 8'h1a;
    13: T64 = 8'h40;
    14: T64 = 8'ha5;
    15: T64 = 8'hdb;
    16: T64 = 8'h3d;
    17: T64 = 8'h14;
    18: T64 = 8'h44;
    19: T64 = 8'h59;
    20: T64 = 8'h82;
    21: T64 = 8'h3f;
    22: T64 = 8'h34;
    23: T64 = 8'h66;
    24: T64 = 8'h18;
    25: T64 = 8'he5;
    26: T64 = 8'h84;
    27: T64 = 8'hf5;
    28: T64 = 8'h50;
    29: T64 = 8'hd8;
    30: T64 = 8'hc3;
    31: T64 = 8'h73;
    32: T64 = 8'h5a;
    33: T64 = 8'ha8;
    34: T64 = 8'h9c;
    35: T64 = 8'hcb;
    36: T64 = 8'hb1;
    37: T64 = 8'h78;
    38: T64 = 8'h2;
    39: T64 = 8'hbe;
    40: T64 = 8'hbc;
    41: T64 = 8'h7;
    42: T64 = 8'h64;
    43: T64 = 8'hb9;
    44: T64 = 8'hae;
    45: T64 = 8'hf3;
    46: T64 = 8'ha2;
    47: T64 = 8'ha;
    48: T64 = 8'hed;
    49: T64 = 8'h12;
    50: T64 = 8'hfd;
    51: T64 = 8'he1;
    52: T64 = 8'h8;
    53: T64 = 8'hd0;
    54: T64 = 8'hac;
    55: T64 = 8'hf4;
    56: T64 = 8'hff;
    57: T64 = 8'h7e;
    58: T64 = 8'h65;
    59: T64 = 8'h4f;
    60: T64 = 8'h91;
    61: T64 = 8'heb;
    62: T64 = 8'he4;
    63: T64 = 8'h79;
    64: T64 = 8'h7b;
    65: T64 = 8'hfb;
    66: T64 = 8'h43;
    67: T64 = 8'hfa;
    68: T64 = 8'ha1;
    69: T64 = 8'h0;
    70: T64 = 8'h6b;
    71: T64 = 8'h61;
    72: T64 = 8'hf1;
    73: T64 = 8'h6f;
    74: T64 = 8'hb5;
    75: T64 = 8'h52;
    76: T64 = 8'hf9;
    77: T64 = 8'h21;
    78: T64 = 8'h45;
    79: T64 = 8'h37;
    80: T64 = 8'h3b;
    81: T64 = 8'h99;
    82: T64 = 8'h1d;
    83: T64 = 8'h9;
    84: T64 = 8'hd5;
    85: T64 = 8'ha7;
    86: T64 = 8'h54;
    87: T64 = 8'h5d;
    88: T64 = 8'h1e;
    89: T64 = 8'h2e;
    90: T64 = 8'h5e;
    91: T64 = 8'h4b;
    92: T64 = 8'h97;
    93: T64 = 8'h72;
    94: T64 = 8'h49;
    95: T64 = 8'hde;
    96: T64 = 8'hc5;
    97: T64 = 8'h60;
    98: T64 = 8'hd2;
    99: T64 = 8'h2d;
    100: T64 = 8'h10;
    101: T64 = 8'he3;
    102: T64 = 8'hf8;
    103: T64 = 8'hca;
    104: T64 = 8'h33;
    105: T64 = 8'h98;
    106: T64 = 8'hfc;
    107: T64 = 8'h7d;
    108: T64 = 8'h51;
    109: T64 = 8'hce;
    110: T64 = 8'hd7;
    111: T64 = 8'hba;
    112: T64 = 8'h27;
    113: T64 = 8'h9e;
    114: T64 = 8'hb2;
    115: T64 = 8'hbb;
    116: T64 = 8'h83;
    117: T64 = 8'h88;
    118: T64 = 8'h1;
    119: T64 = 8'h31;
    120: T64 = 8'h32;
    121: T64 = 8'h11;
    122: T64 = 8'h8d;
    123: T64 = 8'h5b;
    124: T64 = 8'h2f;
    125: T64 = 8'h81;
    126: T64 = 8'h3c;
    127: T64 = 8'h63;
    128: T64 = 8'h9a;
    129: T64 = 8'h23;
    130: T64 = 8'h56;
    131: T64 = 8'hab;
    132: T64 = 8'h69;
    133: T64 = 8'h22;
    134: T64 = 8'h26;
    135: T64 = 8'hc8;
    136: T64 = 8'h93;
    137: T64 = 8'h3a;
    138: T64 = 8'h4d;
    139: T64 = 8'h76;
    140: T64 = 8'had;
    141: T64 = 8'hf6;
    142: T64 = 8'h4c;
    143: T64 = 8'hfe;
    144: T64 = 8'h85;
    145: T64 = 8'he8;
    146: T64 = 8'hc4;
    147: T64 = 8'h90;
    148: T64 = 8'hc6;
    149: T64 = 8'h7c;
    150: T64 = 8'h35;
    151: T64 = 8'h4;
    152: T64 = 8'h6c;
    153: T64 = 8'h4a;
    154: T64 = 8'hdf;
    155: T64 = 8'hea;
    156: T64 = 8'h86;
    157: T64 = 8'he6;
    158: T64 = 8'h9d;
    159: T64 = 8'h8b;
    160: T64 = 8'hbd;
    161: T64 = 8'hcd;
    162: T64 = 8'hc7;
    163: T64 = 8'h80;
    164: T64 = 8'hb0;
    165: T64 = 8'h13;
    166: T64 = 8'hd3;
    167: T64 = 8'hec;
    168: T64 = 8'h7f;
    169: T64 = 8'hc0;
    170: T64 = 8'he7;
    171: T64 = 8'h46;
    172: T64 = 8'he9;
    173: T64 = 8'h58;
    174: T64 = 8'h92;
    175: T64 = 8'h2c;
    176: T64 = 8'hb7;
    177: T64 = 8'hc9;
    178: T64 = 8'h16;
    179: T64 = 8'h53;
    180: T64 = 8'hd;
    181: T64 = 8'hd6;
    182: T64 = 8'h74;
    183: T64 = 8'h6d;
    184: T64 = 8'h9f;
    185: T64 = 8'h20;
    186: T64 = 8'h5f;
    187: T64 = 8'he2;
    188: T64 = 8'h8c;
    189: T64 = 8'hdc;
    190: T64 = 8'h39;
    191: T64 = 8'hc;
    192: T64 = 8'hdd;
    193: T64 = 8'h1f;
    194: T64 = 8'hd1;
    195: T64 = 8'hb6;
    196: T64 = 8'h8f;
    197: T64 = 8'h5c;
    198: T64 = 8'h95;
    199: T64 = 8'hb8;
    200: T64 = 8'h94;
    201: T64 = 8'h3e;
    202: T64 = 8'h71;
    203: T64 = 8'h41;
    204: T64 = 8'h25;
    205: T64 = 8'h1b;
    206: T64 = 8'h6a;
    207: T64 = 8'ha6;
    208: T64 = 8'h3;
    209: T64 = 8'he;
    210: T64 = 8'hcc;
    211: T64 = 8'h48;
    212: T64 = 8'h15;
    213: T64 = 8'h29;
    214: T64 = 8'h38;
    215: T64 = 8'h42;
    216: T64 = 8'h1c;
    217: T64 = 8'hc1;
    218: T64 = 8'h28;
    219: T64 = 8'hd9;
    220: T64 = 8'h19;
    221: T64 = 8'h36;
    222: T64 = 8'hb3;
    223: T64 = 8'h75;
    224: T64 = 8'hee;
    225: T64 = 8'h57;
    226: T64 = 8'hf0;
    227: T64 = 8'h9b;
    228: T64 = 8'hb4;
    229: T64 = 8'haa;
    230: T64 = 8'hf2;
    231: T64 = 8'hd4;
    232: T64 = 8'hbf;
    233: T64 = 8'ha3;
    234: T64 = 8'h4e;
    235: T64 = 8'hda;
    236: T64 = 8'h89;
    237: T64 = 8'hc2;
    238: T64 = 8'haf;
    239: T64 = 8'h6e;
    240: T64 = 8'h2b;
    241: T64 = 8'h77;
    242: T64 = 8'he0;
    243: T64 = 8'h47;
    244: T64 = 8'h7a;
    245: T64 = 8'h8e;
    246: T64 = 8'h2a;
    247: T64 = 8'ha0;
    248: T64 = 8'h68;
    249: T64 = 8'h30;
    250: T64 = 8'hf7;
    251: T64 = 8'h67;
    252: T64 = 8'hf;
    253: T64 = 8'hb;
    254: T64 = 8'h8a;
    255: T64 = 8'hef;
`ifndef SYNTHESIS
    default: T64 = {1{$random}};
`else
    default: T64 = 8'bx;
`endif
  endcase
  always @(*) case (PearsonHasher_0_io_romAddr_1)
    0: T65 = 8'h62;
    1: T65 = 8'h6;
    2: T65 = 8'h55;
    3: T65 = 8'h96;
    4: T65 = 8'h24;
    5: T65 = 8'h17;
    6: T65 = 8'h70;
    7: T65 = 8'ha4;
    8: T65 = 8'h87;
    9: T65 = 8'hcf;
    10: T65 = 8'ha9;
    11: T65 = 8'h5;
    12: T65 = 8'h1a;
    13: T65 = 8'h40;
    14: T65 = 8'ha5;
    15: T65 = 8'hdb;
    16: T65 = 8'h3d;
    17: T65 = 8'h14;
    18: T65 = 8'h44;
    19: T65 = 8'h59;
    20: T65 = 8'h82;
    21: T65 = 8'h3f;
    22: T65 = 8'h34;
    23: T65 = 8'h66;
    24: T65 = 8'h18;
    25: T65 = 8'he5;
    26: T65 = 8'h84;
    27: T65 = 8'hf5;
    28: T65 = 8'h50;
    29: T65 = 8'hd8;
    30: T65 = 8'hc3;
    31: T65 = 8'h73;
    32: T65 = 8'h5a;
    33: T65 = 8'ha8;
    34: T65 = 8'h9c;
    35: T65 = 8'hcb;
    36: T65 = 8'hb1;
    37: T65 = 8'h78;
    38: T65 = 8'h2;
    39: T65 = 8'hbe;
    40: T65 = 8'hbc;
    41: T65 = 8'h7;
    42: T65 = 8'h64;
    43: T65 = 8'hb9;
    44: T65 = 8'hae;
    45: T65 = 8'hf3;
    46: T65 = 8'ha2;
    47: T65 = 8'ha;
    48: T65 = 8'hed;
    49: T65 = 8'h12;
    50: T65 = 8'hfd;
    51: T65 = 8'he1;
    52: T65 = 8'h8;
    53: T65 = 8'hd0;
    54: T65 = 8'hac;
    55: T65 = 8'hf4;
    56: T65 = 8'hff;
    57: T65 = 8'h7e;
    58: T65 = 8'h65;
    59: T65 = 8'h4f;
    60: T65 = 8'h91;
    61: T65 = 8'heb;
    62: T65 = 8'he4;
    63: T65 = 8'h79;
    64: T65 = 8'h7b;
    65: T65 = 8'hfb;
    66: T65 = 8'h43;
    67: T65 = 8'hfa;
    68: T65 = 8'ha1;
    69: T65 = 8'h0;
    70: T65 = 8'h6b;
    71: T65 = 8'h61;
    72: T65 = 8'hf1;
    73: T65 = 8'h6f;
    74: T65 = 8'hb5;
    75: T65 = 8'h52;
    76: T65 = 8'hf9;
    77: T65 = 8'h21;
    78: T65 = 8'h45;
    79: T65 = 8'h37;
    80: T65 = 8'h3b;
    81: T65 = 8'h99;
    82: T65 = 8'h1d;
    83: T65 = 8'h9;
    84: T65 = 8'hd5;
    85: T65 = 8'ha7;
    86: T65 = 8'h54;
    87: T65 = 8'h5d;
    88: T65 = 8'h1e;
    89: T65 = 8'h2e;
    90: T65 = 8'h5e;
    91: T65 = 8'h4b;
    92: T65 = 8'h97;
    93: T65 = 8'h72;
    94: T65 = 8'h49;
    95: T65 = 8'hde;
    96: T65 = 8'hc5;
    97: T65 = 8'h60;
    98: T65 = 8'hd2;
    99: T65 = 8'h2d;
    100: T65 = 8'h10;
    101: T65 = 8'he3;
    102: T65 = 8'hf8;
    103: T65 = 8'hca;
    104: T65 = 8'h33;
    105: T65 = 8'h98;
    106: T65 = 8'hfc;
    107: T65 = 8'h7d;
    108: T65 = 8'h51;
    109: T65 = 8'hce;
    110: T65 = 8'hd7;
    111: T65 = 8'hba;
    112: T65 = 8'h27;
    113: T65 = 8'h9e;
    114: T65 = 8'hb2;
    115: T65 = 8'hbb;
    116: T65 = 8'h83;
    117: T65 = 8'h88;
    118: T65 = 8'h1;
    119: T65 = 8'h31;
    120: T65 = 8'h32;
    121: T65 = 8'h11;
    122: T65 = 8'h8d;
    123: T65 = 8'h5b;
    124: T65 = 8'h2f;
    125: T65 = 8'h81;
    126: T65 = 8'h3c;
    127: T65 = 8'h63;
    128: T65 = 8'h9a;
    129: T65 = 8'h23;
    130: T65 = 8'h56;
    131: T65 = 8'hab;
    132: T65 = 8'h69;
    133: T65 = 8'h22;
    134: T65 = 8'h26;
    135: T65 = 8'hc8;
    136: T65 = 8'h93;
    137: T65 = 8'h3a;
    138: T65 = 8'h4d;
    139: T65 = 8'h76;
    140: T65 = 8'had;
    141: T65 = 8'hf6;
    142: T65 = 8'h4c;
    143: T65 = 8'hfe;
    144: T65 = 8'h85;
    145: T65 = 8'he8;
    146: T65 = 8'hc4;
    147: T65 = 8'h90;
    148: T65 = 8'hc6;
    149: T65 = 8'h7c;
    150: T65 = 8'h35;
    151: T65 = 8'h4;
    152: T65 = 8'h6c;
    153: T65 = 8'h4a;
    154: T65 = 8'hdf;
    155: T65 = 8'hea;
    156: T65 = 8'h86;
    157: T65 = 8'he6;
    158: T65 = 8'h9d;
    159: T65 = 8'h8b;
    160: T65 = 8'hbd;
    161: T65 = 8'hcd;
    162: T65 = 8'hc7;
    163: T65 = 8'h80;
    164: T65 = 8'hb0;
    165: T65 = 8'h13;
    166: T65 = 8'hd3;
    167: T65 = 8'hec;
    168: T65 = 8'h7f;
    169: T65 = 8'hc0;
    170: T65 = 8'he7;
    171: T65 = 8'h46;
    172: T65 = 8'he9;
    173: T65 = 8'h58;
    174: T65 = 8'h92;
    175: T65 = 8'h2c;
    176: T65 = 8'hb7;
    177: T65 = 8'hc9;
    178: T65 = 8'h16;
    179: T65 = 8'h53;
    180: T65 = 8'hd;
    181: T65 = 8'hd6;
    182: T65 = 8'h74;
    183: T65 = 8'h6d;
    184: T65 = 8'h9f;
    185: T65 = 8'h20;
    186: T65 = 8'h5f;
    187: T65 = 8'he2;
    188: T65 = 8'h8c;
    189: T65 = 8'hdc;
    190: T65 = 8'h39;
    191: T65 = 8'hc;
    192: T65 = 8'hdd;
    193: T65 = 8'h1f;
    194: T65 = 8'hd1;
    195: T65 = 8'hb6;
    196: T65 = 8'h8f;
    197: T65 = 8'h5c;
    198: T65 = 8'h95;
    199: T65 = 8'hb8;
    200: T65 = 8'h94;
    201: T65 = 8'h3e;
    202: T65 = 8'h71;
    203: T65 = 8'h41;
    204: T65 = 8'h25;
    205: T65 = 8'h1b;
    206: T65 = 8'h6a;
    207: T65 = 8'ha6;
    208: T65 = 8'h3;
    209: T65 = 8'he;
    210: T65 = 8'hcc;
    211: T65 = 8'h48;
    212: T65 = 8'h15;
    213: T65 = 8'h29;
    214: T65 = 8'h38;
    215: T65 = 8'h42;
    216: T65 = 8'h1c;
    217: T65 = 8'hc1;
    218: T65 = 8'h28;
    219: T65 = 8'hd9;
    220: T65 = 8'h19;
    221: T65 = 8'h36;
    222: T65 = 8'hb3;
    223: T65 = 8'h75;
    224: T65 = 8'hee;
    225: T65 = 8'h57;
    226: T65 = 8'hf0;
    227: T65 = 8'h9b;
    228: T65 = 8'hb4;
    229: T65 = 8'haa;
    230: T65 = 8'hf2;
    231: T65 = 8'hd4;
    232: T65 = 8'hbf;
    233: T65 = 8'ha3;
    234: T65 = 8'h4e;
    235: T65 = 8'hda;
    236: T65 = 8'h89;
    237: T65 = 8'hc2;
    238: T65 = 8'haf;
    239: T65 = 8'h6e;
    240: T65 = 8'h2b;
    241: T65 = 8'h77;
    242: T65 = 8'he0;
    243: T65 = 8'h47;
    244: T65 = 8'h7a;
    245: T65 = 8'h8e;
    246: T65 = 8'h2a;
    247: T65 = 8'ha0;
    248: T65 = 8'h68;
    249: T65 = 8'h30;
    250: T65 = 8'hf7;
    251: T65 = 8'h67;
    252: T65 = 8'hf;
    253: T65 = 8'hb;
    254: T65 = 8'h8a;
    255: T65 = 8'hef;
`ifndef SYNTHESIS
    default: T65 = {1{$random}};
`else
    default: T65 = 8'bx;
`endif
  endcase
  assign T66 = keyLen[3'h5:1'h0];
  assign io_halted = T0;
  assign T0 = T1 & io_lock;
  assign T1 = state == 2'h0;
  assign io_hashOut_bits_tag = keyTag;
  assign T20 = T5 ? io_keyInfo_bits_tag : keyTag;
  assign io_hashOut_bits_len = keyLen;
  assign io_hashOut_bits_hash2 = T48;
  assign T48 = PearsonHasher_1_io_result_bits[4'h9:1'h0];
  assign io_hashOut_bits_hash1 = T49;
  assign T49 = PearsonHasher_0_io_result_bits[4'h9:1'h0];
  assign io_hashOut_valid = T21;
  assign T21 = state == 2'h2;
  assign io_keyInfo_ready = T22;
  assign T22 = T24 & T23;
  assign T23 = io_lock ^ 1'h1;
  assign T24 = state == 2'h0;
  assign io_keyData_ready = T25;
  assign T25 = state == 2'h1;
  assign io_keyWrite = keyWrite;
  assign T50 = reset ? 1'h0 : T26;
  assign T26 = T19 ? 1'h0 : T27;
  assign T27 = T30 ? 1'h1 : T28;
  assign T28 = T9 ? 1'h1 : T29;
  assign T29 = T17 ? 1'h0 : keyWrite;
  assign T30 = T16 & T31;
  assign T31 = T33 & T32;
  assign T32 = byteOff == 2'h3;
  assign byteOff = index[1'h1:1'h0];
  assign T33 = T10 ^ 1'h1;
  assign io_keyWriteData = keyWriteData;
  assign T51 = T52[5'h1f:1'h0];
  assign T52 = reset ? 39'h0 : T34;
  assign T34 = T40 ? T38 : T53;
  assign T53 = {7'h0, T35};
  assign T35 = T36 ? T54 : keyWriteData;
  assign T54 = {24'h0, io_keyData_bits};
  assign T36 = T16 & T37;
  assign T37 = byteOff == 2'h0;
  assign T38 = T55 | T39;
  assign T39 = io_keyData_bits << inputShift;
  assign inputShift = {byteOff, 3'h0};
  assign T55 = {7'h0, keyWriteData};
  assign T40 = T16 & T41;
  assign T41 = T37 ^ 1'h1;
  assign io_keyWriteAddr = keyWriteAddr;
  assign T56 = reset ? 6'h0 : T42;
  assign T42 = T30 ? T45 : T43;
  assign T43 = T9 ? T44 : keyWriteAddr;
  assign T44 = index[3'h7:2'h2];
  assign T45 = index[3'h7:2'h2];
  PearsonHasher PearsonHasher_0(.clk(clk), .reset(reset),
       .io_keyData_valid( hashInputValid ),
       .io_keyData_bits( io_keyData_bits ),
       .io_keyLen( T66 ),
       .io_romAddr_1( PearsonHasher_0_io_romAddr_1 ),
       .io_romAddr_0( PearsonHasher_0_io_romAddr_0 ),
       .io_romData_1( T65 ),
       .io_romData_0( T64 ),
       //.io_result_valid(  )
       .io_result_bits( PearsonHasher_0_io_result_bits ),
       .io_restart( restart )
  );
  PearsonHasher PearsonHasher_1(.clk(clk), .reset(reset),
       .io_keyData_valid( hashInputValid ),
       .io_keyData_bits( io_keyData_bits ),
       .io_keyLen( T62 ),
       .io_romAddr_1( PearsonHasher_1_io_romAddr_1 ),
       .io_romAddr_0( PearsonHasher_1_io_romAddr_0 ),
       .io_romData_1( T61 ),
       .io_romData_0( T60 ),
       //.io_result_valid(  )
       .io_result_bits( PearsonHasher_1_io_result_bits ),
       .io_restart( restart )
  );

  always @(posedge clk) begin
    if(reset) begin
      restart <= 1'h0;
    end else if(T18) begin
      restart <= 1'h1;
    end else if(T8) begin
      restart <= 1'h0;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T18) begin
      state <= 2'h0;
    end else if(T9) begin
      state <= 2'h2;
    end else if(T5) begin
      state <= 2'h1;
    end
    if(T5) begin
      keyLen <= io_keyInfo_bits_len;
    end
    if(reset) begin
      index <= 8'h0;
    end else if(T16) begin
      index <= T15;
    end else if(T5) begin
      index <= 8'h0;
    end
    if(T5) begin
      keyTag <= io_keyInfo_bits_tag;
    end
    if(reset) begin
      keyWrite <= 1'h0;
    end else if(T19) begin
      keyWrite <= 1'h0;
    end else if(T30) begin
      keyWrite <= 1'h1;
    end else if(T9) begin
      keyWrite <= 1'h1;
    end else if(T17) begin
      keyWrite <= 1'h0;
    end
    keyWriteData <= T51;
    if(reset) begin
      keyWriteAddr <= 6'h0;
    end else if(T30) begin
      keyWriteAddr <= T45;
    end else if(T9) begin
      keyWriteAddr <= T44;
    end
  end
endmodule

module KeyCompare(input clk, input reset,
    output[5:0] io_curKeyAddr,
    input [31:0] io_curKeyData,
    output[15:0] io_allKeyAddr,
    input [31:0] io_allKeyData,
    output[9:0] io_lenAddr,
    input [7:0] io_lenData,
    output io_hashIn_ready,
    input  io_hashIn_valid,
    input [9:0] io_hashIn_bits_hash1,
    input [9:0] io_hashIn_bits_hash2,
    input [7:0] io_hashIn_bits_len,
    input [3:0] io_hashIn_bits_tag,
    input  io_hashOut_ready,
    output io_hashOut_valid,
    output[3:0] io_hashOut_bits_tag,
    output[9:0] io_hashOut_bits_hash,
    output io_hashOut_bits_found,
    input  io_findAvailable,
    input  io_resetCounts
);

  reg  hashFound;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg [2:0] state;
  wire[2:0] T10343;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [7:0] curInfo_len;
  wire[7:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  checkFirst;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [3:0] hashCount2;
  wire[3:0] T10344;
  wire[3:0] T39;
  wire[3:0] T40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[3:0] T45;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[3:0] T48;
  wire[3:0] T49;
  reg [3:0] counts_0;
  wire[3:0] T10345;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T52;
  wire[3:0] T53;
  wire[3:0] T10346;
  wire T54;
  wire[4:0] T55;
  wire[4:0] T56;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[3:0] T66;
  wire T67;
  wire[9:0] T68;
  wire[9:0] curHash;
  reg [9:0] curInfo_hash2;
  wire[9:0] T69;
  reg [9:0] curInfo_hash1;
  wire[9:0] T70;
  wire[3:0] T71;
  reg [3:0] counts_2;
  wire[3:0] T10347;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire[1023:0] T76;
  reg [3:0] counts_3;
  wire[3:0] T10348;
  wire[3:0] T77;
  wire[3:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[3:0] T83;
  wire[3:0] T84;
  reg [3:0] counts_4;
  wire[3:0] T10349;
  wire[3:0] T85;
  wire[3:0] T86;
  wire T87;
  wire T88;
  reg [3:0] counts_5;
  wire[3:0] T10350;
  wire[3:0] T89;
  wire[3:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  reg [3:0] counts_6;
  wire[3:0] T10351;
  wire[3:0] T95;
  wire[3:0] T96;
  wire T97;
  wire T98;
  reg [3:0] counts_7;
  wire[3:0] T10352;
  wire[3:0] T99;
  wire[3:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] T108;
  reg [3:0] counts_8;
  wire[3:0] T10353;
  wire[3:0] T109;
  wire[3:0] T110;
  wire T111;
  wire T112;
  reg [3:0] counts_9;
  wire[3:0] T10354;
  wire[3:0] T113;
  wire[3:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire[3:0] T118;
  reg [3:0] counts_10;
  wire[3:0] T10355;
  wire[3:0] T119;
  wire[3:0] T120;
  wire T121;
  wire T122;
  reg [3:0] counts_11;
  wire[3:0] T10356;
  wire[3:0] T123;
  wire[3:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[3:0] T129;
  wire[3:0] T130;
  reg [3:0] counts_12;
  wire[3:0] T10357;
  wire[3:0] T131;
  wire[3:0] T132;
  wire T133;
  wire T134;
  reg [3:0] counts_13;
  wire[3:0] T10358;
  wire[3:0] T135;
  wire[3:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire[3:0] T140;
  reg [3:0] counts_14;
  wire[3:0] T10359;
  wire[3:0] T141;
  wire[3:0] T142;
  wire T143;
  wire T144;
  reg [3:0] counts_15;
  wire[3:0] T10360;
  wire[3:0] T145;
  wire[3:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire[3:0] T153;
  wire[3:0] T154;
  wire[3:0] T155;
  wire[3:0] T156;
  reg [3:0] counts_16;
  wire[3:0] T10361;
  wire[3:0] T157;
  wire[3:0] T158;
  wire T159;
  wire T160;
  reg [3:0] counts_17;
  wire[3:0] T10362;
  wire[3:0] T161;
  wire[3:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire[3:0] T166;
  reg [3:0] counts_18;
  wire[3:0] T10363;
  wire[3:0] T167;
  wire[3:0] T168;
  wire T169;
  wire T170;
  reg [3:0] counts_19;
  wire[3:0] T10364;
  wire[3:0] T171;
  wire[3:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire[3:0] T177;
  wire[3:0] T178;
  reg [3:0] counts_20;
  wire[3:0] T10365;
  wire[3:0] T179;
  wire[3:0] T180;
  wire T181;
  wire T182;
  reg [3:0] counts_21;
  wire[3:0] T10366;
  wire[3:0] T183;
  wire[3:0] T184;
  wire T185;
  wire T186;
  wire T187;
  wire[3:0] T188;
  reg [3:0] counts_22;
  wire[3:0] T10367;
  wire[3:0] T189;
  wire[3:0] T190;
  wire T191;
  wire T192;
  reg [3:0] counts_23;
  wire[3:0] T10368;
  wire[3:0] T193;
  wire[3:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire[3:0] T200;
  wire[3:0] T201;
  wire[3:0] T202;
  reg [3:0] counts_24;
  wire[3:0] T10369;
  wire[3:0] T203;
  wire[3:0] T204;
  wire T205;
  wire T206;
  reg [3:0] counts_25;
  wire[3:0] T10370;
  wire[3:0] T207;
  wire[3:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire[3:0] T212;
  reg [3:0] counts_26;
  wire[3:0] T10371;
  wire[3:0] T213;
  wire[3:0] T214;
  wire T215;
  wire T216;
  reg [3:0] counts_27;
  wire[3:0] T10372;
  wire[3:0] T217;
  wire[3:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] T224;
  reg [3:0] counts_28;
  wire[3:0] T10373;
  wire[3:0] T225;
  wire[3:0] T226;
  wire T227;
  wire T228;
  reg [3:0] counts_29;
  wire[3:0] T10374;
  wire[3:0] T229;
  wire[3:0] T230;
  wire T231;
  wire T232;
  wire T233;
  wire[3:0] T234;
  reg [3:0] counts_30;
  wire[3:0] T10375;
  wire[3:0] T235;
  wire[3:0] T236;
  wire T237;
  wire T238;
  reg [3:0] counts_31;
  wire[3:0] T10376;
  wire[3:0] T239;
  wire[3:0] T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[3:0] T248;
  wire[3:0] T249;
  wire[3:0] T250;
  wire[3:0] T251;
  wire[3:0] T252;
  reg [3:0] counts_32;
  wire[3:0] T10377;
  wire[3:0] T253;
  wire[3:0] T254;
  wire T255;
  wire T256;
  reg [3:0] counts_33;
  wire[3:0] T10378;
  wire[3:0] T257;
  wire[3:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire[3:0] T262;
  reg [3:0] counts_34;
  wire[3:0] T10379;
  wire[3:0] T263;
  wire[3:0] T264;
  wire T265;
  wire T266;
  reg [3:0] counts_35;
  wire[3:0] T10380;
  wire[3:0] T267;
  wire[3:0] T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[3:0] T273;
  wire[3:0] T274;
  reg [3:0] counts_36;
  wire[3:0] T10381;
  wire[3:0] T275;
  wire[3:0] T276;
  wire T277;
  wire T278;
  reg [3:0] counts_37;
  wire[3:0] T10382;
  wire[3:0] T279;
  wire[3:0] T280;
  wire T281;
  wire T282;
  wire T283;
  wire[3:0] T284;
  reg [3:0] counts_38;
  wire[3:0] T10383;
  wire[3:0] T285;
  wire[3:0] T286;
  wire T287;
  wire T288;
  reg [3:0] counts_39;
  wire[3:0] T10384;
  wire[3:0] T289;
  wire[3:0] T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire[3:0] T296;
  wire[3:0] T297;
  wire[3:0] T298;
  reg [3:0] counts_40;
  wire[3:0] T10385;
  wire[3:0] T299;
  wire[3:0] T300;
  wire T301;
  wire T302;
  reg [3:0] counts_41;
  wire[3:0] T10386;
  wire[3:0] T303;
  wire[3:0] T304;
  wire T305;
  wire T306;
  wire T307;
  wire[3:0] T308;
  reg [3:0] counts_42;
  wire[3:0] T10387;
  wire[3:0] T309;
  wire[3:0] T310;
  wire T311;
  wire T312;
  reg [3:0] counts_43;
  wire[3:0] T10388;
  wire[3:0] T313;
  wire[3:0] T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire[3:0] T319;
  wire[3:0] T320;
  reg [3:0] counts_44;
  wire[3:0] T10389;
  wire[3:0] T321;
  wire[3:0] T322;
  wire T323;
  wire T324;
  reg [3:0] counts_45;
  wire[3:0] T10390;
  wire[3:0] T325;
  wire[3:0] T326;
  wire T327;
  wire T328;
  wire T329;
  wire[3:0] T330;
  reg [3:0] counts_46;
  wire[3:0] T10391;
  wire[3:0] T331;
  wire[3:0] T332;
  wire T333;
  wire T334;
  reg [3:0] counts_47;
  wire[3:0] T10392;
  wire[3:0] T335;
  wire[3:0] T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire[3:0] T343;
  wire[3:0] T344;
  wire[3:0] T345;
  wire[3:0] T346;
  reg [3:0] counts_48;
  wire[3:0] T10393;
  wire[3:0] T347;
  wire[3:0] T348;
  wire T349;
  wire T350;
  reg [3:0] counts_49;
  wire[3:0] T10394;
  wire[3:0] T351;
  wire[3:0] T352;
  wire T353;
  wire T354;
  wire T355;
  wire[3:0] T356;
  reg [3:0] counts_50;
  wire[3:0] T10395;
  wire[3:0] T357;
  wire[3:0] T358;
  wire T359;
  wire T360;
  reg [3:0] counts_51;
  wire[3:0] T10396;
  wire[3:0] T361;
  wire[3:0] T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire[3:0] T367;
  wire[3:0] T368;
  reg [3:0] counts_52;
  wire[3:0] T10397;
  wire[3:0] T369;
  wire[3:0] T370;
  wire T371;
  wire T372;
  reg [3:0] counts_53;
  wire[3:0] T10398;
  wire[3:0] T373;
  wire[3:0] T374;
  wire T375;
  wire T376;
  wire T377;
  wire[3:0] T378;
  reg [3:0] counts_54;
  wire[3:0] T10399;
  wire[3:0] T379;
  wire[3:0] T380;
  wire T381;
  wire T382;
  reg [3:0] counts_55;
  wire[3:0] T10400;
  wire[3:0] T383;
  wire[3:0] T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire[3:0] T390;
  wire[3:0] T391;
  wire[3:0] T392;
  reg [3:0] counts_56;
  wire[3:0] T10401;
  wire[3:0] T393;
  wire[3:0] T394;
  wire T395;
  wire T396;
  reg [3:0] counts_57;
  wire[3:0] T10402;
  wire[3:0] T397;
  wire[3:0] T398;
  wire T399;
  wire T400;
  wire T401;
  wire[3:0] T402;
  reg [3:0] counts_58;
  wire[3:0] T10403;
  wire[3:0] T403;
  wire[3:0] T404;
  wire T405;
  wire T406;
  reg [3:0] counts_59;
  wire[3:0] T10404;
  wire[3:0] T407;
  wire[3:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire[3:0] T413;
  wire[3:0] T414;
  reg [3:0] counts_60;
  wire[3:0] T10405;
  wire[3:0] T415;
  wire[3:0] T416;
  wire T417;
  wire T418;
  reg [3:0] counts_61;
  wire[3:0] T10406;
  wire[3:0] T419;
  wire[3:0] T420;
  wire T421;
  wire T422;
  wire T423;
  wire[3:0] T424;
  reg [3:0] counts_62;
  wire[3:0] T10407;
  wire[3:0] T425;
  wire[3:0] T426;
  wire T427;
  wire T428;
  reg [3:0] counts_63;
  wire[3:0] T10408;
  wire[3:0] T429;
  wire[3:0] T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire[3:0] T439;
  wire[3:0] T440;
  wire[3:0] T441;
  wire[3:0] T442;
  wire[3:0] T443;
  wire[3:0] T444;
  reg [3:0] counts_64;
  wire[3:0] T10409;
  wire[3:0] T445;
  wire[3:0] T446;
  wire T447;
  wire T448;
  reg [3:0] counts_65;
  wire[3:0] T10410;
  wire[3:0] T449;
  wire[3:0] T450;
  wire T451;
  wire T452;
  wire T453;
  wire[3:0] T454;
  reg [3:0] counts_66;
  wire[3:0] T10411;
  wire[3:0] T455;
  wire[3:0] T456;
  wire T457;
  wire T458;
  reg [3:0] counts_67;
  wire[3:0] T10412;
  wire[3:0] T459;
  wire[3:0] T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  reg [3:0] counts_68;
  wire[3:0] T10413;
  wire[3:0] T467;
  wire[3:0] T468;
  wire T469;
  wire T470;
  reg [3:0] counts_69;
  wire[3:0] T10414;
  wire[3:0] T471;
  wire[3:0] T472;
  wire T473;
  wire T474;
  wire T475;
  wire[3:0] T476;
  reg [3:0] counts_70;
  wire[3:0] T10415;
  wire[3:0] T477;
  wire[3:0] T478;
  wire T479;
  wire T480;
  reg [3:0] counts_71;
  wire[3:0] T10416;
  wire[3:0] T481;
  wire[3:0] T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[3:0] T488;
  wire[3:0] T489;
  wire[3:0] T490;
  reg [3:0] counts_72;
  wire[3:0] T10417;
  wire[3:0] T491;
  wire[3:0] T492;
  wire T493;
  wire T494;
  reg [3:0] counts_73;
  wire[3:0] T10418;
  wire[3:0] T495;
  wire[3:0] T496;
  wire T497;
  wire T498;
  wire T499;
  wire[3:0] T500;
  reg [3:0] counts_74;
  wire[3:0] T10419;
  wire[3:0] T501;
  wire[3:0] T502;
  wire T503;
  wire T504;
  reg [3:0] counts_75;
  wire[3:0] T10420;
  wire[3:0] T505;
  wire[3:0] T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire[3:0] T511;
  wire[3:0] T512;
  reg [3:0] counts_76;
  wire[3:0] T10421;
  wire[3:0] T513;
  wire[3:0] T514;
  wire T515;
  wire T516;
  reg [3:0] counts_77;
  wire[3:0] T10422;
  wire[3:0] T517;
  wire[3:0] T518;
  wire T519;
  wire T520;
  wire T521;
  wire[3:0] T522;
  reg [3:0] counts_78;
  wire[3:0] T10423;
  wire[3:0] T523;
  wire[3:0] T524;
  wire T525;
  wire T526;
  reg [3:0] counts_79;
  wire[3:0] T10424;
  wire[3:0] T527;
  wire[3:0] T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire[3:0] T535;
  wire[3:0] T536;
  wire[3:0] T537;
  wire[3:0] T538;
  reg [3:0] counts_80;
  wire[3:0] T10425;
  wire[3:0] T539;
  wire[3:0] T540;
  wire T541;
  wire T542;
  reg [3:0] counts_81;
  wire[3:0] T10426;
  wire[3:0] T543;
  wire[3:0] T544;
  wire T545;
  wire T546;
  wire T547;
  wire[3:0] T548;
  reg [3:0] counts_82;
  wire[3:0] T10427;
  wire[3:0] T549;
  wire[3:0] T550;
  wire T551;
  wire T552;
  reg [3:0] counts_83;
  wire[3:0] T10428;
  wire[3:0] T553;
  wire[3:0] T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire[3:0] T559;
  wire[3:0] T560;
  reg [3:0] counts_84;
  wire[3:0] T10429;
  wire[3:0] T561;
  wire[3:0] T562;
  wire T563;
  wire T564;
  reg [3:0] counts_85;
  wire[3:0] T10430;
  wire[3:0] T565;
  wire[3:0] T566;
  wire T567;
  wire T568;
  wire T569;
  wire[3:0] T570;
  reg [3:0] counts_86;
  wire[3:0] T10431;
  wire[3:0] T571;
  wire[3:0] T572;
  wire T573;
  wire T574;
  reg [3:0] counts_87;
  wire[3:0] T10432;
  wire[3:0] T575;
  wire[3:0] T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire[3:0] T582;
  wire[3:0] T583;
  wire[3:0] T584;
  reg [3:0] counts_88;
  wire[3:0] T10433;
  wire[3:0] T585;
  wire[3:0] T586;
  wire T587;
  wire T588;
  reg [3:0] counts_89;
  wire[3:0] T10434;
  wire[3:0] T589;
  wire[3:0] T590;
  wire T591;
  wire T592;
  wire T593;
  wire[3:0] T594;
  reg [3:0] counts_90;
  wire[3:0] T10435;
  wire[3:0] T595;
  wire[3:0] T596;
  wire T597;
  wire T598;
  reg [3:0] counts_91;
  wire[3:0] T10436;
  wire[3:0] T599;
  wire[3:0] T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire[3:0] T605;
  wire[3:0] T606;
  reg [3:0] counts_92;
  wire[3:0] T10437;
  wire[3:0] T607;
  wire[3:0] T608;
  wire T609;
  wire T610;
  reg [3:0] counts_93;
  wire[3:0] T10438;
  wire[3:0] T611;
  wire[3:0] T612;
  wire T613;
  wire T614;
  wire T615;
  wire[3:0] T616;
  reg [3:0] counts_94;
  wire[3:0] T10439;
  wire[3:0] T617;
  wire[3:0] T618;
  wire T619;
  wire T620;
  reg [3:0] counts_95;
  wire[3:0] T10440;
  wire[3:0] T621;
  wire[3:0] T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire[3:0] T630;
  wire[3:0] T631;
  wire[3:0] T632;
  wire[3:0] T633;
  wire[3:0] T634;
  reg [3:0] counts_96;
  wire[3:0] T10441;
  wire[3:0] T635;
  wire[3:0] T636;
  wire T637;
  wire T638;
  reg [3:0] counts_97;
  wire[3:0] T10442;
  wire[3:0] T639;
  wire[3:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[3:0] T644;
  reg [3:0] counts_98;
  wire[3:0] T10443;
  wire[3:0] T645;
  wire[3:0] T646;
  wire T647;
  wire T648;
  reg [3:0] counts_99;
  wire[3:0] T10444;
  wire[3:0] T649;
  wire[3:0] T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire[3:0] T655;
  wire[3:0] T656;
  reg [3:0] counts_100;
  wire[3:0] T10445;
  wire[3:0] T657;
  wire[3:0] T658;
  wire T659;
  wire T660;
  reg [3:0] counts_101;
  wire[3:0] T10446;
  wire[3:0] T661;
  wire[3:0] T662;
  wire T663;
  wire T664;
  wire T665;
  wire[3:0] T666;
  reg [3:0] counts_102;
  wire[3:0] T10447;
  wire[3:0] T667;
  wire[3:0] T668;
  wire T669;
  wire T670;
  reg [3:0] counts_103;
  wire[3:0] T10448;
  wire[3:0] T671;
  wire[3:0] T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire[3:0] T678;
  wire[3:0] T679;
  wire[3:0] T680;
  reg [3:0] counts_104;
  wire[3:0] T10449;
  wire[3:0] T681;
  wire[3:0] T682;
  wire T683;
  wire T684;
  reg [3:0] counts_105;
  wire[3:0] T10450;
  wire[3:0] T685;
  wire[3:0] T686;
  wire T687;
  wire T688;
  wire T689;
  wire[3:0] T690;
  reg [3:0] counts_106;
  wire[3:0] T10451;
  wire[3:0] T691;
  wire[3:0] T692;
  wire T693;
  wire T694;
  reg [3:0] counts_107;
  wire[3:0] T10452;
  wire[3:0] T695;
  wire[3:0] T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire[3:0] T701;
  wire[3:0] T702;
  reg [3:0] counts_108;
  wire[3:0] T10453;
  wire[3:0] T703;
  wire[3:0] T704;
  wire T705;
  wire T706;
  reg [3:0] counts_109;
  wire[3:0] T10454;
  wire[3:0] T707;
  wire[3:0] T708;
  wire T709;
  wire T710;
  wire T711;
  wire[3:0] T712;
  reg [3:0] counts_110;
  wire[3:0] T10455;
  wire[3:0] T713;
  wire[3:0] T714;
  wire T715;
  wire T716;
  reg [3:0] counts_111;
  wire[3:0] T10456;
  wire[3:0] T717;
  wire[3:0] T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire[3:0] T725;
  wire[3:0] T726;
  wire[3:0] T727;
  wire[3:0] T728;
  reg [3:0] counts_112;
  wire[3:0] T10457;
  wire[3:0] T729;
  wire[3:0] T730;
  wire T731;
  wire T732;
  reg [3:0] counts_113;
  wire[3:0] T10458;
  wire[3:0] T733;
  wire[3:0] T734;
  wire T735;
  wire T736;
  wire T737;
  wire[3:0] T738;
  reg [3:0] counts_114;
  wire[3:0] T10459;
  wire[3:0] T739;
  wire[3:0] T740;
  wire T741;
  wire T742;
  reg [3:0] counts_115;
  wire[3:0] T10460;
  wire[3:0] T743;
  wire[3:0] T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire[3:0] T749;
  wire[3:0] T750;
  reg [3:0] counts_116;
  wire[3:0] T10461;
  wire[3:0] T751;
  wire[3:0] T752;
  wire T753;
  wire T754;
  reg [3:0] counts_117;
  wire[3:0] T10462;
  wire[3:0] T755;
  wire[3:0] T756;
  wire T757;
  wire T758;
  wire T759;
  wire[3:0] T760;
  reg [3:0] counts_118;
  wire[3:0] T10463;
  wire[3:0] T761;
  wire[3:0] T762;
  wire T763;
  wire T764;
  reg [3:0] counts_119;
  wire[3:0] T10464;
  wire[3:0] T765;
  wire[3:0] T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[3:0] T772;
  wire[3:0] T773;
  wire[3:0] T774;
  reg [3:0] counts_120;
  wire[3:0] T10465;
  wire[3:0] T775;
  wire[3:0] T776;
  wire T777;
  wire T778;
  reg [3:0] counts_121;
  wire[3:0] T10466;
  wire[3:0] T779;
  wire[3:0] T780;
  wire T781;
  wire T782;
  wire T783;
  wire[3:0] T784;
  reg [3:0] counts_122;
  wire[3:0] T10467;
  wire[3:0] T785;
  wire[3:0] T786;
  wire T787;
  wire T788;
  reg [3:0] counts_123;
  wire[3:0] T10468;
  wire[3:0] T789;
  wire[3:0] T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire[3:0] T795;
  wire[3:0] T796;
  reg [3:0] counts_124;
  wire[3:0] T10469;
  wire[3:0] T797;
  wire[3:0] T798;
  wire T799;
  wire T800;
  reg [3:0] counts_125;
  wire[3:0] T10470;
  wire[3:0] T801;
  wire[3:0] T802;
  wire T803;
  wire T804;
  wire T805;
  wire[3:0] T806;
  reg [3:0] counts_126;
  wire[3:0] T10471;
  wire[3:0] T807;
  wire[3:0] T808;
  wire T809;
  wire T810;
  reg [3:0] counts_127;
  wire[3:0] T10472;
  wire[3:0] T811;
  wire[3:0] T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire[3:0] T822;
  wire[3:0] T823;
  wire[3:0] T824;
  wire[3:0] T825;
  wire[3:0] T826;
  wire[3:0] T827;
  wire[3:0] T828;
  reg [3:0] counts_128;
  wire[3:0] T10473;
  wire[3:0] T829;
  wire[3:0] T830;
  wire T831;
  wire T832;
  reg [3:0] counts_129;
  wire[3:0] T10474;
  wire[3:0] T833;
  wire[3:0] T834;
  wire T835;
  wire T836;
  wire T837;
  wire[3:0] T838;
  reg [3:0] counts_130;
  wire[3:0] T10475;
  wire[3:0] T839;
  wire[3:0] T840;
  wire T841;
  wire T842;
  reg [3:0] counts_131;
  wire[3:0] T10476;
  wire[3:0] T843;
  wire[3:0] T844;
  wire T845;
  wire T846;
  wire T847;
  wire T848;
  wire[3:0] T849;
  wire[3:0] T850;
  reg [3:0] counts_132;
  wire[3:0] T10477;
  wire[3:0] T851;
  wire[3:0] T852;
  wire T853;
  wire T854;
  reg [3:0] counts_133;
  wire[3:0] T10478;
  wire[3:0] T855;
  wire[3:0] T856;
  wire T857;
  wire T858;
  wire T859;
  wire[3:0] T860;
  reg [3:0] counts_134;
  wire[3:0] T10479;
  wire[3:0] T861;
  wire[3:0] T862;
  wire T863;
  wire T864;
  reg [3:0] counts_135;
  wire[3:0] T10480;
  wire[3:0] T865;
  wire[3:0] T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire[3:0] T872;
  wire[3:0] T873;
  wire[3:0] T874;
  reg [3:0] counts_136;
  wire[3:0] T10481;
  wire[3:0] T875;
  wire[3:0] T876;
  wire T877;
  wire T878;
  reg [3:0] counts_137;
  wire[3:0] T10482;
  wire[3:0] T879;
  wire[3:0] T880;
  wire T881;
  wire T882;
  wire T883;
  wire[3:0] T884;
  reg [3:0] counts_138;
  wire[3:0] T10483;
  wire[3:0] T885;
  wire[3:0] T886;
  wire T887;
  wire T888;
  reg [3:0] counts_139;
  wire[3:0] T10484;
  wire[3:0] T889;
  wire[3:0] T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire[3:0] T895;
  wire[3:0] T896;
  reg [3:0] counts_140;
  wire[3:0] T10485;
  wire[3:0] T897;
  wire[3:0] T898;
  wire T899;
  wire T900;
  reg [3:0] counts_141;
  wire[3:0] T10486;
  wire[3:0] T901;
  wire[3:0] T902;
  wire T903;
  wire T904;
  wire T905;
  wire[3:0] T906;
  reg [3:0] counts_142;
  wire[3:0] T10487;
  wire[3:0] T907;
  wire[3:0] T908;
  wire T909;
  wire T910;
  reg [3:0] counts_143;
  wire[3:0] T10488;
  wire[3:0] T911;
  wire[3:0] T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire[3:0] T919;
  wire[3:0] T920;
  wire[3:0] T921;
  wire[3:0] T922;
  reg [3:0] counts_144;
  wire[3:0] T10489;
  wire[3:0] T923;
  wire[3:0] T924;
  wire T925;
  wire T926;
  reg [3:0] counts_145;
  wire[3:0] T10490;
  wire[3:0] T927;
  wire[3:0] T928;
  wire T929;
  wire T930;
  wire T931;
  wire[3:0] T932;
  reg [3:0] counts_146;
  wire[3:0] T10491;
  wire[3:0] T933;
  wire[3:0] T934;
  wire T935;
  wire T936;
  reg [3:0] counts_147;
  wire[3:0] T10492;
  wire[3:0] T937;
  wire[3:0] T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire[3:0] T943;
  wire[3:0] T944;
  reg [3:0] counts_148;
  wire[3:0] T10493;
  wire[3:0] T945;
  wire[3:0] T946;
  wire T947;
  wire T948;
  reg [3:0] counts_149;
  wire[3:0] T10494;
  wire[3:0] T949;
  wire[3:0] T950;
  wire T951;
  wire T952;
  wire T953;
  wire[3:0] T954;
  reg [3:0] counts_150;
  wire[3:0] T10495;
  wire[3:0] T955;
  wire[3:0] T956;
  wire T957;
  wire T958;
  reg [3:0] counts_151;
  wire[3:0] T10496;
  wire[3:0] T959;
  wire[3:0] T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire[3:0] T966;
  wire[3:0] T967;
  wire[3:0] T968;
  reg [3:0] counts_152;
  wire[3:0] T10497;
  wire[3:0] T969;
  wire[3:0] T970;
  wire T971;
  wire T972;
  reg [3:0] counts_153;
  wire[3:0] T10498;
  wire[3:0] T973;
  wire[3:0] T974;
  wire T975;
  wire T976;
  wire T977;
  wire[3:0] T978;
  reg [3:0] counts_154;
  wire[3:0] T10499;
  wire[3:0] T979;
  wire[3:0] T980;
  wire T981;
  wire T982;
  reg [3:0] counts_155;
  wire[3:0] T10500;
  wire[3:0] T983;
  wire[3:0] T984;
  wire T985;
  wire T986;
  wire T987;
  wire T988;
  wire[3:0] T989;
  wire[3:0] T990;
  reg [3:0] counts_156;
  wire[3:0] T10501;
  wire[3:0] T991;
  wire[3:0] T992;
  wire T993;
  wire T994;
  reg [3:0] counts_157;
  wire[3:0] T10502;
  wire[3:0] T995;
  wire[3:0] T996;
  wire T997;
  wire T998;
  wire T999;
  wire[3:0] T1000;
  reg [3:0] counts_158;
  wire[3:0] T10503;
  wire[3:0] T1001;
  wire[3:0] T1002;
  wire T1003;
  wire T1004;
  reg [3:0] counts_159;
  wire[3:0] T10504;
  wire[3:0] T1005;
  wire[3:0] T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire[3:0] T1014;
  wire[3:0] T1015;
  wire[3:0] T1016;
  wire[3:0] T1017;
  wire[3:0] T1018;
  reg [3:0] counts_160;
  wire[3:0] T10505;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire T1021;
  wire T1022;
  reg [3:0] counts_161;
  wire[3:0] T10506;
  wire[3:0] T1023;
  wire[3:0] T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[3:0] T1028;
  reg [3:0] counts_162;
  wire[3:0] T10507;
  wire[3:0] T1029;
  wire[3:0] T1030;
  wire T1031;
  wire T1032;
  reg [3:0] counts_163;
  wire[3:0] T10508;
  wire[3:0] T1033;
  wire[3:0] T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire[3:0] T1039;
  wire[3:0] T1040;
  reg [3:0] counts_164;
  wire[3:0] T10509;
  wire[3:0] T1041;
  wire[3:0] T1042;
  wire T1043;
  wire T1044;
  reg [3:0] counts_165;
  wire[3:0] T10510;
  wire[3:0] T1045;
  wire[3:0] T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire[3:0] T1050;
  reg [3:0] counts_166;
  wire[3:0] T10511;
  wire[3:0] T1051;
  wire[3:0] T1052;
  wire T1053;
  wire T1054;
  reg [3:0] counts_167;
  wire[3:0] T10512;
  wire[3:0] T1055;
  wire[3:0] T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire[3:0] T1062;
  wire[3:0] T1063;
  wire[3:0] T1064;
  reg [3:0] counts_168;
  wire[3:0] T10513;
  wire[3:0] T1065;
  wire[3:0] T1066;
  wire T1067;
  wire T1068;
  reg [3:0] counts_169;
  wire[3:0] T10514;
  wire[3:0] T1069;
  wire[3:0] T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire[3:0] T1074;
  reg [3:0] counts_170;
  wire[3:0] T10515;
  wire[3:0] T1075;
  wire[3:0] T1076;
  wire T1077;
  wire T1078;
  reg [3:0] counts_171;
  wire[3:0] T10516;
  wire[3:0] T1079;
  wire[3:0] T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire[3:0] T1085;
  wire[3:0] T1086;
  reg [3:0] counts_172;
  wire[3:0] T10517;
  wire[3:0] T1087;
  wire[3:0] T1088;
  wire T1089;
  wire T1090;
  reg [3:0] counts_173;
  wire[3:0] T10518;
  wire[3:0] T1091;
  wire[3:0] T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire[3:0] T1096;
  reg [3:0] counts_174;
  wire[3:0] T10519;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire T1099;
  wire T1100;
  reg [3:0] counts_175;
  wire[3:0] T10520;
  wire[3:0] T1101;
  wire[3:0] T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire[3:0] T1109;
  wire[3:0] T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  reg [3:0] counts_176;
  wire[3:0] T10521;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire T1115;
  wire T1116;
  reg [3:0] counts_177;
  wire[3:0] T10522;
  wire[3:0] T1117;
  wire[3:0] T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire[3:0] T1122;
  reg [3:0] counts_178;
  wire[3:0] T10523;
  wire[3:0] T1123;
  wire[3:0] T1124;
  wire T1125;
  wire T1126;
  reg [3:0] counts_179;
  wire[3:0] T10524;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire[3:0] T1133;
  wire[3:0] T1134;
  reg [3:0] counts_180;
  wire[3:0] T10525;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire T1137;
  wire T1138;
  reg [3:0] counts_181;
  wire[3:0] T10526;
  wire[3:0] T1139;
  wire[3:0] T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[3:0] T1144;
  reg [3:0] counts_182;
  wire[3:0] T10527;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire T1147;
  wire T1148;
  reg [3:0] counts_183;
  wire[3:0] T10528;
  wire[3:0] T1149;
  wire[3:0] T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire[3:0] T1156;
  wire[3:0] T1157;
  wire[3:0] T1158;
  reg [3:0] counts_184;
  wire[3:0] T10529;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire T1161;
  wire T1162;
  reg [3:0] counts_185;
  wire[3:0] T10530;
  wire[3:0] T1163;
  wire[3:0] T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire[3:0] T1168;
  reg [3:0] counts_186;
  wire[3:0] T10531;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire T1171;
  wire T1172;
  reg [3:0] counts_187;
  wire[3:0] T10532;
  wire[3:0] T1173;
  wire[3:0] T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire[3:0] T1179;
  wire[3:0] T1180;
  reg [3:0] counts_188;
  wire[3:0] T10533;
  wire[3:0] T1181;
  wire[3:0] T1182;
  wire T1183;
  wire T1184;
  reg [3:0] counts_189;
  wire[3:0] T10534;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire[3:0] T1190;
  reg [3:0] counts_190;
  wire[3:0] T10535;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire T1193;
  wire T1194;
  reg [3:0] counts_191;
  wire[3:0] T10536;
  wire[3:0] T1195;
  wire[3:0] T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire[3:0] T1205;
  wire[3:0] T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  reg [3:0] counts_192;
  wire[3:0] T10537;
  wire[3:0] T1211;
  wire[3:0] T1212;
  wire T1213;
  wire T1214;
  reg [3:0] counts_193;
  wire[3:0] T10538;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire[3:0] T1220;
  reg [3:0] counts_194;
  wire[3:0] T10539;
  wire[3:0] T1221;
  wire[3:0] T1222;
  wire T1223;
  wire T1224;
  reg [3:0] counts_195;
  wire[3:0] T10540;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  reg [3:0] counts_196;
  wire[3:0] T10541;
  wire[3:0] T1233;
  wire[3:0] T1234;
  wire T1235;
  wire T1236;
  reg [3:0] counts_197;
  wire[3:0] T10542;
  wire[3:0] T1237;
  wire[3:0] T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire[3:0] T1242;
  reg [3:0] counts_198;
  wire[3:0] T10543;
  wire[3:0] T1243;
  wire[3:0] T1244;
  wire T1245;
  wire T1246;
  reg [3:0] counts_199;
  wire[3:0] T10544;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire[3:0] T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  reg [3:0] counts_200;
  wire[3:0] T10545;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire T1259;
  wire T1260;
  reg [3:0] counts_201;
  wire[3:0] T10546;
  wire[3:0] T1261;
  wire[3:0] T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire[3:0] T1266;
  reg [3:0] counts_202;
  wire[3:0] T10547;
  wire[3:0] T1267;
  wire[3:0] T1268;
  wire T1269;
  wire T1270;
  reg [3:0] counts_203;
  wire[3:0] T10548;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire[3:0] T1277;
  wire[3:0] T1278;
  reg [3:0] counts_204;
  wire[3:0] T10549;
  wire[3:0] T1279;
  wire[3:0] T1280;
  wire T1281;
  wire T1282;
  reg [3:0] counts_205;
  wire[3:0] T10550;
  wire[3:0] T1283;
  wire[3:0] T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire[3:0] T1288;
  reg [3:0] counts_206;
  wire[3:0] T10551;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire T1291;
  wire T1292;
  reg [3:0] counts_207;
  wire[3:0] T10552;
  wire[3:0] T1293;
  wire[3:0] T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire[3:0] T1301;
  wire[3:0] T1302;
  wire[3:0] T1303;
  wire[3:0] T1304;
  reg [3:0] counts_208;
  wire[3:0] T10553;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire T1307;
  wire T1308;
  reg [3:0] counts_209;
  wire[3:0] T10554;
  wire[3:0] T1309;
  wire[3:0] T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire[3:0] T1314;
  reg [3:0] counts_210;
  wire[3:0] T10555;
  wire[3:0] T1315;
  wire[3:0] T1316;
  wire T1317;
  wire T1318;
  reg [3:0] counts_211;
  wire[3:0] T10556;
  wire[3:0] T1319;
  wire[3:0] T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire[3:0] T1325;
  wire[3:0] T1326;
  reg [3:0] counts_212;
  wire[3:0] T10557;
  wire[3:0] T1327;
  wire[3:0] T1328;
  wire T1329;
  wire T1330;
  reg [3:0] counts_213;
  wire[3:0] T10558;
  wire[3:0] T1331;
  wire[3:0] T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  wire[3:0] T1336;
  reg [3:0] counts_214;
  wire[3:0] T10559;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire T1339;
  wire T1340;
  reg [3:0] counts_215;
  wire[3:0] T10560;
  wire[3:0] T1341;
  wire[3:0] T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[3:0] T1348;
  wire[3:0] T1349;
  wire[3:0] T1350;
  reg [3:0] counts_216;
  wire[3:0] T10561;
  wire[3:0] T1351;
  wire[3:0] T1352;
  wire T1353;
  wire T1354;
  reg [3:0] counts_217;
  wire[3:0] T10562;
  wire[3:0] T1355;
  wire[3:0] T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire[3:0] T1360;
  reg [3:0] counts_218;
  wire[3:0] T10563;
  wire[3:0] T1361;
  wire[3:0] T1362;
  wire T1363;
  wire T1364;
  reg [3:0] counts_219;
  wire[3:0] T10564;
  wire[3:0] T1365;
  wire[3:0] T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire[3:0] T1371;
  wire[3:0] T1372;
  reg [3:0] counts_220;
  wire[3:0] T10565;
  wire[3:0] T1373;
  wire[3:0] T1374;
  wire T1375;
  wire T1376;
  reg [3:0] counts_221;
  wire[3:0] T10566;
  wire[3:0] T1377;
  wire[3:0] T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire[3:0] T1382;
  reg [3:0] counts_222;
  wire[3:0] T10567;
  wire[3:0] T1383;
  wire[3:0] T1384;
  wire T1385;
  wire T1386;
  reg [3:0] counts_223;
  wire[3:0] T10568;
  wire[3:0] T1387;
  wire[3:0] T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[3:0] T1396;
  wire[3:0] T1397;
  wire[3:0] T1398;
  wire[3:0] T1399;
  wire[3:0] T1400;
  reg [3:0] counts_224;
  wire[3:0] T10569;
  wire[3:0] T1401;
  wire[3:0] T1402;
  wire T1403;
  wire T1404;
  reg [3:0] counts_225;
  wire[3:0] T10570;
  wire[3:0] T1405;
  wire[3:0] T1406;
  wire T1407;
  wire T1408;
  wire T1409;
  wire[3:0] T1410;
  reg [3:0] counts_226;
  wire[3:0] T10571;
  wire[3:0] T1411;
  wire[3:0] T1412;
  wire T1413;
  wire T1414;
  reg [3:0] counts_227;
  wire[3:0] T10572;
  wire[3:0] T1415;
  wire[3:0] T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire[3:0] T1421;
  wire[3:0] T1422;
  reg [3:0] counts_228;
  wire[3:0] T10573;
  wire[3:0] T1423;
  wire[3:0] T1424;
  wire T1425;
  wire T1426;
  reg [3:0] counts_229;
  wire[3:0] T10574;
  wire[3:0] T1427;
  wire[3:0] T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[3:0] T1432;
  reg [3:0] counts_230;
  wire[3:0] T10575;
  wire[3:0] T1433;
  wire[3:0] T1434;
  wire T1435;
  wire T1436;
  reg [3:0] counts_231;
  wire[3:0] T10576;
  wire[3:0] T1437;
  wire[3:0] T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire T1442;
  wire T1443;
  wire[3:0] T1444;
  wire[3:0] T1445;
  wire[3:0] T1446;
  reg [3:0] counts_232;
  wire[3:0] T10577;
  wire[3:0] T1447;
  wire[3:0] T1448;
  wire T1449;
  wire T1450;
  reg [3:0] counts_233;
  wire[3:0] T10578;
  wire[3:0] T1451;
  wire[3:0] T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire[3:0] T1456;
  reg [3:0] counts_234;
  wire[3:0] T10579;
  wire[3:0] T1457;
  wire[3:0] T1458;
  wire T1459;
  wire T1460;
  reg [3:0] counts_235;
  wire[3:0] T10580;
  wire[3:0] T1461;
  wire[3:0] T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire[3:0] T1467;
  wire[3:0] T1468;
  reg [3:0] counts_236;
  wire[3:0] T10581;
  wire[3:0] T1469;
  wire[3:0] T1470;
  wire T1471;
  wire T1472;
  reg [3:0] counts_237;
  wire[3:0] T10582;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire T1475;
  wire T1476;
  wire T1477;
  wire[3:0] T1478;
  reg [3:0] counts_238;
  wire[3:0] T10583;
  wire[3:0] T1479;
  wire[3:0] T1480;
  wire T1481;
  wire T1482;
  reg [3:0] counts_239;
  wire[3:0] T10584;
  wire[3:0] T1483;
  wire[3:0] T1484;
  wire T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire[3:0] T1491;
  wire[3:0] T1492;
  wire[3:0] T1493;
  wire[3:0] T1494;
  reg [3:0] counts_240;
  wire[3:0] T10585;
  wire[3:0] T1495;
  wire[3:0] T1496;
  wire T1497;
  wire T1498;
  reg [3:0] counts_241;
  wire[3:0] T10586;
  wire[3:0] T1499;
  wire[3:0] T1500;
  wire T1501;
  wire T1502;
  wire T1503;
  wire[3:0] T1504;
  reg [3:0] counts_242;
  wire[3:0] T10587;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire T1507;
  wire T1508;
  reg [3:0] counts_243;
  wire[3:0] T10588;
  wire[3:0] T1509;
  wire[3:0] T1510;
  wire T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire[3:0] T1515;
  wire[3:0] T1516;
  reg [3:0] counts_244;
  wire[3:0] T10589;
  wire[3:0] T1517;
  wire[3:0] T1518;
  wire T1519;
  wire T1520;
  reg [3:0] counts_245;
  wire[3:0] T10590;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire T1523;
  wire T1524;
  wire T1525;
  wire[3:0] T1526;
  reg [3:0] counts_246;
  wire[3:0] T10591;
  wire[3:0] T1527;
  wire[3:0] T1528;
  wire T1529;
  wire T1530;
  reg [3:0] counts_247;
  wire[3:0] T10592;
  wire[3:0] T1531;
  wire[3:0] T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[3:0] T1540;
  reg [3:0] counts_248;
  wire[3:0] T10593;
  wire[3:0] T1541;
  wire[3:0] T1542;
  wire T1543;
  wire T1544;
  reg [3:0] counts_249;
  wire[3:0] T10594;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire T1547;
  wire T1548;
  wire T1549;
  wire[3:0] T1550;
  reg [3:0] counts_250;
  wire[3:0] T10595;
  wire[3:0] T1551;
  wire[3:0] T1552;
  wire T1553;
  wire T1554;
  reg [3:0] counts_251;
  wire[3:0] T10596;
  wire[3:0] T1555;
  wire[3:0] T1556;
  wire T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  reg [3:0] counts_252;
  wire[3:0] T10597;
  wire[3:0] T1563;
  wire[3:0] T1564;
  wire T1565;
  wire T1566;
  reg [3:0] counts_253;
  wire[3:0] T10598;
  wire[3:0] T1567;
  wire[3:0] T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire[3:0] T1572;
  reg [3:0] counts_254;
  wire[3:0] T10599;
  wire[3:0] T1573;
  wire[3:0] T1574;
  wire T1575;
  wire T1576;
  reg [3:0] counts_255;
  wire[3:0] T10600;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire T1579;
  wire T1580;
  wire T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire T1585;
  wire T1586;
  wire T1587;
  wire T1588;
  wire[3:0] T1589;
  wire[3:0] T1590;
  wire[3:0] T1591;
  wire[3:0] T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[3:0] T1596;
  reg [3:0] counts_256;
  wire[3:0] T10601;
  wire[3:0] T1597;
  wire[3:0] T1598;
  wire T1599;
  wire T1600;
  reg [3:0] counts_257;
  wire[3:0] T10602;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire T1603;
  wire T1604;
  wire T1605;
  wire[3:0] T1606;
  reg [3:0] counts_258;
  wire[3:0] T10603;
  wire[3:0] T1607;
  wire[3:0] T1608;
  wire T1609;
  wire T1610;
  reg [3:0] counts_259;
  wire[3:0] T10604;
  wire[3:0] T1611;
  wire[3:0] T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  reg [3:0] counts_260;
  wire[3:0] T10605;
  wire[3:0] T1619;
  wire[3:0] T1620;
  wire T1621;
  wire T1622;
  reg [3:0] counts_261;
  wire[3:0] T10606;
  wire[3:0] T1623;
  wire[3:0] T1624;
  wire T1625;
  wire T1626;
  wire T1627;
  wire[3:0] T1628;
  reg [3:0] counts_262;
  wire[3:0] T10607;
  wire[3:0] T1629;
  wire[3:0] T1630;
  wire T1631;
  wire T1632;
  reg [3:0] counts_263;
  wire[3:0] T10608;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire T1635;
  wire T1636;
  wire T1637;
  wire T1638;
  wire T1639;
  wire[3:0] T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  reg [3:0] counts_264;
  wire[3:0] T10609;
  wire[3:0] T1643;
  wire[3:0] T1644;
  wire T1645;
  wire T1646;
  reg [3:0] counts_265;
  wire[3:0] T10610;
  wire[3:0] T1647;
  wire[3:0] T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire[3:0] T1652;
  reg [3:0] counts_266;
  wire[3:0] T10611;
  wire[3:0] T1653;
  wire[3:0] T1654;
  wire T1655;
  wire T1656;
  reg [3:0] counts_267;
  wire[3:0] T10612;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire T1659;
  wire T1660;
  wire T1661;
  wire T1662;
  wire[3:0] T1663;
  wire[3:0] T1664;
  reg [3:0] counts_268;
  wire[3:0] T10613;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire T1667;
  wire T1668;
  reg [3:0] counts_269;
  wire[3:0] T10614;
  wire[3:0] T1669;
  wire[3:0] T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire[3:0] T1674;
  reg [3:0] counts_270;
  wire[3:0] T10615;
  wire[3:0] T1675;
  wire[3:0] T1676;
  wire T1677;
  wire T1678;
  reg [3:0] counts_271;
  wire[3:0] T10616;
  wire[3:0] T1679;
  wire[3:0] T1680;
  wire T1681;
  wire T1682;
  wire T1683;
  wire T1684;
  wire T1685;
  wire T1686;
  wire[3:0] T1687;
  wire[3:0] T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  reg [3:0] counts_272;
  wire[3:0] T10617;
  wire[3:0] T1691;
  wire[3:0] T1692;
  wire T1693;
  wire T1694;
  reg [3:0] counts_273;
  wire[3:0] T10618;
  wire[3:0] T1695;
  wire[3:0] T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire[3:0] T1700;
  reg [3:0] counts_274;
  wire[3:0] T10619;
  wire[3:0] T1701;
  wire[3:0] T1702;
  wire T1703;
  wire T1704;
  reg [3:0] counts_275;
  wire[3:0] T10620;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire T1707;
  wire T1708;
  wire T1709;
  wire T1710;
  wire[3:0] T1711;
  wire[3:0] T1712;
  reg [3:0] counts_276;
  wire[3:0] T10621;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire T1715;
  wire T1716;
  reg [3:0] counts_277;
  wire[3:0] T10622;
  wire[3:0] T1717;
  wire[3:0] T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire[3:0] T1722;
  reg [3:0] counts_278;
  wire[3:0] T10623;
  wire[3:0] T1723;
  wire[3:0] T1724;
  wire T1725;
  wire T1726;
  reg [3:0] counts_279;
  wire[3:0] T10624;
  wire[3:0] T1727;
  wire[3:0] T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire T1732;
  wire T1733;
  wire[3:0] T1734;
  wire[3:0] T1735;
  wire[3:0] T1736;
  reg [3:0] counts_280;
  wire[3:0] T10625;
  wire[3:0] T1737;
  wire[3:0] T1738;
  wire T1739;
  wire T1740;
  reg [3:0] counts_281;
  wire[3:0] T10626;
  wire[3:0] T1741;
  wire[3:0] T1742;
  wire T1743;
  wire T1744;
  wire T1745;
  wire[3:0] T1746;
  reg [3:0] counts_282;
  wire[3:0] T10627;
  wire[3:0] T1747;
  wire[3:0] T1748;
  wire T1749;
  wire T1750;
  reg [3:0] counts_283;
  wire[3:0] T10628;
  wire[3:0] T1751;
  wire[3:0] T1752;
  wire T1753;
  wire T1754;
  wire T1755;
  wire T1756;
  wire[3:0] T1757;
  wire[3:0] T1758;
  reg [3:0] counts_284;
  wire[3:0] T10629;
  wire[3:0] T1759;
  wire[3:0] T1760;
  wire T1761;
  wire T1762;
  reg [3:0] counts_285;
  wire[3:0] T10630;
  wire[3:0] T1763;
  wire[3:0] T1764;
  wire T1765;
  wire T1766;
  wire T1767;
  wire[3:0] T1768;
  reg [3:0] counts_286;
  wire[3:0] T10631;
  wire[3:0] T1769;
  wire[3:0] T1770;
  wire T1771;
  wire T1772;
  reg [3:0] counts_287;
  wire[3:0] T10632;
  wire[3:0] T1773;
  wire[3:0] T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire T1778;
  wire T1779;
  wire T1780;
  wire T1781;
  wire[3:0] T1782;
  wire[3:0] T1783;
  wire[3:0] T1784;
  wire[3:0] T1785;
  wire[3:0] T1786;
  reg [3:0] counts_288;
  wire[3:0] T10633;
  wire[3:0] T1787;
  wire[3:0] T1788;
  wire T1789;
  wire T1790;
  reg [3:0] counts_289;
  wire[3:0] T10634;
  wire[3:0] T1791;
  wire[3:0] T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire[3:0] T1796;
  reg [3:0] counts_290;
  wire[3:0] T10635;
  wire[3:0] T1797;
  wire[3:0] T1798;
  wire T1799;
  wire T1800;
  reg [3:0] counts_291;
  wire[3:0] T10636;
  wire[3:0] T1801;
  wire[3:0] T1802;
  wire T1803;
  wire T1804;
  wire T1805;
  wire T1806;
  wire[3:0] T1807;
  wire[3:0] T1808;
  reg [3:0] counts_292;
  wire[3:0] T10637;
  wire[3:0] T1809;
  wire[3:0] T1810;
  wire T1811;
  wire T1812;
  reg [3:0] counts_293;
  wire[3:0] T10638;
  wire[3:0] T1813;
  wire[3:0] T1814;
  wire T1815;
  wire T1816;
  wire T1817;
  wire[3:0] T1818;
  reg [3:0] counts_294;
  wire[3:0] T10639;
  wire[3:0] T1819;
  wire[3:0] T1820;
  wire T1821;
  wire T1822;
  reg [3:0] counts_295;
  wire[3:0] T10640;
  wire[3:0] T1823;
  wire[3:0] T1824;
  wire T1825;
  wire T1826;
  wire T1827;
  wire T1828;
  wire T1829;
  wire[3:0] T1830;
  wire[3:0] T1831;
  wire[3:0] T1832;
  reg [3:0] counts_296;
  wire[3:0] T10641;
  wire[3:0] T1833;
  wire[3:0] T1834;
  wire T1835;
  wire T1836;
  reg [3:0] counts_297;
  wire[3:0] T10642;
  wire[3:0] T1837;
  wire[3:0] T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire[3:0] T1842;
  reg [3:0] counts_298;
  wire[3:0] T10643;
  wire[3:0] T1843;
  wire[3:0] T1844;
  wire T1845;
  wire T1846;
  reg [3:0] counts_299;
  wire[3:0] T10644;
  wire[3:0] T1847;
  wire[3:0] T1848;
  wire T1849;
  wire T1850;
  wire T1851;
  wire T1852;
  wire[3:0] T1853;
  wire[3:0] T1854;
  reg [3:0] counts_300;
  wire[3:0] T10645;
  wire[3:0] T1855;
  wire[3:0] T1856;
  wire T1857;
  wire T1858;
  reg [3:0] counts_301;
  wire[3:0] T10646;
  wire[3:0] T1859;
  wire[3:0] T1860;
  wire T1861;
  wire T1862;
  wire T1863;
  wire[3:0] T1864;
  reg [3:0] counts_302;
  wire[3:0] T10647;
  wire[3:0] T1865;
  wire[3:0] T1866;
  wire T1867;
  wire T1868;
  reg [3:0] counts_303;
  wire[3:0] T10648;
  wire[3:0] T1869;
  wire[3:0] T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire T1876;
  wire[3:0] T1877;
  wire[3:0] T1878;
  wire[3:0] T1879;
  wire[3:0] T1880;
  reg [3:0] counts_304;
  wire[3:0] T10649;
  wire[3:0] T1881;
  wire[3:0] T1882;
  wire T1883;
  wire T1884;
  reg [3:0] counts_305;
  wire[3:0] T10650;
  wire[3:0] T1885;
  wire[3:0] T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire[3:0] T1890;
  reg [3:0] counts_306;
  wire[3:0] T10651;
  wire[3:0] T1891;
  wire[3:0] T1892;
  wire T1893;
  wire T1894;
  reg [3:0] counts_307;
  wire[3:0] T10652;
  wire[3:0] T1895;
  wire[3:0] T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire T1900;
  wire[3:0] T1901;
  wire[3:0] T1902;
  reg [3:0] counts_308;
  wire[3:0] T10653;
  wire[3:0] T1903;
  wire[3:0] T1904;
  wire T1905;
  wire T1906;
  reg [3:0] counts_309;
  wire[3:0] T10654;
  wire[3:0] T1907;
  wire[3:0] T1908;
  wire T1909;
  wire T1910;
  wire T1911;
  wire[3:0] T1912;
  reg [3:0] counts_310;
  wire[3:0] T10655;
  wire[3:0] T1913;
  wire[3:0] T1914;
  wire T1915;
  wire T1916;
  reg [3:0] counts_311;
  wire[3:0] T10656;
  wire[3:0] T1917;
  wire[3:0] T1918;
  wire T1919;
  wire T1920;
  wire T1921;
  wire T1922;
  wire T1923;
  wire[3:0] T1924;
  wire[3:0] T1925;
  wire[3:0] T1926;
  reg [3:0] counts_312;
  wire[3:0] T10657;
  wire[3:0] T1927;
  wire[3:0] T1928;
  wire T1929;
  wire T1930;
  reg [3:0] counts_313;
  wire[3:0] T10658;
  wire[3:0] T1931;
  wire[3:0] T1932;
  wire T1933;
  wire T1934;
  wire T1935;
  wire[3:0] T1936;
  reg [3:0] counts_314;
  wire[3:0] T10659;
  wire[3:0] T1937;
  wire[3:0] T1938;
  wire T1939;
  wire T1940;
  reg [3:0] counts_315;
  wire[3:0] T10660;
  wire[3:0] T1941;
  wire[3:0] T1942;
  wire T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire[3:0] T1947;
  wire[3:0] T1948;
  reg [3:0] counts_316;
  wire[3:0] T10661;
  wire[3:0] T1949;
  wire[3:0] T1950;
  wire T1951;
  wire T1952;
  reg [3:0] counts_317;
  wire[3:0] T10662;
  wire[3:0] T1953;
  wire[3:0] T1954;
  wire T1955;
  wire T1956;
  wire T1957;
  wire[3:0] T1958;
  reg [3:0] counts_318;
  wire[3:0] T10663;
  wire[3:0] T1959;
  wire[3:0] T1960;
  wire T1961;
  wire T1962;
  reg [3:0] counts_319;
  wire[3:0] T10664;
  wire[3:0] T1963;
  wire[3:0] T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire T1972;
  wire[3:0] T1973;
  wire[3:0] T1974;
  wire[3:0] T1975;
  wire[3:0] T1976;
  wire[3:0] T1977;
  wire[3:0] T1978;
  reg [3:0] counts_320;
  wire[3:0] T10665;
  wire[3:0] T1979;
  wire[3:0] T1980;
  wire T1981;
  wire T1982;
  reg [3:0] counts_321;
  wire[3:0] T10666;
  wire[3:0] T1983;
  wire[3:0] T1984;
  wire T1985;
  wire T1986;
  wire T1987;
  wire[3:0] T1988;
  reg [3:0] counts_322;
  wire[3:0] T10667;
  wire[3:0] T1989;
  wire[3:0] T1990;
  wire T1991;
  wire T1992;
  reg [3:0] counts_323;
  wire[3:0] T10668;
  wire[3:0] T1993;
  wire[3:0] T1994;
  wire T1995;
  wire T1996;
  wire T1997;
  wire T1998;
  wire[3:0] T1999;
  wire[3:0] T2000;
  reg [3:0] counts_324;
  wire[3:0] T10669;
  wire[3:0] T2001;
  wire[3:0] T2002;
  wire T2003;
  wire T2004;
  reg [3:0] counts_325;
  wire[3:0] T10670;
  wire[3:0] T2005;
  wire[3:0] T2006;
  wire T2007;
  wire T2008;
  wire T2009;
  wire[3:0] T2010;
  reg [3:0] counts_326;
  wire[3:0] T10671;
  wire[3:0] T2011;
  wire[3:0] T2012;
  wire T2013;
  wire T2014;
  reg [3:0] counts_327;
  wire[3:0] T10672;
  wire[3:0] T2015;
  wire[3:0] T2016;
  wire T2017;
  wire T2018;
  wire T2019;
  wire T2020;
  wire T2021;
  wire[3:0] T2022;
  wire[3:0] T2023;
  wire[3:0] T2024;
  reg [3:0] counts_328;
  wire[3:0] T10673;
  wire[3:0] T2025;
  wire[3:0] T2026;
  wire T2027;
  wire T2028;
  reg [3:0] counts_329;
  wire[3:0] T10674;
  wire[3:0] T2029;
  wire[3:0] T2030;
  wire T2031;
  wire T2032;
  wire T2033;
  wire[3:0] T2034;
  reg [3:0] counts_330;
  wire[3:0] T10675;
  wire[3:0] T2035;
  wire[3:0] T2036;
  wire T2037;
  wire T2038;
  reg [3:0] counts_331;
  wire[3:0] T10676;
  wire[3:0] T2039;
  wire[3:0] T2040;
  wire T2041;
  wire T2042;
  wire T2043;
  wire T2044;
  wire[3:0] T2045;
  wire[3:0] T2046;
  reg [3:0] counts_332;
  wire[3:0] T10677;
  wire[3:0] T2047;
  wire[3:0] T2048;
  wire T2049;
  wire T2050;
  reg [3:0] counts_333;
  wire[3:0] T10678;
  wire[3:0] T2051;
  wire[3:0] T2052;
  wire T2053;
  wire T2054;
  wire T2055;
  wire[3:0] T2056;
  reg [3:0] counts_334;
  wire[3:0] T10679;
  wire[3:0] T2057;
  wire[3:0] T2058;
  wire T2059;
  wire T2060;
  reg [3:0] counts_335;
  wire[3:0] T10680;
  wire[3:0] T2061;
  wire[3:0] T2062;
  wire T2063;
  wire T2064;
  wire T2065;
  wire T2066;
  wire T2067;
  wire T2068;
  wire[3:0] T2069;
  wire[3:0] T2070;
  wire[3:0] T2071;
  wire[3:0] T2072;
  reg [3:0] counts_336;
  wire[3:0] T10681;
  wire[3:0] T2073;
  wire[3:0] T2074;
  wire T2075;
  wire T2076;
  reg [3:0] counts_337;
  wire[3:0] T10682;
  wire[3:0] T2077;
  wire[3:0] T2078;
  wire T2079;
  wire T2080;
  wire T2081;
  wire[3:0] T2082;
  reg [3:0] counts_338;
  wire[3:0] T10683;
  wire[3:0] T2083;
  wire[3:0] T2084;
  wire T2085;
  wire T2086;
  reg [3:0] counts_339;
  wire[3:0] T10684;
  wire[3:0] T2087;
  wire[3:0] T2088;
  wire T2089;
  wire T2090;
  wire T2091;
  wire T2092;
  wire[3:0] T2093;
  wire[3:0] T2094;
  reg [3:0] counts_340;
  wire[3:0] T10685;
  wire[3:0] T2095;
  wire[3:0] T2096;
  wire T2097;
  wire T2098;
  reg [3:0] counts_341;
  wire[3:0] T10686;
  wire[3:0] T2099;
  wire[3:0] T2100;
  wire T2101;
  wire T2102;
  wire T2103;
  wire[3:0] T2104;
  reg [3:0] counts_342;
  wire[3:0] T10687;
  wire[3:0] T2105;
  wire[3:0] T2106;
  wire T2107;
  wire T2108;
  reg [3:0] counts_343;
  wire[3:0] T10688;
  wire[3:0] T2109;
  wire[3:0] T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire T2115;
  wire[3:0] T2116;
  wire[3:0] T2117;
  wire[3:0] T2118;
  reg [3:0] counts_344;
  wire[3:0] T10689;
  wire[3:0] T2119;
  wire[3:0] T2120;
  wire T2121;
  wire T2122;
  reg [3:0] counts_345;
  wire[3:0] T10690;
  wire[3:0] T2123;
  wire[3:0] T2124;
  wire T2125;
  wire T2126;
  wire T2127;
  wire[3:0] T2128;
  reg [3:0] counts_346;
  wire[3:0] T10691;
  wire[3:0] T2129;
  wire[3:0] T2130;
  wire T2131;
  wire T2132;
  reg [3:0] counts_347;
  wire[3:0] T10692;
  wire[3:0] T2133;
  wire[3:0] T2134;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire[3:0] T2139;
  wire[3:0] T2140;
  reg [3:0] counts_348;
  wire[3:0] T10693;
  wire[3:0] T2141;
  wire[3:0] T2142;
  wire T2143;
  wire T2144;
  reg [3:0] counts_349;
  wire[3:0] T10694;
  wire[3:0] T2145;
  wire[3:0] T2146;
  wire T2147;
  wire T2148;
  wire T2149;
  wire[3:0] T2150;
  reg [3:0] counts_350;
  wire[3:0] T10695;
  wire[3:0] T2151;
  wire[3:0] T2152;
  wire T2153;
  wire T2154;
  reg [3:0] counts_351;
  wire[3:0] T10696;
  wire[3:0] T2155;
  wire[3:0] T2156;
  wire T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire[3:0] T2164;
  wire[3:0] T2165;
  wire[3:0] T2166;
  wire[3:0] T2167;
  wire[3:0] T2168;
  reg [3:0] counts_352;
  wire[3:0] T10697;
  wire[3:0] T2169;
  wire[3:0] T2170;
  wire T2171;
  wire T2172;
  reg [3:0] counts_353;
  wire[3:0] T10698;
  wire[3:0] T2173;
  wire[3:0] T2174;
  wire T2175;
  wire T2176;
  wire T2177;
  wire[3:0] T2178;
  reg [3:0] counts_354;
  wire[3:0] T10699;
  wire[3:0] T2179;
  wire[3:0] T2180;
  wire T2181;
  wire T2182;
  reg [3:0] counts_355;
  wire[3:0] T10700;
  wire[3:0] T2183;
  wire[3:0] T2184;
  wire T2185;
  wire T2186;
  wire T2187;
  wire T2188;
  wire[3:0] T2189;
  wire[3:0] T2190;
  reg [3:0] counts_356;
  wire[3:0] T10701;
  wire[3:0] T2191;
  wire[3:0] T2192;
  wire T2193;
  wire T2194;
  reg [3:0] counts_357;
  wire[3:0] T10702;
  wire[3:0] T2195;
  wire[3:0] T2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire[3:0] T2200;
  reg [3:0] counts_358;
  wire[3:0] T10703;
  wire[3:0] T2201;
  wire[3:0] T2202;
  wire T2203;
  wire T2204;
  reg [3:0] counts_359;
  wire[3:0] T10704;
  wire[3:0] T2205;
  wire[3:0] T2206;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  wire T2211;
  wire[3:0] T2212;
  wire[3:0] T2213;
  wire[3:0] T2214;
  reg [3:0] counts_360;
  wire[3:0] T10705;
  wire[3:0] T2215;
  wire[3:0] T2216;
  wire T2217;
  wire T2218;
  reg [3:0] counts_361;
  wire[3:0] T10706;
  wire[3:0] T2219;
  wire[3:0] T2220;
  wire T2221;
  wire T2222;
  wire T2223;
  wire[3:0] T2224;
  reg [3:0] counts_362;
  wire[3:0] T10707;
  wire[3:0] T2225;
  wire[3:0] T2226;
  wire T2227;
  wire T2228;
  reg [3:0] counts_363;
  wire[3:0] T10708;
  wire[3:0] T2229;
  wire[3:0] T2230;
  wire T2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire[3:0] T2235;
  wire[3:0] T2236;
  reg [3:0] counts_364;
  wire[3:0] T10709;
  wire[3:0] T2237;
  wire[3:0] T2238;
  wire T2239;
  wire T2240;
  reg [3:0] counts_365;
  wire[3:0] T10710;
  wire[3:0] T2241;
  wire[3:0] T2242;
  wire T2243;
  wire T2244;
  wire T2245;
  wire[3:0] T2246;
  reg [3:0] counts_366;
  wire[3:0] T10711;
  wire[3:0] T2247;
  wire[3:0] T2248;
  wire T2249;
  wire T2250;
  reg [3:0] counts_367;
  wire[3:0] T10712;
  wire[3:0] T2251;
  wire[3:0] T2252;
  wire T2253;
  wire T2254;
  wire T2255;
  wire T2256;
  wire T2257;
  wire T2258;
  wire[3:0] T2259;
  wire[3:0] T2260;
  wire[3:0] T2261;
  wire[3:0] T2262;
  reg [3:0] counts_368;
  wire[3:0] T10713;
  wire[3:0] T2263;
  wire[3:0] T2264;
  wire T2265;
  wire T2266;
  reg [3:0] counts_369;
  wire[3:0] T10714;
  wire[3:0] T2267;
  wire[3:0] T2268;
  wire T2269;
  wire T2270;
  wire T2271;
  wire[3:0] T2272;
  reg [3:0] counts_370;
  wire[3:0] T10715;
  wire[3:0] T2273;
  wire[3:0] T2274;
  wire T2275;
  wire T2276;
  reg [3:0] counts_371;
  wire[3:0] T10716;
  wire[3:0] T2277;
  wire[3:0] T2278;
  wire T2279;
  wire T2280;
  wire T2281;
  wire T2282;
  wire[3:0] T2283;
  wire[3:0] T2284;
  reg [3:0] counts_372;
  wire[3:0] T10717;
  wire[3:0] T2285;
  wire[3:0] T2286;
  wire T2287;
  wire T2288;
  reg [3:0] counts_373;
  wire[3:0] T10718;
  wire[3:0] T2289;
  wire[3:0] T2290;
  wire T2291;
  wire T2292;
  wire T2293;
  wire[3:0] T2294;
  reg [3:0] counts_374;
  wire[3:0] T10719;
  wire[3:0] T2295;
  wire[3:0] T2296;
  wire T2297;
  wire T2298;
  reg [3:0] counts_375;
  wire[3:0] T10720;
  wire[3:0] T2299;
  wire[3:0] T2300;
  wire T2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire T2305;
  wire[3:0] T2306;
  wire[3:0] T2307;
  wire[3:0] T2308;
  reg [3:0] counts_376;
  wire[3:0] T10721;
  wire[3:0] T2309;
  wire[3:0] T2310;
  wire T2311;
  wire T2312;
  reg [3:0] counts_377;
  wire[3:0] T10722;
  wire[3:0] T2313;
  wire[3:0] T2314;
  wire T2315;
  wire T2316;
  wire T2317;
  wire[3:0] T2318;
  reg [3:0] counts_378;
  wire[3:0] T10723;
  wire[3:0] T2319;
  wire[3:0] T2320;
  wire T2321;
  wire T2322;
  reg [3:0] counts_379;
  wire[3:0] T10724;
  wire[3:0] T2323;
  wire[3:0] T2324;
  wire T2325;
  wire T2326;
  wire T2327;
  wire T2328;
  wire[3:0] T2329;
  wire[3:0] T2330;
  reg [3:0] counts_380;
  wire[3:0] T10725;
  wire[3:0] T2331;
  wire[3:0] T2332;
  wire T2333;
  wire T2334;
  reg [3:0] counts_381;
  wire[3:0] T10726;
  wire[3:0] T2335;
  wire[3:0] T2336;
  wire T2337;
  wire T2338;
  wire T2339;
  wire[3:0] T2340;
  reg [3:0] counts_382;
  wire[3:0] T10727;
  wire[3:0] T2341;
  wire[3:0] T2342;
  wire T2343;
  wire T2344;
  reg [3:0] counts_383;
  wire[3:0] T10728;
  wire[3:0] T2345;
  wire[3:0] T2346;
  wire T2347;
  wire T2348;
  wire T2349;
  wire T2350;
  wire T2351;
  wire T2352;
  wire T2353;
  wire T2354;
  wire T2355;
  wire[3:0] T2356;
  wire[3:0] T2357;
  wire[3:0] T2358;
  wire[3:0] T2359;
  wire[3:0] T2360;
  wire[3:0] T2361;
  wire[3:0] T2362;
  reg [3:0] counts_384;
  wire[3:0] T10729;
  wire[3:0] T2363;
  wire[3:0] T2364;
  wire T2365;
  wire T2366;
  reg [3:0] counts_385;
  wire[3:0] T10730;
  wire[3:0] T2367;
  wire[3:0] T2368;
  wire T2369;
  wire T2370;
  wire T2371;
  wire[3:0] T2372;
  reg [3:0] counts_386;
  wire[3:0] T10731;
  wire[3:0] T2373;
  wire[3:0] T2374;
  wire T2375;
  wire T2376;
  reg [3:0] counts_387;
  wire[3:0] T10732;
  wire[3:0] T2377;
  wire[3:0] T2378;
  wire T2379;
  wire T2380;
  wire T2381;
  wire T2382;
  wire[3:0] T2383;
  wire[3:0] T2384;
  reg [3:0] counts_388;
  wire[3:0] T10733;
  wire[3:0] T2385;
  wire[3:0] T2386;
  wire T2387;
  wire T2388;
  reg [3:0] counts_389;
  wire[3:0] T10734;
  wire[3:0] T2389;
  wire[3:0] T2390;
  wire T2391;
  wire T2392;
  wire T2393;
  wire[3:0] T2394;
  reg [3:0] counts_390;
  wire[3:0] T10735;
  wire[3:0] T2395;
  wire[3:0] T2396;
  wire T2397;
  wire T2398;
  reg [3:0] counts_391;
  wire[3:0] T10736;
  wire[3:0] T2399;
  wire[3:0] T2400;
  wire T2401;
  wire T2402;
  wire T2403;
  wire T2404;
  wire T2405;
  wire[3:0] T2406;
  wire[3:0] T2407;
  wire[3:0] T2408;
  reg [3:0] counts_392;
  wire[3:0] T10737;
  wire[3:0] T2409;
  wire[3:0] T2410;
  wire T2411;
  wire T2412;
  reg [3:0] counts_393;
  wire[3:0] T10738;
  wire[3:0] T2413;
  wire[3:0] T2414;
  wire T2415;
  wire T2416;
  wire T2417;
  wire[3:0] T2418;
  reg [3:0] counts_394;
  wire[3:0] T10739;
  wire[3:0] T2419;
  wire[3:0] T2420;
  wire T2421;
  wire T2422;
  reg [3:0] counts_395;
  wire[3:0] T10740;
  wire[3:0] T2423;
  wire[3:0] T2424;
  wire T2425;
  wire T2426;
  wire T2427;
  wire T2428;
  wire[3:0] T2429;
  wire[3:0] T2430;
  reg [3:0] counts_396;
  wire[3:0] T10741;
  wire[3:0] T2431;
  wire[3:0] T2432;
  wire T2433;
  wire T2434;
  reg [3:0] counts_397;
  wire[3:0] T10742;
  wire[3:0] T2435;
  wire[3:0] T2436;
  wire T2437;
  wire T2438;
  wire T2439;
  wire[3:0] T2440;
  reg [3:0] counts_398;
  wire[3:0] T10743;
  wire[3:0] T2441;
  wire[3:0] T2442;
  wire T2443;
  wire T2444;
  reg [3:0] counts_399;
  wire[3:0] T10744;
  wire[3:0] T2445;
  wire[3:0] T2446;
  wire T2447;
  wire T2448;
  wire T2449;
  wire T2450;
  wire T2451;
  wire T2452;
  wire[3:0] T2453;
  wire[3:0] T2454;
  wire[3:0] T2455;
  wire[3:0] T2456;
  reg [3:0] counts_400;
  wire[3:0] T10745;
  wire[3:0] T2457;
  wire[3:0] T2458;
  wire T2459;
  wire T2460;
  reg [3:0] counts_401;
  wire[3:0] T10746;
  wire[3:0] T2461;
  wire[3:0] T2462;
  wire T2463;
  wire T2464;
  wire T2465;
  wire[3:0] T2466;
  reg [3:0] counts_402;
  wire[3:0] T10747;
  wire[3:0] T2467;
  wire[3:0] T2468;
  wire T2469;
  wire T2470;
  reg [3:0] counts_403;
  wire[3:0] T10748;
  wire[3:0] T2471;
  wire[3:0] T2472;
  wire T2473;
  wire T2474;
  wire T2475;
  wire T2476;
  wire[3:0] T2477;
  wire[3:0] T2478;
  reg [3:0] counts_404;
  wire[3:0] T10749;
  wire[3:0] T2479;
  wire[3:0] T2480;
  wire T2481;
  wire T2482;
  reg [3:0] counts_405;
  wire[3:0] T10750;
  wire[3:0] T2483;
  wire[3:0] T2484;
  wire T2485;
  wire T2486;
  wire T2487;
  wire[3:0] T2488;
  reg [3:0] counts_406;
  wire[3:0] T10751;
  wire[3:0] T2489;
  wire[3:0] T2490;
  wire T2491;
  wire T2492;
  reg [3:0] counts_407;
  wire[3:0] T10752;
  wire[3:0] T2493;
  wire[3:0] T2494;
  wire T2495;
  wire T2496;
  wire T2497;
  wire T2498;
  wire T2499;
  wire[3:0] T2500;
  wire[3:0] T2501;
  wire[3:0] T2502;
  reg [3:0] counts_408;
  wire[3:0] T10753;
  wire[3:0] T2503;
  wire[3:0] T2504;
  wire T2505;
  wire T2506;
  reg [3:0] counts_409;
  wire[3:0] T10754;
  wire[3:0] T2507;
  wire[3:0] T2508;
  wire T2509;
  wire T2510;
  wire T2511;
  wire[3:0] T2512;
  reg [3:0] counts_410;
  wire[3:0] T10755;
  wire[3:0] T2513;
  wire[3:0] T2514;
  wire T2515;
  wire T2516;
  reg [3:0] counts_411;
  wire[3:0] T10756;
  wire[3:0] T2517;
  wire[3:0] T2518;
  wire T2519;
  wire T2520;
  wire T2521;
  wire T2522;
  wire[3:0] T2523;
  wire[3:0] T2524;
  reg [3:0] counts_412;
  wire[3:0] T10757;
  wire[3:0] T2525;
  wire[3:0] T2526;
  wire T2527;
  wire T2528;
  reg [3:0] counts_413;
  wire[3:0] T10758;
  wire[3:0] T2529;
  wire[3:0] T2530;
  wire T2531;
  wire T2532;
  wire T2533;
  wire[3:0] T2534;
  reg [3:0] counts_414;
  wire[3:0] T10759;
  wire[3:0] T2535;
  wire[3:0] T2536;
  wire T2537;
  wire T2538;
  reg [3:0] counts_415;
  wire[3:0] T10760;
  wire[3:0] T2539;
  wire[3:0] T2540;
  wire T2541;
  wire T2542;
  wire T2543;
  wire T2544;
  wire T2545;
  wire T2546;
  wire T2547;
  wire[3:0] T2548;
  wire[3:0] T2549;
  wire[3:0] T2550;
  wire[3:0] T2551;
  wire[3:0] T2552;
  reg [3:0] counts_416;
  wire[3:0] T10761;
  wire[3:0] T2553;
  wire[3:0] T2554;
  wire T2555;
  wire T2556;
  reg [3:0] counts_417;
  wire[3:0] T10762;
  wire[3:0] T2557;
  wire[3:0] T2558;
  wire T2559;
  wire T2560;
  wire T2561;
  wire[3:0] T2562;
  reg [3:0] counts_418;
  wire[3:0] T10763;
  wire[3:0] T2563;
  wire[3:0] T2564;
  wire T2565;
  wire T2566;
  reg [3:0] counts_419;
  wire[3:0] T10764;
  wire[3:0] T2567;
  wire[3:0] T2568;
  wire T2569;
  wire T2570;
  wire T2571;
  wire T2572;
  wire[3:0] T2573;
  wire[3:0] T2574;
  reg [3:0] counts_420;
  wire[3:0] T10765;
  wire[3:0] T2575;
  wire[3:0] T2576;
  wire T2577;
  wire T2578;
  reg [3:0] counts_421;
  wire[3:0] T10766;
  wire[3:0] T2579;
  wire[3:0] T2580;
  wire T2581;
  wire T2582;
  wire T2583;
  wire[3:0] T2584;
  reg [3:0] counts_422;
  wire[3:0] T10767;
  wire[3:0] T2585;
  wire[3:0] T2586;
  wire T2587;
  wire T2588;
  reg [3:0] counts_423;
  wire[3:0] T10768;
  wire[3:0] T2589;
  wire[3:0] T2590;
  wire T2591;
  wire T2592;
  wire T2593;
  wire T2594;
  wire T2595;
  wire[3:0] T2596;
  wire[3:0] T2597;
  wire[3:0] T2598;
  reg [3:0] counts_424;
  wire[3:0] T10769;
  wire[3:0] T2599;
  wire[3:0] T2600;
  wire T2601;
  wire T2602;
  reg [3:0] counts_425;
  wire[3:0] T10770;
  wire[3:0] T2603;
  wire[3:0] T2604;
  wire T2605;
  wire T2606;
  wire T2607;
  wire[3:0] T2608;
  reg [3:0] counts_426;
  wire[3:0] T10771;
  wire[3:0] T2609;
  wire[3:0] T2610;
  wire T2611;
  wire T2612;
  reg [3:0] counts_427;
  wire[3:0] T10772;
  wire[3:0] T2613;
  wire[3:0] T2614;
  wire T2615;
  wire T2616;
  wire T2617;
  wire T2618;
  wire[3:0] T2619;
  wire[3:0] T2620;
  reg [3:0] counts_428;
  wire[3:0] T10773;
  wire[3:0] T2621;
  wire[3:0] T2622;
  wire T2623;
  wire T2624;
  reg [3:0] counts_429;
  wire[3:0] T10774;
  wire[3:0] T2625;
  wire[3:0] T2626;
  wire T2627;
  wire T2628;
  wire T2629;
  wire[3:0] T2630;
  reg [3:0] counts_430;
  wire[3:0] T10775;
  wire[3:0] T2631;
  wire[3:0] T2632;
  wire T2633;
  wire T2634;
  reg [3:0] counts_431;
  wire[3:0] T10776;
  wire[3:0] T2635;
  wire[3:0] T2636;
  wire T2637;
  wire T2638;
  wire T2639;
  wire T2640;
  wire T2641;
  wire T2642;
  wire[3:0] T2643;
  wire[3:0] T2644;
  wire[3:0] T2645;
  wire[3:0] T2646;
  reg [3:0] counts_432;
  wire[3:0] T10777;
  wire[3:0] T2647;
  wire[3:0] T2648;
  wire T2649;
  wire T2650;
  reg [3:0] counts_433;
  wire[3:0] T10778;
  wire[3:0] T2651;
  wire[3:0] T2652;
  wire T2653;
  wire T2654;
  wire T2655;
  wire[3:0] T2656;
  reg [3:0] counts_434;
  wire[3:0] T10779;
  wire[3:0] T2657;
  wire[3:0] T2658;
  wire T2659;
  wire T2660;
  reg [3:0] counts_435;
  wire[3:0] T10780;
  wire[3:0] T2661;
  wire[3:0] T2662;
  wire T2663;
  wire T2664;
  wire T2665;
  wire T2666;
  wire[3:0] T2667;
  wire[3:0] T2668;
  reg [3:0] counts_436;
  wire[3:0] T10781;
  wire[3:0] T2669;
  wire[3:0] T2670;
  wire T2671;
  wire T2672;
  reg [3:0] counts_437;
  wire[3:0] T10782;
  wire[3:0] T2673;
  wire[3:0] T2674;
  wire T2675;
  wire T2676;
  wire T2677;
  wire[3:0] T2678;
  reg [3:0] counts_438;
  wire[3:0] T10783;
  wire[3:0] T2679;
  wire[3:0] T2680;
  wire T2681;
  wire T2682;
  reg [3:0] counts_439;
  wire[3:0] T10784;
  wire[3:0] T2683;
  wire[3:0] T2684;
  wire T2685;
  wire T2686;
  wire T2687;
  wire T2688;
  wire T2689;
  wire[3:0] T2690;
  wire[3:0] T2691;
  wire[3:0] T2692;
  reg [3:0] counts_440;
  wire[3:0] T10785;
  wire[3:0] T2693;
  wire[3:0] T2694;
  wire T2695;
  wire T2696;
  reg [3:0] counts_441;
  wire[3:0] T10786;
  wire[3:0] T2697;
  wire[3:0] T2698;
  wire T2699;
  wire T2700;
  wire T2701;
  wire[3:0] T2702;
  reg [3:0] counts_442;
  wire[3:0] T10787;
  wire[3:0] T2703;
  wire[3:0] T2704;
  wire T2705;
  wire T2706;
  reg [3:0] counts_443;
  wire[3:0] T10788;
  wire[3:0] T2707;
  wire[3:0] T2708;
  wire T2709;
  wire T2710;
  wire T2711;
  wire T2712;
  wire[3:0] T2713;
  wire[3:0] T2714;
  reg [3:0] counts_444;
  wire[3:0] T10789;
  wire[3:0] T2715;
  wire[3:0] T2716;
  wire T2717;
  wire T2718;
  reg [3:0] counts_445;
  wire[3:0] T10790;
  wire[3:0] T2719;
  wire[3:0] T2720;
  wire T2721;
  wire T2722;
  wire T2723;
  wire[3:0] T2724;
  reg [3:0] counts_446;
  wire[3:0] T10791;
  wire[3:0] T2725;
  wire[3:0] T2726;
  wire T2727;
  wire T2728;
  reg [3:0] counts_447;
  wire[3:0] T10792;
  wire[3:0] T2729;
  wire[3:0] T2730;
  wire T2731;
  wire T2732;
  wire T2733;
  wire T2734;
  wire T2735;
  wire T2736;
  wire T2737;
  wire T2738;
  wire[3:0] T2739;
  wire[3:0] T2740;
  wire[3:0] T2741;
  wire[3:0] T2742;
  wire[3:0] T2743;
  wire[3:0] T2744;
  reg [3:0] counts_448;
  wire[3:0] T10793;
  wire[3:0] T2745;
  wire[3:0] T2746;
  wire T2747;
  wire T2748;
  reg [3:0] counts_449;
  wire[3:0] T10794;
  wire[3:0] T2749;
  wire[3:0] T2750;
  wire T2751;
  wire T2752;
  wire T2753;
  wire[3:0] T2754;
  reg [3:0] counts_450;
  wire[3:0] T10795;
  wire[3:0] T2755;
  wire[3:0] T2756;
  wire T2757;
  wire T2758;
  reg [3:0] counts_451;
  wire[3:0] T10796;
  wire[3:0] T2759;
  wire[3:0] T2760;
  wire T2761;
  wire T2762;
  wire T2763;
  wire T2764;
  wire[3:0] T2765;
  wire[3:0] T2766;
  reg [3:0] counts_452;
  wire[3:0] T10797;
  wire[3:0] T2767;
  wire[3:0] T2768;
  wire T2769;
  wire T2770;
  reg [3:0] counts_453;
  wire[3:0] T10798;
  wire[3:0] T2771;
  wire[3:0] T2772;
  wire T2773;
  wire T2774;
  wire T2775;
  wire[3:0] T2776;
  reg [3:0] counts_454;
  wire[3:0] T10799;
  wire[3:0] T2777;
  wire[3:0] T2778;
  wire T2779;
  wire T2780;
  reg [3:0] counts_455;
  wire[3:0] T10800;
  wire[3:0] T2781;
  wire[3:0] T2782;
  wire T2783;
  wire T2784;
  wire T2785;
  wire T2786;
  wire T2787;
  wire[3:0] T2788;
  wire[3:0] T2789;
  wire[3:0] T2790;
  reg [3:0] counts_456;
  wire[3:0] T10801;
  wire[3:0] T2791;
  wire[3:0] T2792;
  wire T2793;
  wire T2794;
  reg [3:0] counts_457;
  wire[3:0] T10802;
  wire[3:0] T2795;
  wire[3:0] T2796;
  wire T2797;
  wire T2798;
  wire T2799;
  wire[3:0] T2800;
  reg [3:0] counts_458;
  wire[3:0] T10803;
  wire[3:0] T2801;
  wire[3:0] T2802;
  wire T2803;
  wire T2804;
  reg [3:0] counts_459;
  wire[3:0] T10804;
  wire[3:0] T2805;
  wire[3:0] T2806;
  wire T2807;
  wire T2808;
  wire T2809;
  wire T2810;
  wire[3:0] T2811;
  wire[3:0] T2812;
  reg [3:0] counts_460;
  wire[3:0] T10805;
  wire[3:0] T2813;
  wire[3:0] T2814;
  wire T2815;
  wire T2816;
  reg [3:0] counts_461;
  wire[3:0] T10806;
  wire[3:0] T2817;
  wire[3:0] T2818;
  wire T2819;
  wire T2820;
  wire T2821;
  wire[3:0] T2822;
  reg [3:0] counts_462;
  wire[3:0] T10807;
  wire[3:0] T2823;
  wire[3:0] T2824;
  wire T2825;
  wire T2826;
  reg [3:0] counts_463;
  wire[3:0] T10808;
  wire[3:0] T2827;
  wire[3:0] T2828;
  wire T2829;
  wire T2830;
  wire T2831;
  wire T2832;
  wire T2833;
  wire T2834;
  wire[3:0] T2835;
  wire[3:0] T2836;
  wire[3:0] T2837;
  wire[3:0] T2838;
  reg [3:0] counts_464;
  wire[3:0] T10809;
  wire[3:0] T2839;
  wire[3:0] T2840;
  wire T2841;
  wire T2842;
  reg [3:0] counts_465;
  wire[3:0] T10810;
  wire[3:0] T2843;
  wire[3:0] T2844;
  wire T2845;
  wire T2846;
  wire T2847;
  wire[3:0] T2848;
  reg [3:0] counts_466;
  wire[3:0] T10811;
  wire[3:0] T2849;
  wire[3:0] T2850;
  wire T2851;
  wire T2852;
  reg [3:0] counts_467;
  wire[3:0] T10812;
  wire[3:0] T2853;
  wire[3:0] T2854;
  wire T2855;
  wire T2856;
  wire T2857;
  wire T2858;
  wire[3:0] T2859;
  wire[3:0] T2860;
  reg [3:0] counts_468;
  wire[3:0] T10813;
  wire[3:0] T2861;
  wire[3:0] T2862;
  wire T2863;
  wire T2864;
  reg [3:0] counts_469;
  wire[3:0] T10814;
  wire[3:0] T2865;
  wire[3:0] T2866;
  wire T2867;
  wire T2868;
  wire T2869;
  wire[3:0] T2870;
  reg [3:0] counts_470;
  wire[3:0] T10815;
  wire[3:0] T2871;
  wire[3:0] T2872;
  wire T2873;
  wire T2874;
  reg [3:0] counts_471;
  wire[3:0] T10816;
  wire[3:0] T2875;
  wire[3:0] T2876;
  wire T2877;
  wire T2878;
  wire T2879;
  wire T2880;
  wire T2881;
  wire[3:0] T2882;
  wire[3:0] T2883;
  wire[3:0] T2884;
  reg [3:0] counts_472;
  wire[3:0] T10817;
  wire[3:0] T2885;
  wire[3:0] T2886;
  wire T2887;
  wire T2888;
  reg [3:0] counts_473;
  wire[3:0] T10818;
  wire[3:0] T2889;
  wire[3:0] T2890;
  wire T2891;
  wire T2892;
  wire T2893;
  wire[3:0] T2894;
  reg [3:0] counts_474;
  wire[3:0] T10819;
  wire[3:0] T2895;
  wire[3:0] T2896;
  wire T2897;
  wire T2898;
  reg [3:0] counts_475;
  wire[3:0] T10820;
  wire[3:0] T2899;
  wire[3:0] T2900;
  wire T2901;
  wire T2902;
  wire T2903;
  wire T2904;
  wire[3:0] T2905;
  wire[3:0] T2906;
  reg [3:0] counts_476;
  wire[3:0] T10821;
  wire[3:0] T2907;
  wire[3:0] T2908;
  wire T2909;
  wire T2910;
  reg [3:0] counts_477;
  wire[3:0] T10822;
  wire[3:0] T2911;
  wire[3:0] T2912;
  wire T2913;
  wire T2914;
  wire T2915;
  wire[3:0] T2916;
  reg [3:0] counts_478;
  wire[3:0] T10823;
  wire[3:0] T2917;
  wire[3:0] T2918;
  wire T2919;
  wire T2920;
  reg [3:0] counts_479;
  wire[3:0] T10824;
  wire[3:0] T2921;
  wire[3:0] T2922;
  wire T2923;
  wire T2924;
  wire T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire T2929;
  wire[3:0] T2930;
  wire[3:0] T2931;
  wire[3:0] T2932;
  wire[3:0] T2933;
  wire[3:0] T2934;
  reg [3:0] counts_480;
  wire[3:0] T10825;
  wire[3:0] T2935;
  wire[3:0] T2936;
  wire T2937;
  wire T2938;
  reg [3:0] counts_481;
  wire[3:0] T10826;
  wire[3:0] T2939;
  wire[3:0] T2940;
  wire T2941;
  wire T2942;
  wire T2943;
  wire[3:0] T2944;
  reg [3:0] counts_482;
  wire[3:0] T10827;
  wire[3:0] T2945;
  wire[3:0] T2946;
  wire T2947;
  wire T2948;
  reg [3:0] counts_483;
  wire[3:0] T10828;
  wire[3:0] T2949;
  wire[3:0] T2950;
  wire T2951;
  wire T2952;
  wire T2953;
  wire T2954;
  wire[3:0] T2955;
  wire[3:0] T2956;
  reg [3:0] counts_484;
  wire[3:0] T10829;
  wire[3:0] T2957;
  wire[3:0] T2958;
  wire T2959;
  wire T2960;
  reg [3:0] counts_485;
  wire[3:0] T10830;
  wire[3:0] T2961;
  wire[3:0] T2962;
  wire T2963;
  wire T2964;
  wire T2965;
  wire[3:0] T2966;
  reg [3:0] counts_486;
  wire[3:0] T10831;
  wire[3:0] T2967;
  wire[3:0] T2968;
  wire T2969;
  wire T2970;
  reg [3:0] counts_487;
  wire[3:0] T10832;
  wire[3:0] T2971;
  wire[3:0] T2972;
  wire T2973;
  wire T2974;
  wire T2975;
  wire T2976;
  wire T2977;
  wire[3:0] T2978;
  wire[3:0] T2979;
  wire[3:0] T2980;
  reg [3:0] counts_488;
  wire[3:0] T10833;
  wire[3:0] T2981;
  wire[3:0] T2982;
  wire T2983;
  wire T2984;
  reg [3:0] counts_489;
  wire[3:0] T10834;
  wire[3:0] T2985;
  wire[3:0] T2986;
  wire T2987;
  wire T2988;
  wire T2989;
  wire[3:0] T2990;
  reg [3:0] counts_490;
  wire[3:0] T10835;
  wire[3:0] T2991;
  wire[3:0] T2992;
  wire T2993;
  wire T2994;
  reg [3:0] counts_491;
  wire[3:0] T10836;
  wire[3:0] T2995;
  wire[3:0] T2996;
  wire T2997;
  wire T2998;
  wire T2999;
  wire T3000;
  wire[3:0] T3001;
  wire[3:0] T3002;
  reg [3:0] counts_492;
  wire[3:0] T10837;
  wire[3:0] T3003;
  wire[3:0] T3004;
  wire T3005;
  wire T3006;
  reg [3:0] counts_493;
  wire[3:0] T10838;
  wire[3:0] T3007;
  wire[3:0] T3008;
  wire T3009;
  wire T3010;
  wire T3011;
  wire[3:0] T3012;
  reg [3:0] counts_494;
  wire[3:0] T10839;
  wire[3:0] T3013;
  wire[3:0] T3014;
  wire T3015;
  wire T3016;
  reg [3:0] counts_495;
  wire[3:0] T10840;
  wire[3:0] T3017;
  wire[3:0] T3018;
  wire T3019;
  wire T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  wire T3024;
  wire[3:0] T3025;
  wire[3:0] T3026;
  wire[3:0] T3027;
  wire[3:0] T3028;
  reg [3:0] counts_496;
  wire[3:0] T10841;
  wire[3:0] T3029;
  wire[3:0] T3030;
  wire T3031;
  wire T3032;
  reg [3:0] counts_497;
  wire[3:0] T10842;
  wire[3:0] T3033;
  wire[3:0] T3034;
  wire T3035;
  wire T3036;
  wire T3037;
  wire[3:0] T3038;
  reg [3:0] counts_498;
  wire[3:0] T10843;
  wire[3:0] T3039;
  wire[3:0] T3040;
  wire T3041;
  wire T3042;
  reg [3:0] counts_499;
  wire[3:0] T10844;
  wire[3:0] T3043;
  wire[3:0] T3044;
  wire T3045;
  wire T3046;
  wire T3047;
  wire T3048;
  wire[3:0] T3049;
  wire[3:0] T3050;
  reg [3:0] counts_500;
  wire[3:0] T10845;
  wire[3:0] T3051;
  wire[3:0] T3052;
  wire T3053;
  wire T3054;
  reg [3:0] counts_501;
  wire[3:0] T10846;
  wire[3:0] T3055;
  wire[3:0] T3056;
  wire T3057;
  wire T3058;
  wire T3059;
  wire[3:0] T3060;
  reg [3:0] counts_502;
  wire[3:0] T10847;
  wire[3:0] T3061;
  wire[3:0] T3062;
  wire T3063;
  wire T3064;
  reg [3:0] counts_503;
  wire[3:0] T10848;
  wire[3:0] T3065;
  wire[3:0] T3066;
  wire T3067;
  wire T3068;
  wire T3069;
  wire T3070;
  wire T3071;
  wire[3:0] T3072;
  wire[3:0] T3073;
  wire[3:0] T3074;
  reg [3:0] counts_504;
  wire[3:0] T10849;
  wire[3:0] T3075;
  wire[3:0] T3076;
  wire T3077;
  wire T3078;
  reg [3:0] counts_505;
  wire[3:0] T10850;
  wire[3:0] T3079;
  wire[3:0] T3080;
  wire T3081;
  wire T3082;
  wire T3083;
  wire[3:0] T3084;
  reg [3:0] counts_506;
  wire[3:0] T10851;
  wire[3:0] T3085;
  wire[3:0] T3086;
  wire T3087;
  wire T3088;
  reg [3:0] counts_507;
  wire[3:0] T10852;
  wire[3:0] T3089;
  wire[3:0] T3090;
  wire T3091;
  wire T3092;
  wire T3093;
  wire T3094;
  wire[3:0] T3095;
  wire[3:0] T3096;
  reg [3:0] counts_508;
  wire[3:0] T10853;
  wire[3:0] T3097;
  wire[3:0] T3098;
  wire T3099;
  wire T3100;
  reg [3:0] counts_509;
  wire[3:0] T10854;
  wire[3:0] T3101;
  wire[3:0] T3102;
  wire T3103;
  wire T3104;
  wire T3105;
  wire[3:0] T3106;
  reg [3:0] counts_510;
  wire[3:0] T10855;
  wire[3:0] T3107;
  wire[3:0] T3108;
  wire T3109;
  wire T3110;
  reg [3:0] counts_511;
  wire[3:0] T10856;
  wire[3:0] T3111;
  wire[3:0] T3112;
  wire T3113;
  wire T3114;
  wire T3115;
  wire T3116;
  wire T3117;
  wire T3118;
  wire T3119;
  wire T3120;
  wire T3121;
  wire T3122;
  wire T3123;
  wire[3:0] T3124;
  wire[3:0] T3125;
  wire[3:0] T3126;
  wire[3:0] T3127;
  wire[3:0] T3128;
  wire[3:0] T3129;
  wire[3:0] T3130;
  wire[3:0] T3131;
  wire[3:0] T3132;
  reg [3:0] counts_512;
  wire[3:0] T10857;
  wire[3:0] T3133;
  wire[3:0] T3134;
  wire T3135;
  wire T3136;
  reg [3:0] counts_513;
  wire[3:0] T10858;
  wire[3:0] T3137;
  wire[3:0] T3138;
  wire T3139;
  wire T3140;
  wire T3141;
  wire[3:0] T3142;
  reg [3:0] counts_514;
  wire[3:0] T10859;
  wire[3:0] T3143;
  wire[3:0] T3144;
  wire T3145;
  wire T3146;
  reg [3:0] counts_515;
  wire[3:0] T10860;
  wire[3:0] T3147;
  wire[3:0] T3148;
  wire T3149;
  wire T3150;
  wire T3151;
  wire T3152;
  wire[3:0] T3153;
  wire[3:0] T3154;
  reg [3:0] counts_516;
  wire[3:0] T10861;
  wire[3:0] T3155;
  wire[3:0] T3156;
  wire T3157;
  wire T3158;
  reg [3:0] counts_517;
  wire[3:0] T10862;
  wire[3:0] T3159;
  wire[3:0] T3160;
  wire T3161;
  wire T3162;
  wire T3163;
  wire[3:0] T3164;
  reg [3:0] counts_518;
  wire[3:0] T10863;
  wire[3:0] T3165;
  wire[3:0] T3166;
  wire T3167;
  wire T3168;
  reg [3:0] counts_519;
  wire[3:0] T10864;
  wire[3:0] T3169;
  wire[3:0] T3170;
  wire T3171;
  wire T3172;
  wire T3173;
  wire T3174;
  wire T3175;
  wire[3:0] T3176;
  wire[3:0] T3177;
  wire[3:0] T3178;
  reg [3:0] counts_520;
  wire[3:0] T10865;
  wire[3:0] T3179;
  wire[3:0] T3180;
  wire T3181;
  wire T3182;
  reg [3:0] counts_521;
  wire[3:0] T10866;
  wire[3:0] T3183;
  wire[3:0] T3184;
  wire T3185;
  wire T3186;
  wire T3187;
  wire[3:0] T3188;
  reg [3:0] counts_522;
  wire[3:0] T10867;
  wire[3:0] T3189;
  wire[3:0] T3190;
  wire T3191;
  wire T3192;
  reg [3:0] counts_523;
  wire[3:0] T10868;
  wire[3:0] T3193;
  wire[3:0] T3194;
  wire T3195;
  wire T3196;
  wire T3197;
  wire T3198;
  wire[3:0] T3199;
  wire[3:0] T3200;
  reg [3:0] counts_524;
  wire[3:0] T10869;
  wire[3:0] T3201;
  wire[3:0] T3202;
  wire T3203;
  wire T3204;
  reg [3:0] counts_525;
  wire[3:0] T10870;
  wire[3:0] T3205;
  wire[3:0] T3206;
  wire T3207;
  wire T3208;
  wire T3209;
  wire[3:0] T3210;
  reg [3:0] counts_526;
  wire[3:0] T10871;
  wire[3:0] T3211;
  wire[3:0] T3212;
  wire T3213;
  wire T3214;
  reg [3:0] counts_527;
  wire[3:0] T10872;
  wire[3:0] T3215;
  wire[3:0] T3216;
  wire T3217;
  wire T3218;
  wire T3219;
  wire T3220;
  wire T3221;
  wire T3222;
  wire[3:0] T3223;
  wire[3:0] T3224;
  wire[3:0] T3225;
  wire[3:0] T3226;
  reg [3:0] counts_528;
  wire[3:0] T10873;
  wire[3:0] T3227;
  wire[3:0] T3228;
  wire T3229;
  wire T3230;
  reg [3:0] counts_529;
  wire[3:0] T10874;
  wire[3:0] T3231;
  wire[3:0] T3232;
  wire T3233;
  wire T3234;
  wire T3235;
  wire[3:0] T3236;
  reg [3:0] counts_530;
  wire[3:0] T10875;
  wire[3:0] T3237;
  wire[3:0] T3238;
  wire T3239;
  wire T3240;
  reg [3:0] counts_531;
  wire[3:0] T10876;
  wire[3:0] T3241;
  wire[3:0] T3242;
  wire T3243;
  wire T3244;
  wire T3245;
  wire T3246;
  wire[3:0] T3247;
  wire[3:0] T3248;
  reg [3:0] counts_532;
  wire[3:0] T10877;
  wire[3:0] T3249;
  wire[3:0] T3250;
  wire T3251;
  wire T3252;
  reg [3:0] counts_533;
  wire[3:0] T10878;
  wire[3:0] T3253;
  wire[3:0] T3254;
  wire T3255;
  wire T3256;
  wire T3257;
  wire[3:0] T3258;
  reg [3:0] counts_534;
  wire[3:0] T10879;
  wire[3:0] T3259;
  wire[3:0] T3260;
  wire T3261;
  wire T3262;
  reg [3:0] counts_535;
  wire[3:0] T10880;
  wire[3:0] T3263;
  wire[3:0] T3264;
  wire T3265;
  wire T3266;
  wire T3267;
  wire T3268;
  wire T3269;
  wire[3:0] T3270;
  wire[3:0] T3271;
  wire[3:0] T3272;
  reg [3:0] counts_536;
  wire[3:0] T10881;
  wire[3:0] T3273;
  wire[3:0] T3274;
  wire T3275;
  wire T3276;
  reg [3:0] counts_537;
  wire[3:0] T10882;
  wire[3:0] T3277;
  wire[3:0] T3278;
  wire T3279;
  wire T3280;
  wire T3281;
  wire[3:0] T3282;
  reg [3:0] counts_538;
  wire[3:0] T10883;
  wire[3:0] T3283;
  wire[3:0] T3284;
  wire T3285;
  wire T3286;
  reg [3:0] counts_539;
  wire[3:0] T10884;
  wire[3:0] T3287;
  wire[3:0] T3288;
  wire T3289;
  wire T3290;
  wire T3291;
  wire T3292;
  wire[3:0] T3293;
  wire[3:0] T3294;
  reg [3:0] counts_540;
  wire[3:0] T10885;
  wire[3:0] T3295;
  wire[3:0] T3296;
  wire T3297;
  wire T3298;
  reg [3:0] counts_541;
  wire[3:0] T10886;
  wire[3:0] T3299;
  wire[3:0] T3300;
  wire T3301;
  wire T3302;
  wire T3303;
  wire[3:0] T3304;
  reg [3:0] counts_542;
  wire[3:0] T10887;
  wire[3:0] T3305;
  wire[3:0] T3306;
  wire T3307;
  wire T3308;
  reg [3:0] counts_543;
  wire[3:0] T10888;
  wire[3:0] T3309;
  wire[3:0] T3310;
  wire T3311;
  wire T3312;
  wire T3313;
  wire T3314;
  wire T3315;
  wire T3316;
  wire T3317;
  wire[3:0] T3318;
  wire[3:0] T3319;
  wire[3:0] T3320;
  wire[3:0] T3321;
  wire[3:0] T3322;
  reg [3:0] counts_544;
  wire[3:0] T10889;
  wire[3:0] T3323;
  wire[3:0] T3324;
  wire T3325;
  wire T3326;
  reg [3:0] counts_545;
  wire[3:0] T10890;
  wire[3:0] T3327;
  wire[3:0] T3328;
  wire T3329;
  wire T3330;
  wire T3331;
  wire[3:0] T3332;
  reg [3:0] counts_546;
  wire[3:0] T10891;
  wire[3:0] T3333;
  wire[3:0] T3334;
  wire T3335;
  wire T3336;
  reg [3:0] counts_547;
  wire[3:0] T10892;
  wire[3:0] T3337;
  wire[3:0] T3338;
  wire T3339;
  wire T3340;
  wire T3341;
  wire T3342;
  wire[3:0] T3343;
  wire[3:0] T3344;
  reg [3:0] counts_548;
  wire[3:0] T10893;
  wire[3:0] T3345;
  wire[3:0] T3346;
  wire T3347;
  wire T3348;
  reg [3:0] counts_549;
  wire[3:0] T10894;
  wire[3:0] T3349;
  wire[3:0] T3350;
  wire T3351;
  wire T3352;
  wire T3353;
  wire[3:0] T3354;
  reg [3:0] counts_550;
  wire[3:0] T10895;
  wire[3:0] T3355;
  wire[3:0] T3356;
  wire T3357;
  wire T3358;
  reg [3:0] counts_551;
  wire[3:0] T10896;
  wire[3:0] T3359;
  wire[3:0] T3360;
  wire T3361;
  wire T3362;
  wire T3363;
  wire T3364;
  wire T3365;
  wire[3:0] T3366;
  wire[3:0] T3367;
  wire[3:0] T3368;
  reg [3:0] counts_552;
  wire[3:0] T10897;
  wire[3:0] T3369;
  wire[3:0] T3370;
  wire T3371;
  wire T3372;
  reg [3:0] counts_553;
  wire[3:0] T10898;
  wire[3:0] T3373;
  wire[3:0] T3374;
  wire T3375;
  wire T3376;
  wire T3377;
  wire[3:0] T3378;
  reg [3:0] counts_554;
  wire[3:0] T10899;
  wire[3:0] T3379;
  wire[3:0] T3380;
  wire T3381;
  wire T3382;
  reg [3:0] counts_555;
  wire[3:0] T10900;
  wire[3:0] T3383;
  wire[3:0] T3384;
  wire T3385;
  wire T3386;
  wire T3387;
  wire T3388;
  wire[3:0] T3389;
  wire[3:0] T3390;
  reg [3:0] counts_556;
  wire[3:0] T10901;
  wire[3:0] T3391;
  wire[3:0] T3392;
  wire T3393;
  wire T3394;
  reg [3:0] counts_557;
  wire[3:0] T10902;
  wire[3:0] T3395;
  wire[3:0] T3396;
  wire T3397;
  wire T3398;
  wire T3399;
  wire[3:0] T3400;
  reg [3:0] counts_558;
  wire[3:0] T10903;
  wire[3:0] T3401;
  wire[3:0] T3402;
  wire T3403;
  wire T3404;
  reg [3:0] counts_559;
  wire[3:0] T10904;
  wire[3:0] T3405;
  wire[3:0] T3406;
  wire T3407;
  wire T3408;
  wire T3409;
  wire T3410;
  wire T3411;
  wire T3412;
  wire[3:0] T3413;
  wire[3:0] T3414;
  wire[3:0] T3415;
  wire[3:0] T3416;
  reg [3:0] counts_560;
  wire[3:0] T10905;
  wire[3:0] T3417;
  wire[3:0] T3418;
  wire T3419;
  wire T3420;
  reg [3:0] counts_561;
  wire[3:0] T10906;
  wire[3:0] T3421;
  wire[3:0] T3422;
  wire T3423;
  wire T3424;
  wire T3425;
  wire[3:0] T3426;
  reg [3:0] counts_562;
  wire[3:0] T10907;
  wire[3:0] T3427;
  wire[3:0] T3428;
  wire T3429;
  wire T3430;
  reg [3:0] counts_563;
  wire[3:0] T10908;
  wire[3:0] T3431;
  wire[3:0] T3432;
  wire T3433;
  wire T3434;
  wire T3435;
  wire T3436;
  wire[3:0] T3437;
  wire[3:0] T3438;
  reg [3:0] counts_564;
  wire[3:0] T10909;
  wire[3:0] T3439;
  wire[3:0] T3440;
  wire T3441;
  wire T3442;
  reg [3:0] counts_565;
  wire[3:0] T10910;
  wire[3:0] T3443;
  wire[3:0] T3444;
  wire T3445;
  wire T3446;
  wire T3447;
  wire[3:0] T3448;
  reg [3:0] counts_566;
  wire[3:0] T10911;
  wire[3:0] T3449;
  wire[3:0] T3450;
  wire T3451;
  wire T3452;
  reg [3:0] counts_567;
  wire[3:0] T10912;
  wire[3:0] T3453;
  wire[3:0] T3454;
  wire T3455;
  wire T3456;
  wire T3457;
  wire T3458;
  wire T3459;
  wire[3:0] T3460;
  wire[3:0] T3461;
  wire[3:0] T3462;
  reg [3:0] counts_568;
  wire[3:0] T10913;
  wire[3:0] T3463;
  wire[3:0] T3464;
  wire T3465;
  wire T3466;
  reg [3:0] counts_569;
  wire[3:0] T10914;
  wire[3:0] T3467;
  wire[3:0] T3468;
  wire T3469;
  wire T3470;
  wire T3471;
  wire[3:0] T3472;
  reg [3:0] counts_570;
  wire[3:0] T10915;
  wire[3:0] T3473;
  wire[3:0] T3474;
  wire T3475;
  wire T3476;
  reg [3:0] counts_571;
  wire[3:0] T10916;
  wire[3:0] T3477;
  wire[3:0] T3478;
  wire T3479;
  wire T3480;
  wire T3481;
  wire T3482;
  wire[3:0] T3483;
  wire[3:0] T3484;
  reg [3:0] counts_572;
  wire[3:0] T10917;
  wire[3:0] T3485;
  wire[3:0] T3486;
  wire T3487;
  wire T3488;
  reg [3:0] counts_573;
  wire[3:0] T10918;
  wire[3:0] T3489;
  wire[3:0] T3490;
  wire T3491;
  wire T3492;
  wire T3493;
  wire[3:0] T3494;
  reg [3:0] counts_574;
  wire[3:0] T10919;
  wire[3:0] T3495;
  wire[3:0] T3496;
  wire T3497;
  wire T3498;
  reg [3:0] counts_575;
  wire[3:0] T10920;
  wire[3:0] T3499;
  wire[3:0] T3500;
  wire T3501;
  wire T3502;
  wire T3503;
  wire T3504;
  wire T3505;
  wire T3506;
  wire T3507;
  wire T3508;
  wire[3:0] T3509;
  wire[3:0] T3510;
  wire[3:0] T3511;
  wire[3:0] T3512;
  wire[3:0] T3513;
  wire[3:0] T3514;
  reg [3:0] counts_576;
  wire[3:0] T10921;
  wire[3:0] T3515;
  wire[3:0] T3516;
  wire T3517;
  wire T3518;
  reg [3:0] counts_577;
  wire[3:0] T10922;
  wire[3:0] T3519;
  wire[3:0] T3520;
  wire T3521;
  wire T3522;
  wire T3523;
  wire[3:0] T3524;
  reg [3:0] counts_578;
  wire[3:0] T10923;
  wire[3:0] T3525;
  wire[3:0] T3526;
  wire T3527;
  wire T3528;
  reg [3:0] counts_579;
  wire[3:0] T10924;
  wire[3:0] T3529;
  wire[3:0] T3530;
  wire T3531;
  wire T3532;
  wire T3533;
  wire T3534;
  wire[3:0] T3535;
  wire[3:0] T3536;
  reg [3:0] counts_580;
  wire[3:0] T10925;
  wire[3:0] T3537;
  wire[3:0] T3538;
  wire T3539;
  wire T3540;
  reg [3:0] counts_581;
  wire[3:0] T10926;
  wire[3:0] T3541;
  wire[3:0] T3542;
  wire T3543;
  wire T3544;
  wire T3545;
  wire[3:0] T3546;
  reg [3:0] counts_582;
  wire[3:0] T10927;
  wire[3:0] T3547;
  wire[3:0] T3548;
  wire T3549;
  wire T3550;
  reg [3:0] counts_583;
  wire[3:0] T10928;
  wire[3:0] T3551;
  wire[3:0] T3552;
  wire T3553;
  wire T3554;
  wire T3555;
  wire T3556;
  wire T3557;
  wire[3:0] T3558;
  wire[3:0] T3559;
  wire[3:0] T3560;
  reg [3:0] counts_584;
  wire[3:0] T10929;
  wire[3:0] T3561;
  wire[3:0] T3562;
  wire T3563;
  wire T3564;
  reg [3:0] counts_585;
  wire[3:0] T10930;
  wire[3:0] T3565;
  wire[3:0] T3566;
  wire T3567;
  wire T3568;
  wire T3569;
  wire[3:0] T3570;
  reg [3:0] counts_586;
  wire[3:0] T10931;
  wire[3:0] T3571;
  wire[3:0] T3572;
  wire T3573;
  wire T3574;
  reg [3:0] counts_587;
  wire[3:0] T10932;
  wire[3:0] T3575;
  wire[3:0] T3576;
  wire T3577;
  wire T3578;
  wire T3579;
  wire T3580;
  wire[3:0] T3581;
  wire[3:0] T3582;
  reg [3:0] counts_588;
  wire[3:0] T10933;
  wire[3:0] T3583;
  wire[3:0] T3584;
  wire T3585;
  wire T3586;
  reg [3:0] counts_589;
  wire[3:0] T10934;
  wire[3:0] T3587;
  wire[3:0] T3588;
  wire T3589;
  wire T3590;
  wire T3591;
  wire[3:0] T3592;
  reg [3:0] counts_590;
  wire[3:0] T10935;
  wire[3:0] T3593;
  wire[3:0] T3594;
  wire T3595;
  wire T3596;
  reg [3:0] counts_591;
  wire[3:0] T10936;
  wire[3:0] T3597;
  wire[3:0] T3598;
  wire T3599;
  wire T3600;
  wire T3601;
  wire T3602;
  wire T3603;
  wire T3604;
  wire[3:0] T3605;
  wire[3:0] T3606;
  wire[3:0] T3607;
  wire[3:0] T3608;
  reg [3:0] counts_592;
  wire[3:0] T10937;
  wire[3:0] T3609;
  wire[3:0] T3610;
  wire T3611;
  wire T3612;
  reg [3:0] counts_593;
  wire[3:0] T10938;
  wire[3:0] T3613;
  wire[3:0] T3614;
  wire T3615;
  wire T3616;
  wire T3617;
  wire[3:0] T3618;
  reg [3:0] counts_594;
  wire[3:0] T10939;
  wire[3:0] T3619;
  wire[3:0] T3620;
  wire T3621;
  wire T3622;
  reg [3:0] counts_595;
  wire[3:0] T10940;
  wire[3:0] T3623;
  wire[3:0] T3624;
  wire T3625;
  wire T3626;
  wire T3627;
  wire T3628;
  wire[3:0] T3629;
  wire[3:0] T3630;
  reg [3:0] counts_596;
  wire[3:0] T10941;
  wire[3:0] T3631;
  wire[3:0] T3632;
  wire T3633;
  wire T3634;
  reg [3:0] counts_597;
  wire[3:0] T10942;
  wire[3:0] T3635;
  wire[3:0] T3636;
  wire T3637;
  wire T3638;
  wire T3639;
  wire[3:0] T3640;
  reg [3:0] counts_598;
  wire[3:0] T10943;
  wire[3:0] T3641;
  wire[3:0] T3642;
  wire T3643;
  wire T3644;
  reg [3:0] counts_599;
  wire[3:0] T10944;
  wire[3:0] T3645;
  wire[3:0] T3646;
  wire T3647;
  wire T3648;
  wire T3649;
  wire T3650;
  wire T3651;
  wire[3:0] T3652;
  wire[3:0] T3653;
  wire[3:0] T3654;
  reg [3:0] counts_600;
  wire[3:0] T10945;
  wire[3:0] T3655;
  wire[3:0] T3656;
  wire T3657;
  wire T3658;
  reg [3:0] counts_601;
  wire[3:0] T10946;
  wire[3:0] T3659;
  wire[3:0] T3660;
  wire T3661;
  wire T3662;
  wire T3663;
  wire[3:0] T3664;
  reg [3:0] counts_602;
  wire[3:0] T10947;
  wire[3:0] T3665;
  wire[3:0] T3666;
  wire T3667;
  wire T3668;
  reg [3:0] counts_603;
  wire[3:0] T10948;
  wire[3:0] T3669;
  wire[3:0] T3670;
  wire T3671;
  wire T3672;
  wire T3673;
  wire T3674;
  wire[3:0] T3675;
  wire[3:0] T3676;
  reg [3:0] counts_604;
  wire[3:0] T10949;
  wire[3:0] T3677;
  wire[3:0] T3678;
  wire T3679;
  wire T3680;
  reg [3:0] counts_605;
  wire[3:0] T10950;
  wire[3:0] T3681;
  wire[3:0] T3682;
  wire T3683;
  wire T3684;
  wire T3685;
  wire[3:0] T3686;
  reg [3:0] counts_606;
  wire[3:0] T10951;
  wire[3:0] T3687;
  wire[3:0] T3688;
  wire T3689;
  wire T3690;
  reg [3:0] counts_607;
  wire[3:0] T10952;
  wire[3:0] T3691;
  wire[3:0] T3692;
  wire T3693;
  wire T3694;
  wire T3695;
  wire T3696;
  wire T3697;
  wire T3698;
  wire T3699;
  wire[3:0] T3700;
  wire[3:0] T3701;
  wire[3:0] T3702;
  wire[3:0] T3703;
  wire[3:0] T3704;
  reg [3:0] counts_608;
  wire[3:0] T10953;
  wire[3:0] T3705;
  wire[3:0] T3706;
  wire T3707;
  wire T3708;
  reg [3:0] counts_609;
  wire[3:0] T10954;
  wire[3:0] T3709;
  wire[3:0] T3710;
  wire T3711;
  wire T3712;
  wire T3713;
  wire[3:0] T3714;
  reg [3:0] counts_610;
  wire[3:0] T10955;
  wire[3:0] T3715;
  wire[3:0] T3716;
  wire T3717;
  wire T3718;
  reg [3:0] counts_611;
  wire[3:0] T10956;
  wire[3:0] T3719;
  wire[3:0] T3720;
  wire T3721;
  wire T3722;
  wire T3723;
  wire T3724;
  wire[3:0] T3725;
  wire[3:0] T3726;
  reg [3:0] counts_612;
  wire[3:0] T10957;
  wire[3:0] T3727;
  wire[3:0] T3728;
  wire T3729;
  wire T3730;
  reg [3:0] counts_613;
  wire[3:0] T10958;
  wire[3:0] T3731;
  wire[3:0] T3732;
  wire T3733;
  wire T3734;
  wire T3735;
  wire[3:0] T3736;
  reg [3:0] counts_614;
  wire[3:0] T10959;
  wire[3:0] T3737;
  wire[3:0] T3738;
  wire T3739;
  wire T3740;
  reg [3:0] counts_615;
  wire[3:0] T10960;
  wire[3:0] T3741;
  wire[3:0] T3742;
  wire T3743;
  wire T3744;
  wire T3745;
  wire T3746;
  wire T3747;
  wire[3:0] T3748;
  wire[3:0] T3749;
  wire[3:0] T3750;
  reg [3:0] counts_616;
  wire[3:0] T10961;
  wire[3:0] T3751;
  wire[3:0] T3752;
  wire T3753;
  wire T3754;
  reg [3:0] counts_617;
  wire[3:0] T10962;
  wire[3:0] T3755;
  wire[3:0] T3756;
  wire T3757;
  wire T3758;
  wire T3759;
  wire[3:0] T3760;
  reg [3:0] counts_618;
  wire[3:0] T10963;
  wire[3:0] T3761;
  wire[3:0] T3762;
  wire T3763;
  wire T3764;
  reg [3:0] counts_619;
  wire[3:0] T10964;
  wire[3:0] T3765;
  wire[3:0] T3766;
  wire T3767;
  wire T3768;
  wire T3769;
  wire T3770;
  wire[3:0] T3771;
  wire[3:0] T3772;
  reg [3:0] counts_620;
  wire[3:0] T10965;
  wire[3:0] T3773;
  wire[3:0] T3774;
  wire T3775;
  wire T3776;
  reg [3:0] counts_621;
  wire[3:0] T10966;
  wire[3:0] T3777;
  wire[3:0] T3778;
  wire T3779;
  wire T3780;
  wire T3781;
  wire[3:0] T3782;
  reg [3:0] counts_622;
  wire[3:0] T10967;
  wire[3:0] T3783;
  wire[3:0] T3784;
  wire T3785;
  wire T3786;
  reg [3:0] counts_623;
  wire[3:0] T10968;
  wire[3:0] T3787;
  wire[3:0] T3788;
  wire T3789;
  wire T3790;
  wire T3791;
  wire T3792;
  wire T3793;
  wire T3794;
  wire[3:0] T3795;
  wire[3:0] T3796;
  wire[3:0] T3797;
  wire[3:0] T3798;
  reg [3:0] counts_624;
  wire[3:0] T10969;
  wire[3:0] T3799;
  wire[3:0] T3800;
  wire T3801;
  wire T3802;
  reg [3:0] counts_625;
  wire[3:0] T10970;
  wire[3:0] T3803;
  wire[3:0] T3804;
  wire T3805;
  wire T3806;
  wire T3807;
  wire[3:0] T3808;
  reg [3:0] counts_626;
  wire[3:0] T10971;
  wire[3:0] T3809;
  wire[3:0] T3810;
  wire T3811;
  wire T3812;
  reg [3:0] counts_627;
  wire[3:0] T10972;
  wire[3:0] T3813;
  wire[3:0] T3814;
  wire T3815;
  wire T3816;
  wire T3817;
  wire T3818;
  wire[3:0] T3819;
  wire[3:0] T3820;
  reg [3:0] counts_628;
  wire[3:0] T10973;
  wire[3:0] T3821;
  wire[3:0] T3822;
  wire T3823;
  wire T3824;
  reg [3:0] counts_629;
  wire[3:0] T10974;
  wire[3:0] T3825;
  wire[3:0] T3826;
  wire T3827;
  wire T3828;
  wire T3829;
  wire[3:0] T3830;
  reg [3:0] counts_630;
  wire[3:0] T10975;
  wire[3:0] T3831;
  wire[3:0] T3832;
  wire T3833;
  wire T3834;
  reg [3:0] counts_631;
  wire[3:0] T10976;
  wire[3:0] T3835;
  wire[3:0] T3836;
  wire T3837;
  wire T3838;
  wire T3839;
  wire T3840;
  wire T3841;
  wire[3:0] T3842;
  wire[3:0] T3843;
  wire[3:0] T3844;
  reg [3:0] counts_632;
  wire[3:0] T10977;
  wire[3:0] T3845;
  wire[3:0] T3846;
  wire T3847;
  wire T3848;
  reg [3:0] counts_633;
  wire[3:0] T10978;
  wire[3:0] T3849;
  wire[3:0] T3850;
  wire T3851;
  wire T3852;
  wire T3853;
  wire[3:0] T3854;
  reg [3:0] counts_634;
  wire[3:0] T10979;
  wire[3:0] T3855;
  wire[3:0] T3856;
  wire T3857;
  wire T3858;
  reg [3:0] counts_635;
  wire[3:0] T10980;
  wire[3:0] T3859;
  wire[3:0] T3860;
  wire T3861;
  wire T3862;
  wire T3863;
  wire T3864;
  wire[3:0] T3865;
  wire[3:0] T3866;
  reg [3:0] counts_636;
  wire[3:0] T10981;
  wire[3:0] T3867;
  wire[3:0] T3868;
  wire T3869;
  wire T3870;
  reg [3:0] counts_637;
  wire[3:0] T10982;
  wire[3:0] T3871;
  wire[3:0] T3872;
  wire T3873;
  wire T3874;
  wire T3875;
  wire[3:0] T3876;
  reg [3:0] counts_638;
  wire[3:0] T10983;
  wire[3:0] T3877;
  wire[3:0] T3878;
  wire T3879;
  wire T3880;
  reg [3:0] counts_639;
  wire[3:0] T10984;
  wire[3:0] T3881;
  wire[3:0] T3882;
  wire T3883;
  wire T3884;
  wire T3885;
  wire T3886;
  wire T3887;
  wire T3888;
  wire T3889;
  wire T3890;
  wire T3891;
  wire[3:0] T3892;
  wire[3:0] T3893;
  wire[3:0] T3894;
  wire[3:0] T3895;
  wire[3:0] T3896;
  wire[3:0] T3897;
  wire[3:0] T3898;
  reg [3:0] counts_640;
  wire[3:0] T10985;
  wire[3:0] T3899;
  wire[3:0] T3900;
  wire T3901;
  wire T3902;
  reg [3:0] counts_641;
  wire[3:0] T10986;
  wire[3:0] T3903;
  wire[3:0] T3904;
  wire T3905;
  wire T3906;
  wire T3907;
  wire[3:0] T3908;
  reg [3:0] counts_642;
  wire[3:0] T10987;
  wire[3:0] T3909;
  wire[3:0] T3910;
  wire T3911;
  wire T3912;
  reg [3:0] counts_643;
  wire[3:0] T10988;
  wire[3:0] T3913;
  wire[3:0] T3914;
  wire T3915;
  wire T3916;
  wire T3917;
  wire T3918;
  wire[3:0] T3919;
  wire[3:0] T3920;
  reg [3:0] counts_644;
  wire[3:0] T10989;
  wire[3:0] T3921;
  wire[3:0] T3922;
  wire T3923;
  wire T3924;
  reg [3:0] counts_645;
  wire[3:0] T10990;
  wire[3:0] T3925;
  wire[3:0] T3926;
  wire T3927;
  wire T3928;
  wire T3929;
  wire[3:0] T3930;
  reg [3:0] counts_646;
  wire[3:0] T10991;
  wire[3:0] T3931;
  wire[3:0] T3932;
  wire T3933;
  wire T3934;
  reg [3:0] counts_647;
  wire[3:0] T10992;
  wire[3:0] T3935;
  wire[3:0] T3936;
  wire T3937;
  wire T3938;
  wire T3939;
  wire T3940;
  wire T3941;
  wire[3:0] T3942;
  wire[3:0] T3943;
  wire[3:0] T3944;
  reg [3:0] counts_648;
  wire[3:0] T10993;
  wire[3:0] T3945;
  wire[3:0] T3946;
  wire T3947;
  wire T3948;
  reg [3:0] counts_649;
  wire[3:0] T10994;
  wire[3:0] T3949;
  wire[3:0] T3950;
  wire T3951;
  wire T3952;
  wire T3953;
  wire[3:0] T3954;
  reg [3:0] counts_650;
  wire[3:0] T10995;
  wire[3:0] T3955;
  wire[3:0] T3956;
  wire T3957;
  wire T3958;
  reg [3:0] counts_651;
  wire[3:0] T10996;
  wire[3:0] T3959;
  wire[3:0] T3960;
  wire T3961;
  wire T3962;
  wire T3963;
  wire T3964;
  wire[3:0] T3965;
  wire[3:0] T3966;
  reg [3:0] counts_652;
  wire[3:0] T10997;
  wire[3:0] T3967;
  wire[3:0] T3968;
  wire T3969;
  wire T3970;
  reg [3:0] counts_653;
  wire[3:0] T10998;
  wire[3:0] T3971;
  wire[3:0] T3972;
  wire T3973;
  wire T3974;
  wire T3975;
  wire[3:0] T3976;
  reg [3:0] counts_654;
  wire[3:0] T10999;
  wire[3:0] T3977;
  wire[3:0] T3978;
  wire T3979;
  wire T3980;
  reg [3:0] counts_655;
  wire[3:0] T11000;
  wire[3:0] T3981;
  wire[3:0] T3982;
  wire T3983;
  wire T3984;
  wire T3985;
  wire T3986;
  wire T3987;
  wire T3988;
  wire[3:0] T3989;
  wire[3:0] T3990;
  wire[3:0] T3991;
  wire[3:0] T3992;
  reg [3:0] counts_656;
  wire[3:0] T11001;
  wire[3:0] T3993;
  wire[3:0] T3994;
  wire T3995;
  wire T3996;
  reg [3:0] counts_657;
  wire[3:0] T11002;
  wire[3:0] T3997;
  wire[3:0] T3998;
  wire T3999;
  wire T4000;
  wire T4001;
  wire[3:0] T4002;
  reg [3:0] counts_658;
  wire[3:0] T11003;
  wire[3:0] T4003;
  wire[3:0] T4004;
  wire T4005;
  wire T4006;
  reg [3:0] counts_659;
  wire[3:0] T11004;
  wire[3:0] T4007;
  wire[3:0] T4008;
  wire T4009;
  wire T4010;
  wire T4011;
  wire T4012;
  wire[3:0] T4013;
  wire[3:0] T4014;
  reg [3:0] counts_660;
  wire[3:0] T11005;
  wire[3:0] T4015;
  wire[3:0] T4016;
  wire T4017;
  wire T4018;
  reg [3:0] counts_661;
  wire[3:0] T11006;
  wire[3:0] T4019;
  wire[3:0] T4020;
  wire T4021;
  wire T4022;
  wire T4023;
  wire[3:0] T4024;
  reg [3:0] counts_662;
  wire[3:0] T11007;
  wire[3:0] T4025;
  wire[3:0] T4026;
  wire T4027;
  wire T4028;
  reg [3:0] counts_663;
  wire[3:0] T11008;
  wire[3:0] T4029;
  wire[3:0] T4030;
  wire T4031;
  wire T4032;
  wire T4033;
  wire T4034;
  wire T4035;
  wire[3:0] T4036;
  wire[3:0] T4037;
  wire[3:0] T4038;
  reg [3:0] counts_664;
  wire[3:0] T11009;
  wire[3:0] T4039;
  wire[3:0] T4040;
  wire T4041;
  wire T4042;
  reg [3:0] counts_665;
  wire[3:0] T11010;
  wire[3:0] T4043;
  wire[3:0] T4044;
  wire T4045;
  wire T4046;
  wire T4047;
  wire[3:0] T4048;
  reg [3:0] counts_666;
  wire[3:0] T11011;
  wire[3:0] T4049;
  wire[3:0] T4050;
  wire T4051;
  wire T4052;
  reg [3:0] counts_667;
  wire[3:0] T11012;
  wire[3:0] T4053;
  wire[3:0] T4054;
  wire T4055;
  wire T4056;
  wire T4057;
  wire T4058;
  wire[3:0] T4059;
  wire[3:0] T4060;
  reg [3:0] counts_668;
  wire[3:0] T11013;
  wire[3:0] T4061;
  wire[3:0] T4062;
  wire T4063;
  wire T4064;
  reg [3:0] counts_669;
  wire[3:0] T11014;
  wire[3:0] T4065;
  wire[3:0] T4066;
  wire T4067;
  wire T4068;
  wire T4069;
  wire[3:0] T4070;
  reg [3:0] counts_670;
  wire[3:0] T11015;
  wire[3:0] T4071;
  wire[3:0] T4072;
  wire T4073;
  wire T4074;
  reg [3:0] counts_671;
  wire[3:0] T11016;
  wire[3:0] T4075;
  wire[3:0] T4076;
  wire T4077;
  wire T4078;
  wire T4079;
  wire T4080;
  wire T4081;
  wire T4082;
  wire T4083;
  wire[3:0] T4084;
  wire[3:0] T4085;
  wire[3:0] T4086;
  wire[3:0] T4087;
  wire[3:0] T4088;
  reg [3:0] counts_672;
  wire[3:0] T11017;
  wire[3:0] T4089;
  wire[3:0] T4090;
  wire T4091;
  wire T4092;
  reg [3:0] counts_673;
  wire[3:0] T11018;
  wire[3:0] T4093;
  wire[3:0] T4094;
  wire T4095;
  wire T4096;
  wire T4097;
  wire[3:0] T4098;
  reg [3:0] counts_674;
  wire[3:0] T11019;
  wire[3:0] T4099;
  wire[3:0] T4100;
  wire T4101;
  wire T4102;
  reg [3:0] counts_675;
  wire[3:0] T11020;
  wire[3:0] T4103;
  wire[3:0] T4104;
  wire T4105;
  wire T4106;
  wire T4107;
  wire T4108;
  wire[3:0] T4109;
  wire[3:0] T4110;
  reg [3:0] counts_676;
  wire[3:0] T11021;
  wire[3:0] T4111;
  wire[3:0] T4112;
  wire T4113;
  wire T4114;
  reg [3:0] counts_677;
  wire[3:0] T11022;
  wire[3:0] T4115;
  wire[3:0] T4116;
  wire T4117;
  wire T4118;
  wire T4119;
  wire[3:0] T4120;
  reg [3:0] counts_678;
  wire[3:0] T11023;
  wire[3:0] T4121;
  wire[3:0] T4122;
  wire T4123;
  wire T4124;
  reg [3:0] counts_679;
  wire[3:0] T11024;
  wire[3:0] T4125;
  wire[3:0] T4126;
  wire T4127;
  wire T4128;
  wire T4129;
  wire T4130;
  wire T4131;
  wire[3:0] T4132;
  wire[3:0] T4133;
  wire[3:0] T4134;
  reg [3:0] counts_680;
  wire[3:0] T11025;
  wire[3:0] T4135;
  wire[3:0] T4136;
  wire T4137;
  wire T4138;
  reg [3:0] counts_681;
  wire[3:0] T11026;
  wire[3:0] T4139;
  wire[3:0] T4140;
  wire T4141;
  wire T4142;
  wire T4143;
  wire[3:0] T4144;
  reg [3:0] counts_682;
  wire[3:0] T11027;
  wire[3:0] T4145;
  wire[3:0] T4146;
  wire T4147;
  wire T4148;
  reg [3:0] counts_683;
  wire[3:0] T11028;
  wire[3:0] T4149;
  wire[3:0] T4150;
  wire T4151;
  wire T4152;
  wire T4153;
  wire T4154;
  wire[3:0] T4155;
  wire[3:0] T4156;
  reg [3:0] counts_684;
  wire[3:0] T11029;
  wire[3:0] T4157;
  wire[3:0] T4158;
  wire T4159;
  wire T4160;
  reg [3:0] counts_685;
  wire[3:0] T11030;
  wire[3:0] T4161;
  wire[3:0] T4162;
  wire T4163;
  wire T4164;
  wire T4165;
  wire[3:0] T4166;
  reg [3:0] counts_686;
  wire[3:0] T11031;
  wire[3:0] T4167;
  wire[3:0] T4168;
  wire T4169;
  wire T4170;
  reg [3:0] counts_687;
  wire[3:0] T11032;
  wire[3:0] T4171;
  wire[3:0] T4172;
  wire T4173;
  wire T4174;
  wire T4175;
  wire T4176;
  wire T4177;
  wire T4178;
  wire[3:0] T4179;
  wire[3:0] T4180;
  wire[3:0] T4181;
  wire[3:0] T4182;
  reg [3:0] counts_688;
  wire[3:0] T11033;
  wire[3:0] T4183;
  wire[3:0] T4184;
  wire T4185;
  wire T4186;
  reg [3:0] counts_689;
  wire[3:0] T11034;
  wire[3:0] T4187;
  wire[3:0] T4188;
  wire T4189;
  wire T4190;
  wire T4191;
  wire[3:0] T4192;
  reg [3:0] counts_690;
  wire[3:0] T11035;
  wire[3:0] T4193;
  wire[3:0] T4194;
  wire T4195;
  wire T4196;
  reg [3:0] counts_691;
  wire[3:0] T11036;
  wire[3:0] T4197;
  wire[3:0] T4198;
  wire T4199;
  wire T4200;
  wire T4201;
  wire T4202;
  wire[3:0] T4203;
  wire[3:0] T4204;
  reg [3:0] counts_692;
  wire[3:0] T11037;
  wire[3:0] T4205;
  wire[3:0] T4206;
  wire T4207;
  wire T4208;
  reg [3:0] counts_693;
  wire[3:0] T11038;
  wire[3:0] T4209;
  wire[3:0] T4210;
  wire T4211;
  wire T4212;
  wire T4213;
  wire[3:0] T4214;
  reg [3:0] counts_694;
  wire[3:0] T11039;
  wire[3:0] T4215;
  wire[3:0] T4216;
  wire T4217;
  wire T4218;
  reg [3:0] counts_695;
  wire[3:0] T11040;
  wire[3:0] T4219;
  wire[3:0] T4220;
  wire T4221;
  wire T4222;
  wire T4223;
  wire T4224;
  wire T4225;
  wire[3:0] T4226;
  wire[3:0] T4227;
  wire[3:0] T4228;
  reg [3:0] counts_696;
  wire[3:0] T11041;
  wire[3:0] T4229;
  wire[3:0] T4230;
  wire T4231;
  wire T4232;
  reg [3:0] counts_697;
  wire[3:0] T11042;
  wire[3:0] T4233;
  wire[3:0] T4234;
  wire T4235;
  wire T4236;
  wire T4237;
  wire[3:0] T4238;
  reg [3:0] counts_698;
  wire[3:0] T11043;
  wire[3:0] T4239;
  wire[3:0] T4240;
  wire T4241;
  wire T4242;
  reg [3:0] counts_699;
  wire[3:0] T11044;
  wire[3:0] T4243;
  wire[3:0] T4244;
  wire T4245;
  wire T4246;
  wire T4247;
  wire T4248;
  wire[3:0] T4249;
  wire[3:0] T4250;
  reg [3:0] counts_700;
  wire[3:0] T11045;
  wire[3:0] T4251;
  wire[3:0] T4252;
  wire T4253;
  wire T4254;
  reg [3:0] counts_701;
  wire[3:0] T11046;
  wire[3:0] T4255;
  wire[3:0] T4256;
  wire T4257;
  wire T4258;
  wire T4259;
  wire[3:0] T4260;
  reg [3:0] counts_702;
  wire[3:0] T11047;
  wire[3:0] T4261;
  wire[3:0] T4262;
  wire T4263;
  wire T4264;
  reg [3:0] counts_703;
  wire[3:0] T11048;
  wire[3:0] T4265;
  wire[3:0] T4266;
  wire T4267;
  wire T4268;
  wire T4269;
  wire T4270;
  wire T4271;
  wire T4272;
  wire T4273;
  wire T4274;
  wire[3:0] T4275;
  wire[3:0] T4276;
  wire[3:0] T4277;
  wire[3:0] T4278;
  wire[3:0] T4279;
  wire[3:0] T4280;
  reg [3:0] counts_704;
  wire[3:0] T11049;
  wire[3:0] T4281;
  wire[3:0] T4282;
  wire T4283;
  wire T4284;
  reg [3:0] counts_705;
  wire[3:0] T11050;
  wire[3:0] T4285;
  wire[3:0] T4286;
  wire T4287;
  wire T4288;
  wire T4289;
  wire[3:0] T4290;
  reg [3:0] counts_706;
  wire[3:0] T11051;
  wire[3:0] T4291;
  wire[3:0] T4292;
  wire T4293;
  wire T4294;
  reg [3:0] counts_707;
  wire[3:0] T11052;
  wire[3:0] T4295;
  wire[3:0] T4296;
  wire T4297;
  wire T4298;
  wire T4299;
  wire T4300;
  wire[3:0] T4301;
  wire[3:0] T4302;
  reg [3:0] counts_708;
  wire[3:0] T11053;
  wire[3:0] T4303;
  wire[3:0] T4304;
  wire T4305;
  wire T4306;
  reg [3:0] counts_709;
  wire[3:0] T11054;
  wire[3:0] T4307;
  wire[3:0] T4308;
  wire T4309;
  wire T4310;
  wire T4311;
  wire[3:0] T4312;
  reg [3:0] counts_710;
  wire[3:0] T11055;
  wire[3:0] T4313;
  wire[3:0] T4314;
  wire T4315;
  wire T4316;
  reg [3:0] counts_711;
  wire[3:0] T11056;
  wire[3:0] T4317;
  wire[3:0] T4318;
  wire T4319;
  wire T4320;
  wire T4321;
  wire T4322;
  wire T4323;
  wire[3:0] T4324;
  wire[3:0] T4325;
  wire[3:0] T4326;
  reg [3:0] counts_712;
  wire[3:0] T11057;
  wire[3:0] T4327;
  wire[3:0] T4328;
  wire T4329;
  wire T4330;
  reg [3:0] counts_713;
  wire[3:0] T11058;
  wire[3:0] T4331;
  wire[3:0] T4332;
  wire T4333;
  wire T4334;
  wire T4335;
  wire[3:0] T4336;
  reg [3:0] counts_714;
  wire[3:0] T11059;
  wire[3:0] T4337;
  wire[3:0] T4338;
  wire T4339;
  wire T4340;
  reg [3:0] counts_715;
  wire[3:0] T11060;
  wire[3:0] T4341;
  wire[3:0] T4342;
  wire T4343;
  wire T4344;
  wire T4345;
  wire T4346;
  wire[3:0] T4347;
  wire[3:0] T4348;
  reg [3:0] counts_716;
  wire[3:0] T11061;
  wire[3:0] T4349;
  wire[3:0] T4350;
  wire T4351;
  wire T4352;
  reg [3:0] counts_717;
  wire[3:0] T11062;
  wire[3:0] T4353;
  wire[3:0] T4354;
  wire T4355;
  wire T4356;
  wire T4357;
  wire[3:0] T4358;
  reg [3:0] counts_718;
  wire[3:0] T11063;
  wire[3:0] T4359;
  wire[3:0] T4360;
  wire T4361;
  wire T4362;
  reg [3:0] counts_719;
  wire[3:0] T11064;
  wire[3:0] T4363;
  wire[3:0] T4364;
  wire T4365;
  wire T4366;
  wire T4367;
  wire T4368;
  wire T4369;
  wire T4370;
  wire[3:0] T4371;
  wire[3:0] T4372;
  wire[3:0] T4373;
  wire[3:0] T4374;
  reg [3:0] counts_720;
  wire[3:0] T11065;
  wire[3:0] T4375;
  wire[3:0] T4376;
  wire T4377;
  wire T4378;
  reg [3:0] counts_721;
  wire[3:0] T11066;
  wire[3:0] T4379;
  wire[3:0] T4380;
  wire T4381;
  wire T4382;
  wire T4383;
  wire[3:0] T4384;
  reg [3:0] counts_722;
  wire[3:0] T11067;
  wire[3:0] T4385;
  wire[3:0] T4386;
  wire T4387;
  wire T4388;
  reg [3:0] counts_723;
  wire[3:0] T11068;
  wire[3:0] T4389;
  wire[3:0] T4390;
  wire T4391;
  wire T4392;
  wire T4393;
  wire T4394;
  wire[3:0] T4395;
  wire[3:0] T4396;
  reg [3:0] counts_724;
  wire[3:0] T11069;
  wire[3:0] T4397;
  wire[3:0] T4398;
  wire T4399;
  wire T4400;
  reg [3:0] counts_725;
  wire[3:0] T11070;
  wire[3:0] T4401;
  wire[3:0] T4402;
  wire T4403;
  wire T4404;
  wire T4405;
  wire[3:0] T4406;
  reg [3:0] counts_726;
  wire[3:0] T11071;
  wire[3:0] T4407;
  wire[3:0] T4408;
  wire T4409;
  wire T4410;
  reg [3:0] counts_727;
  wire[3:0] T11072;
  wire[3:0] T4411;
  wire[3:0] T4412;
  wire T4413;
  wire T4414;
  wire T4415;
  wire T4416;
  wire T4417;
  wire[3:0] T4418;
  wire[3:0] T4419;
  wire[3:0] T4420;
  reg [3:0] counts_728;
  wire[3:0] T11073;
  wire[3:0] T4421;
  wire[3:0] T4422;
  wire T4423;
  wire T4424;
  reg [3:0] counts_729;
  wire[3:0] T11074;
  wire[3:0] T4425;
  wire[3:0] T4426;
  wire T4427;
  wire T4428;
  wire T4429;
  wire[3:0] T4430;
  reg [3:0] counts_730;
  wire[3:0] T11075;
  wire[3:0] T4431;
  wire[3:0] T4432;
  wire T4433;
  wire T4434;
  reg [3:0] counts_731;
  wire[3:0] T11076;
  wire[3:0] T4435;
  wire[3:0] T4436;
  wire T4437;
  wire T4438;
  wire T4439;
  wire T4440;
  wire[3:0] T4441;
  wire[3:0] T4442;
  reg [3:0] counts_732;
  wire[3:0] T11077;
  wire[3:0] T4443;
  wire[3:0] T4444;
  wire T4445;
  wire T4446;
  reg [3:0] counts_733;
  wire[3:0] T11078;
  wire[3:0] T4447;
  wire[3:0] T4448;
  wire T4449;
  wire T4450;
  wire T4451;
  wire[3:0] T4452;
  reg [3:0] counts_734;
  wire[3:0] T11079;
  wire[3:0] T4453;
  wire[3:0] T4454;
  wire T4455;
  wire T4456;
  reg [3:0] counts_735;
  wire[3:0] T11080;
  wire[3:0] T4457;
  wire[3:0] T4458;
  wire T4459;
  wire T4460;
  wire T4461;
  wire T4462;
  wire T4463;
  wire T4464;
  wire T4465;
  wire[3:0] T4466;
  wire[3:0] T4467;
  wire[3:0] T4468;
  wire[3:0] T4469;
  wire[3:0] T4470;
  reg [3:0] counts_736;
  wire[3:0] T11081;
  wire[3:0] T4471;
  wire[3:0] T4472;
  wire T4473;
  wire T4474;
  reg [3:0] counts_737;
  wire[3:0] T11082;
  wire[3:0] T4475;
  wire[3:0] T4476;
  wire T4477;
  wire T4478;
  wire T4479;
  wire[3:0] T4480;
  reg [3:0] counts_738;
  wire[3:0] T11083;
  wire[3:0] T4481;
  wire[3:0] T4482;
  wire T4483;
  wire T4484;
  reg [3:0] counts_739;
  wire[3:0] T11084;
  wire[3:0] T4485;
  wire[3:0] T4486;
  wire T4487;
  wire T4488;
  wire T4489;
  wire T4490;
  wire[3:0] T4491;
  wire[3:0] T4492;
  reg [3:0] counts_740;
  wire[3:0] T11085;
  wire[3:0] T4493;
  wire[3:0] T4494;
  wire T4495;
  wire T4496;
  reg [3:0] counts_741;
  wire[3:0] T11086;
  wire[3:0] T4497;
  wire[3:0] T4498;
  wire T4499;
  wire T4500;
  wire T4501;
  wire[3:0] T4502;
  reg [3:0] counts_742;
  wire[3:0] T11087;
  wire[3:0] T4503;
  wire[3:0] T4504;
  wire T4505;
  wire T4506;
  reg [3:0] counts_743;
  wire[3:0] T11088;
  wire[3:0] T4507;
  wire[3:0] T4508;
  wire T4509;
  wire T4510;
  wire T4511;
  wire T4512;
  wire T4513;
  wire[3:0] T4514;
  wire[3:0] T4515;
  wire[3:0] T4516;
  reg [3:0] counts_744;
  wire[3:0] T11089;
  wire[3:0] T4517;
  wire[3:0] T4518;
  wire T4519;
  wire T4520;
  reg [3:0] counts_745;
  wire[3:0] T11090;
  wire[3:0] T4521;
  wire[3:0] T4522;
  wire T4523;
  wire T4524;
  wire T4525;
  wire[3:0] T4526;
  reg [3:0] counts_746;
  wire[3:0] T11091;
  wire[3:0] T4527;
  wire[3:0] T4528;
  wire T4529;
  wire T4530;
  reg [3:0] counts_747;
  wire[3:0] T11092;
  wire[3:0] T4531;
  wire[3:0] T4532;
  wire T4533;
  wire T4534;
  wire T4535;
  wire T4536;
  wire[3:0] T4537;
  wire[3:0] T4538;
  reg [3:0] counts_748;
  wire[3:0] T11093;
  wire[3:0] T4539;
  wire[3:0] T4540;
  wire T4541;
  wire T4542;
  reg [3:0] counts_749;
  wire[3:0] T11094;
  wire[3:0] T4543;
  wire[3:0] T4544;
  wire T4545;
  wire T4546;
  wire T4547;
  wire[3:0] T4548;
  reg [3:0] counts_750;
  wire[3:0] T11095;
  wire[3:0] T4549;
  wire[3:0] T4550;
  wire T4551;
  wire T4552;
  reg [3:0] counts_751;
  wire[3:0] T11096;
  wire[3:0] T4553;
  wire[3:0] T4554;
  wire T4555;
  wire T4556;
  wire T4557;
  wire T4558;
  wire T4559;
  wire T4560;
  wire[3:0] T4561;
  wire[3:0] T4562;
  wire[3:0] T4563;
  wire[3:0] T4564;
  reg [3:0] counts_752;
  wire[3:0] T11097;
  wire[3:0] T4565;
  wire[3:0] T4566;
  wire T4567;
  wire T4568;
  reg [3:0] counts_753;
  wire[3:0] T11098;
  wire[3:0] T4569;
  wire[3:0] T4570;
  wire T4571;
  wire T4572;
  wire T4573;
  wire[3:0] T4574;
  reg [3:0] counts_754;
  wire[3:0] T11099;
  wire[3:0] T4575;
  wire[3:0] T4576;
  wire T4577;
  wire T4578;
  reg [3:0] counts_755;
  wire[3:0] T11100;
  wire[3:0] T4579;
  wire[3:0] T4580;
  wire T4581;
  wire T4582;
  wire T4583;
  wire T4584;
  wire[3:0] T4585;
  wire[3:0] T4586;
  reg [3:0] counts_756;
  wire[3:0] T11101;
  wire[3:0] T4587;
  wire[3:0] T4588;
  wire T4589;
  wire T4590;
  reg [3:0] counts_757;
  wire[3:0] T11102;
  wire[3:0] T4591;
  wire[3:0] T4592;
  wire T4593;
  wire T4594;
  wire T4595;
  wire[3:0] T4596;
  reg [3:0] counts_758;
  wire[3:0] T11103;
  wire[3:0] T4597;
  wire[3:0] T4598;
  wire T4599;
  wire T4600;
  reg [3:0] counts_759;
  wire[3:0] T11104;
  wire[3:0] T4601;
  wire[3:0] T4602;
  wire T4603;
  wire T4604;
  wire T4605;
  wire T4606;
  wire T4607;
  wire[3:0] T4608;
  wire[3:0] T4609;
  wire[3:0] T4610;
  reg [3:0] counts_760;
  wire[3:0] T11105;
  wire[3:0] T4611;
  wire[3:0] T4612;
  wire T4613;
  wire T4614;
  reg [3:0] counts_761;
  wire[3:0] T11106;
  wire[3:0] T4615;
  wire[3:0] T4616;
  wire T4617;
  wire T4618;
  wire T4619;
  wire[3:0] T4620;
  reg [3:0] counts_762;
  wire[3:0] T11107;
  wire[3:0] T4621;
  wire[3:0] T4622;
  wire T4623;
  wire T4624;
  reg [3:0] counts_763;
  wire[3:0] T11108;
  wire[3:0] T4625;
  wire[3:0] T4626;
  wire T4627;
  wire T4628;
  wire T4629;
  wire T4630;
  wire[3:0] T4631;
  wire[3:0] T4632;
  reg [3:0] counts_764;
  wire[3:0] T11109;
  wire[3:0] T4633;
  wire[3:0] T4634;
  wire T4635;
  wire T4636;
  reg [3:0] counts_765;
  wire[3:0] T11110;
  wire[3:0] T4637;
  wire[3:0] T4638;
  wire T4639;
  wire T4640;
  wire T4641;
  wire[3:0] T4642;
  reg [3:0] counts_766;
  wire[3:0] T11111;
  wire[3:0] T4643;
  wire[3:0] T4644;
  wire T4645;
  wire T4646;
  reg [3:0] counts_767;
  wire[3:0] T11112;
  wire[3:0] T4647;
  wire[3:0] T4648;
  wire T4649;
  wire T4650;
  wire T4651;
  wire T4652;
  wire T4653;
  wire T4654;
  wire T4655;
  wire T4656;
  wire T4657;
  wire T4658;
  wire[3:0] T4659;
  wire[3:0] T4660;
  wire[3:0] T4661;
  wire[3:0] T4662;
  wire[3:0] T4663;
  wire[3:0] T4664;
  wire[3:0] T4665;
  wire[3:0] T4666;
  reg [3:0] counts_768;
  wire[3:0] T11113;
  wire[3:0] T4667;
  wire[3:0] T4668;
  wire T4669;
  wire T4670;
  reg [3:0] counts_769;
  wire[3:0] T11114;
  wire[3:0] T4671;
  wire[3:0] T4672;
  wire T4673;
  wire T4674;
  wire T4675;
  wire[3:0] T4676;
  reg [3:0] counts_770;
  wire[3:0] T11115;
  wire[3:0] T4677;
  wire[3:0] T4678;
  wire T4679;
  wire T4680;
  reg [3:0] counts_771;
  wire[3:0] T11116;
  wire[3:0] T4681;
  wire[3:0] T4682;
  wire T4683;
  wire T4684;
  wire T4685;
  wire T4686;
  wire[3:0] T4687;
  wire[3:0] T4688;
  reg [3:0] counts_772;
  wire[3:0] T11117;
  wire[3:0] T4689;
  wire[3:0] T4690;
  wire T4691;
  wire T4692;
  reg [3:0] counts_773;
  wire[3:0] T11118;
  wire[3:0] T4693;
  wire[3:0] T4694;
  wire T4695;
  wire T4696;
  wire T4697;
  wire[3:0] T4698;
  reg [3:0] counts_774;
  wire[3:0] T11119;
  wire[3:0] T4699;
  wire[3:0] T4700;
  wire T4701;
  wire T4702;
  reg [3:0] counts_775;
  wire[3:0] T11120;
  wire[3:0] T4703;
  wire[3:0] T4704;
  wire T4705;
  wire T4706;
  wire T4707;
  wire T4708;
  wire T4709;
  wire[3:0] T4710;
  wire[3:0] T4711;
  wire[3:0] T4712;
  reg [3:0] counts_776;
  wire[3:0] T11121;
  wire[3:0] T4713;
  wire[3:0] T4714;
  wire T4715;
  wire T4716;
  reg [3:0] counts_777;
  wire[3:0] T11122;
  wire[3:0] T4717;
  wire[3:0] T4718;
  wire T4719;
  wire T4720;
  wire T4721;
  wire[3:0] T4722;
  reg [3:0] counts_778;
  wire[3:0] T11123;
  wire[3:0] T4723;
  wire[3:0] T4724;
  wire T4725;
  wire T4726;
  reg [3:0] counts_779;
  wire[3:0] T11124;
  wire[3:0] T4727;
  wire[3:0] T4728;
  wire T4729;
  wire T4730;
  wire T4731;
  wire T4732;
  wire[3:0] T4733;
  wire[3:0] T4734;
  reg [3:0] counts_780;
  wire[3:0] T11125;
  wire[3:0] T4735;
  wire[3:0] T4736;
  wire T4737;
  wire T4738;
  reg [3:0] counts_781;
  wire[3:0] T11126;
  wire[3:0] T4739;
  wire[3:0] T4740;
  wire T4741;
  wire T4742;
  wire T4743;
  wire[3:0] T4744;
  reg [3:0] counts_782;
  wire[3:0] T11127;
  wire[3:0] T4745;
  wire[3:0] T4746;
  wire T4747;
  wire T4748;
  reg [3:0] counts_783;
  wire[3:0] T11128;
  wire[3:0] T4749;
  wire[3:0] T4750;
  wire T4751;
  wire T4752;
  wire T4753;
  wire T4754;
  wire T4755;
  wire T4756;
  wire[3:0] T4757;
  wire[3:0] T4758;
  wire[3:0] T4759;
  wire[3:0] T4760;
  reg [3:0] counts_784;
  wire[3:0] T11129;
  wire[3:0] T4761;
  wire[3:0] T4762;
  wire T4763;
  wire T4764;
  reg [3:0] counts_785;
  wire[3:0] T11130;
  wire[3:0] T4765;
  wire[3:0] T4766;
  wire T4767;
  wire T4768;
  wire T4769;
  wire[3:0] T4770;
  reg [3:0] counts_786;
  wire[3:0] T11131;
  wire[3:0] T4771;
  wire[3:0] T4772;
  wire T4773;
  wire T4774;
  reg [3:0] counts_787;
  wire[3:0] T11132;
  wire[3:0] T4775;
  wire[3:0] T4776;
  wire T4777;
  wire T4778;
  wire T4779;
  wire T4780;
  wire[3:0] T4781;
  wire[3:0] T4782;
  reg [3:0] counts_788;
  wire[3:0] T11133;
  wire[3:0] T4783;
  wire[3:0] T4784;
  wire T4785;
  wire T4786;
  reg [3:0] counts_789;
  wire[3:0] T11134;
  wire[3:0] T4787;
  wire[3:0] T4788;
  wire T4789;
  wire T4790;
  wire T4791;
  wire[3:0] T4792;
  reg [3:0] counts_790;
  wire[3:0] T11135;
  wire[3:0] T4793;
  wire[3:0] T4794;
  wire T4795;
  wire T4796;
  reg [3:0] counts_791;
  wire[3:0] T11136;
  wire[3:0] T4797;
  wire[3:0] T4798;
  wire T4799;
  wire T4800;
  wire T4801;
  wire T4802;
  wire T4803;
  wire[3:0] T4804;
  wire[3:0] T4805;
  wire[3:0] T4806;
  reg [3:0] counts_792;
  wire[3:0] T11137;
  wire[3:0] T4807;
  wire[3:0] T4808;
  wire T4809;
  wire T4810;
  reg [3:0] counts_793;
  wire[3:0] T11138;
  wire[3:0] T4811;
  wire[3:0] T4812;
  wire T4813;
  wire T4814;
  wire T4815;
  wire[3:0] T4816;
  reg [3:0] counts_794;
  wire[3:0] T11139;
  wire[3:0] T4817;
  wire[3:0] T4818;
  wire T4819;
  wire T4820;
  reg [3:0] counts_795;
  wire[3:0] T11140;
  wire[3:0] T4821;
  wire[3:0] T4822;
  wire T4823;
  wire T4824;
  wire T4825;
  wire T4826;
  wire[3:0] T4827;
  wire[3:0] T4828;
  reg [3:0] counts_796;
  wire[3:0] T11141;
  wire[3:0] T4829;
  wire[3:0] T4830;
  wire T4831;
  wire T4832;
  reg [3:0] counts_797;
  wire[3:0] T11142;
  wire[3:0] T4833;
  wire[3:0] T4834;
  wire T4835;
  wire T4836;
  wire T4837;
  wire[3:0] T4838;
  reg [3:0] counts_798;
  wire[3:0] T11143;
  wire[3:0] T4839;
  wire[3:0] T4840;
  wire T4841;
  wire T4842;
  reg [3:0] counts_799;
  wire[3:0] T11144;
  wire[3:0] T4843;
  wire[3:0] T4844;
  wire T4845;
  wire T4846;
  wire T4847;
  wire T4848;
  wire T4849;
  wire T4850;
  wire T4851;
  wire[3:0] T4852;
  wire[3:0] T4853;
  wire[3:0] T4854;
  wire[3:0] T4855;
  wire[3:0] T4856;
  reg [3:0] counts_800;
  wire[3:0] T11145;
  wire[3:0] T4857;
  wire[3:0] T4858;
  wire T4859;
  wire T4860;
  reg [3:0] counts_801;
  wire[3:0] T11146;
  wire[3:0] T4861;
  wire[3:0] T4862;
  wire T4863;
  wire T4864;
  wire T4865;
  wire[3:0] T4866;
  reg [3:0] counts_802;
  wire[3:0] T11147;
  wire[3:0] T4867;
  wire[3:0] T4868;
  wire T4869;
  wire T4870;
  reg [3:0] counts_803;
  wire[3:0] T11148;
  wire[3:0] T4871;
  wire[3:0] T4872;
  wire T4873;
  wire T4874;
  wire T4875;
  wire T4876;
  wire[3:0] T4877;
  wire[3:0] T4878;
  reg [3:0] counts_804;
  wire[3:0] T11149;
  wire[3:0] T4879;
  wire[3:0] T4880;
  wire T4881;
  wire T4882;
  reg [3:0] counts_805;
  wire[3:0] T11150;
  wire[3:0] T4883;
  wire[3:0] T4884;
  wire T4885;
  wire T4886;
  wire T4887;
  wire[3:0] T4888;
  reg [3:0] counts_806;
  wire[3:0] T11151;
  wire[3:0] T4889;
  wire[3:0] T4890;
  wire T4891;
  wire T4892;
  reg [3:0] counts_807;
  wire[3:0] T11152;
  wire[3:0] T4893;
  wire[3:0] T4894;
  wire T4895;
  wire T4896;
  wire T4897;
  wire T4898;
  wire T4899;
  wire[3:0] T4900;
  wire[3:0] T4901;
  wire[3:0] T4902;
  reg [3:0] counts_808;
  wire[3:0] T11153;
  wire[3:0] T4903;
  wire[3:0] T4904;
  wire T4905;
  wire T4906;
  reg [3:0] counts_809;
  wire[3:0] T11154;
  wire[3:0] T4907;
  wire[3:0] T4908;
  wire T4909;
  wire T4910;
  wire T4911;
  wire[3:0] T4912;
  reg [3:0] counts_810;
  wire[3:0] T11155;
  wire[3:0] T4913;
  wire[3:0] T4914;
  wire T4915;
  wire T4916;
  reg [3:0] counts_811;
  wire[3:0] T11156;
  wire[3:0] T4917;
  wire[3:0] T4918;
  wire T4919;
  wire T4920;
  wire T4921;
  wire T4922;
  wire[3:0] T4923;
  wire[3:0] T4924;
  reg [3:0] counts_812;
  wire[3:0] T11157;
  wire[3:0] T4925;
  wire[3:0] T4926;
  wire T4927;
  wire T4928;
  reg [3:0] counts_813;
  wire[3:0] T11158;
  wire[3:0] T4929;
  wire[3:0] T4930;
  wire T4931;
  wire T4932;
  wire T4933;
  wire[3:0] T4934;
  reg [3:0] counts_814;
  wire[3:0] T11159;
  wire[3:0] T4935;
  wire[3:0] T4936;
  wire T4937;
  wire T4938;
  reg [3:0] counts_815;
  wire[3:0] T11160;
  wire[3:0] T4939;
  wire[3:0] T4940;
  wire T4941;
  wire T4942;
  wire T4943;
  wire T4944;
  wire T4945;
  wire T4946;
  wire[3:0] T4947;
  wire[3:0] T4948;
  wire[3:0] T4949;
  wire[3:0] T4950;
  reg [3:0] counts_816;
  wire[3:0] T11161;
  wire[3:0] T4951;
  wire[3:0] T4952;
  wire T4953;
  wire T4954;
  reg [3:0] counts_817;
  wire[3:0] T11162;
  wire[3:0] T4955;
  wire[3:0] T4956;
  wire T4957;
  wire T4958;
  wire T4959;
  wire[3:0] T4960;
  reg [3:0] counts_818;
  wire[3:0] T11163;
  wire[3:0] T4961;
  wire[3:0] T4962;
  wire T4963;
  wire T4964;
  reg [3:0] counts_819;
  wire[3:0] T11164;
  wire[3:0] T4965;
  wire[3:0] T4966;
  wire T4967;
  wire T4968;
  wire T4969;
  wire T4970;
  wire[3:0] T4971;
  wire[3:0] T4972;
  reg [3:0] counts_820;
  wire[3:0] T11165;
  wire[3:0] T4973;
  wire[3:0] T4974;
  wire T4975;
  wire T4976;
  reg [3:0] counts_821;
  wire[3:0] T11166;
  wire[3:0] T4977;
  wire[3:0] T4978;
  wire T4979;
  wire T4980;
  wire T4981;
  wire[3:0] T4982;
  reg [3:0] counts_822;
  wire[3:0] T11167;
  wire[3:0] T4983;
  wire[3:0] T4984;
  wire T4985;
  wire T4986;
  reg [3:0] counts_823;
  wire[3:0] T11168;
  wire[3:0] T4987;
  wire[3:0] T4988;
  wire T4989;
  wire T4990;
  wire T4991;
  wire T4992;
  wire T4993;
  wire[3:0] T4994;
  wire[3:0] T4995;
  wire[3:0] T4996;
  reg [3:0] counts_824;
  wire[3:0] T11169;
  wire[3:0] T4997;
  wire[3:0] T4998;
  wire T4999;
  wire T5000;
  reg [3:0] counts_825;
  wire[3:0] T11170;
  wire[3:0] T5001;
  wire[3:0] T5002;
  wire T5003;
  wire T5004;
  wire T5005;
  wire[3:0] T5006;
  reg [3:0] counts_826;
  wire[3:0] T11171;
  wire[3:0] T5007;
  wire[3:0] T5008;
  wire T5009;
  wire T5010;
  reg [3:0] counts_827;
  wire[3:0] T11172;
  wire[3:0] T5011;
  wire[3:0] T5012;
  wire T5013;
  wire T5014;
  wire T5015;
  wire T5016;
  wire[3:0] T5017;
  wire[3:0] T5018;
  reg [3:0] counts_828;
  wire[3:0] T11173;
  wire[3:0] T5019;
  wire[3:0] T5020;
  wire T5021;
  wire T5022;
  reg [3:0] counts_829;
  wire[3:0] T11174;
  wire[3:0] T5023;
  wire[3:0] T5024;
  wire T5025;
  wire T5026;
  wire T5027;
  wire[3:0] T5028;
  reg [3:0] counts_830;
  wire[3:0] T11175;
  wire[3:0] T5029;
  wire[3:0] T5030;
  wire T5031;
  wire T5032;
  reg [3:0] counts_831;
  wire[3:0] T11176;
  wire[3:0] T5033;
  wire[3:0] T5034;
  wire T5035;
  wire T5036;
  wire T5037;
  wire T5038;
  wire T5039;
  wire T5040;
  wire T5041;
  wire T5042;
  wire[3:0] T5043;
  wire[3:0] T5044;
  wire[3:0] T5045;
  wire[3:0] T5046;
  wire[3:0] T5047;
  wire[3:0] T5048;
  reg [3:0] counts_832;
  wire[3:0] T11177;
  wire[3:0] T5049;
  wire[3:0] T5050;
  wire T5051;
  wire T5052;
  reg [3:0] counts_833;
  wire[3:0] T11178;
  wire[3:0] T5053;
  wire[3:0] T5054;
  wire T5055;
  wire T5056;
  wire T5057;
  wire[3:0] T5058;
  reg [3:0] counts_834;
  wire[3:0] T11179;
  wire[3:0] T5059;
  wire[3:0] T5060;
  wire T5061;
  wire T5062;
  reg [3:0] counts_835;
  wire[3:0] T11180;
  wire[3:0] T5063;
  wire[3:0] T5064;
  wire T5065;
  wire T5066;
  wire T5067;
  wire T5068;
  wire[3:0] T5069;
  wire[3:0] T5070;
  reg [3:0] counts_836;
  wire[3:0] T11181;
  wire[3:0] T5071;
  wire[3:0] T5072;
  wire T5073;
  wire T5074;
  reg [3:0] counts_837;
  wire[3:0] T11182;
  wire[3:0] T5075;
  wire[3:0] T5076;
  wire T5077;
  wire T5078;
  wire T5079;
  wire[3:0] T5080;
  reg [3:0] counts_838;
  wire[3:0] T11183;
  wire[3:0] T5081;
  wire[3:0] T5082;
  wire T5083;
  wire T5084;
  reg [3:0] counts_839;
  wire[3:0] T11184;
  wire[3:0] T5085;
  wire[3:0] T5086;
  wire T5087;
  wire T5088;
  wire T5089;
  wire T5090;
  wire T5091;
  wire[3:0] T5092;
  wire[3:0] T5093;
  wire[3:0] T5094;
  reg [3:0] counts_840;
  wire[3:0] T11185;
  wire[3:0] T5095;
  wire[3:0] T5096;
  wire T5097;
  wire T5098;
  reg [3:0] counts_841;
  wire[3:0] T11186;
  wire[3:0] T5099;
  wire[3:0] T5100;
  wire T5101;
  wire T5102;
  wire T5103;
  wire[3:0] T5104;
  reg [3:0] counts_842;
  wire[3:0] T11187;
  wire[3:0] T5105;
  wire[3:0] T5106;
  wire T5107;
  wire T5108;
  reg [3:0] counts_843;
  wire[3:0] T11188;
  wire[3:0] T5109;
  wire[3:0] T5110;
  wire T5111;
  wire T5112;
  wire T5113;
  wire T5114;
  wire[3:0] T5115;
  wire[3:0] T5116;
  reg [3:0] counts_844;
  wire[3:0] T11189;
  wire[3:0] T5117;
  wire[3:0] T5118;
  wire T5119;
  wire T5120;
  reg [3:0] counts_845;
  wire[3:0] T11190;
  wire[3:0] T5121;
  wire[3:0] T5122;
  wire T5123;
  wire T5124;
  wire T5125;
  wire[3:0] T5126;
  reg [3:0] counts_846;
  wire[3:0] T11191;
  wire[3:0] T5127;
  wire[3:0] T5128;
  wire T5129;
  wire T5130;
  reg [3:0] counts_847;
  wire[3:0] T11192;
  wire[3:0] T5131;
  wire[3:0] T5132;
  wire T5133;
  wire T5134;
  wire T5135;
  wire T5136;
  wire T5137;
  wire T5138;
  wire[3:0] T5139;
  wire[3:0] T5140;
  wire[3:0] T5141;
  wire[3:0] T5142;
  reg [3:0] counts_848;
  wire[3:0] T11193;
  wire[3:0] T5143;
  wire[3:0] T5144;
  wire T5145;
  wire T5146;
  reg [3:0] counts_849;
  wire[3:0] T11194;
  wire[3:0] T5147;
  wire[3:0] T5148;
  wire T5149;
  wire T5150;
  wire T5151;
  wire[3:0] T5152;
  reg [3:0] counts_850;
  wire[3:0] T11195;
  wire[3:0] T5153;
  wire[3:0] T5154;
  wire T5155;
  wire T5156;
  reg [3:0] counts_851;
  wire[3:0] T11196;
  wire[3:0] T5157;
  wire[3:0] T5158;
  wire T5159;
  wire T5160;
  wire T5161;
  wire T5162;
  wire[3:0] T5163;
  wire[3:0] T5164;
  reg [3:0] counts_852;
  wire[3:0] T11197;
  wire[3:0] T5165;
  wire[3:0] T5166;
  wire T5167;
  wire T5168;
  reg [3:0] counts_853;
  wire[3:0] T11198;
  wire[3:0] T5169;
  wire[3:0] T5170;
  wire T5171;
  wire T5172;
  wire T5173;
  wire[3:0] T5174;
  reg [3:0] counts_854;
  wire[3:0] T11199;
  wire[3:0] T5175;
  wire[3:0] T5176;
  wire T5177;
  wire T5178;
  reg [3:0] counts_855;
  wire[3:0] T11200;
  wire[3:0] T5179;
  wire[3:0] T5180;
  wire T5181;
  wire T5182;
  wire T5183;
  wire T5184;
  wire T5185;
  wire[3:0] T5186;
  wire[3:0] T5187;
  wire[3:0] T5188;
  reg [3:0] counts_856;
  wire[3:0] T11201;
  wire[3:0] T5189;
  wire[3:0] T5190;
  wire T5191;
  wire T5192;
  reg [3:0] counts_857;
  wire[3:0] T11202;
  wire[3:0] T5193;
  wire[3:0] T5194;
  wire T5195;
  wire T5196;
  wire T5197;
  wire[3:0] T5198;
  reg [3:0] counts_858;
  wire[3:0] T11203;
  wire[3:0] T5199;
  wire[3:0] T5200;
  wire T5201;
  wire T5202;
  reg [3:0] counts_859;
  wire[3:0] T11204;
  wire[3:0] T5203;
  wire[3:0] T5204;
  wire T5205;
  wire T5206;
  wire T5207;
  wire T5208;
  wire[3:0] T5209;
  wire[3:0] T5210;
  reg [3:0] counts_860;
  wire[3:0] T11205;
  wire[3:0] T5211;
  wire[3:0] T5212;
  wire T5213;
  wire T5214;
  reg [3:0] counts_861;
  wire[3:0] T11206;
  wire[3:0] T5215;
  wire[3:0] T5216;
  wire T5217;
  wire T5218;
  wire T5219;
  wire[3:0] T5220;
  reg [3:0] counts_862;
  wire[3:0] T11207;
  wire[3:0] T5221;
  wire[3:0] T5222;
  wire T5223;
  wire T5224;
  reg [3:0] counts_863;
  wire[3:0] T11208;
  wire[3:0] T5225;
  wire[3:0] T5226;
  wire T5227;
  wire T5228;
  wire T5229;
  wire T5230;
  wire T5231;
  wire T5232;
  wire T5233;
  wire[3:0] T5234;
  wire[3:0] T5235;
  wire[3:0] T5236;
  wire[3:0] T5237;
  wire[3:0] T5238;
  reg [3:0] counts_864;
  wire[3:0] T11209;
  wire[3:0] T5239;
  wire[3:0] T5240;
  wire T5241;
  wire T5242;
  reg [3:0] counts_865;
  wire[3:0] T11210;
  wire[3:0] T5243;
  wire[3:0] T5244;
  wire T5245;
  wire T5246;
  wire T5247;
  wire[3:0] T5248;
  reg [3:0] counts_866;
  wire[3:0] T11211;
  wire[3:0] T5249;
  wire[3:0] T5250;
  wire T5251;
  wire T5252;
  reg [3:0] counts_867;
  wire[3:0] T11212;
  wire[3:0] T5253;
  wire[3:0] T5254;
  wire T5255;
  wire T5256;
  wire T5257;
  wire T5258;
  wire[3:0] T5259;
  wire[3:0] T5260;
  reg [3:0] counts_868;
  wire[3:0] T11213;
  wire[3:0] T5261;
  wire[3:0] T5262;
  wire T5263;
  wire T5264;
  reg [3:0] counts_869;
  wire[3:0] T11214;
  wire[3:0] T5265;
  wire[3:0] T5266;
  wire T5267;
  wire T5268;
  wire T5269;
  wire[3:0] T5270;
  reg [3:0] counts_870;
  wire[3:0] T11215;
  wire[3:0] T5271;
  wire[3:0] T5272;
  wire T5273;
  wire T5274;
  reg [3:0] counts_871;
  wire[3:0] T11216;
  wire[3:0] T5275;
  wire[3:0] T5276;
  wire T5277;
  wire T5278;
  wire T5279;
  wire T5280;
  wire T5281;
  wire[3:0] T5282;
  wire[3:0] T5283;
  wire[3:0] T5284;
  reg [3:0] counts_872;
  wire[3:0] T11217;
  wire[3:0] T5285;
  wire[3:0] T5286;
  wire T5287;
  wire T5288;
  reg [3:0] counts_873;
  wire[3:0] T11218;
  wire[3:0] T5289;
  wire[3:0] T5290;
  wire T5291;
  wire T5292;
  wire T5293;
  wire[3:0] T5294;
  reg [3:0] counts_874;
  wire[3:0] T11219;
  wire[3:0] T5295;
  wire[3:0] T5296;
  wire T5297;
  wire T5298;
  reg [3:0] counts_875;
  wire[3:0] T11220;
  wire[3:0] T5299;
  wire[3:0] T5300;
  wire T5301;
  wire T5302;
  wire T5303;
  wire T5304;
  wire[3:0] T5305;
  wire[3:0] T5306;
  reg [3:0] counts_876;
  wire[3:0] T11221;
  wire[3:0] T5307;
  wire[3:0] T5308;
  wire T5309;
  wire T5310;
  reg [3:0] counts_877;
  wire[3:0] T11222;
  wire[3:0] T5311;
  wire[3:0] T5312;
  wire T5313;
  wire T5314;
  wire T5315;
  wire[3:0] T5316;
  reg [3:0] counts_878;
  wire[3:0] T11223;
  wire[3:0] T5317;
  wire[3:0] T5318;
  wire T5319;
  wire T5320;
  reg [3:0] counts_879;
  wire[3:0] T11224;
  wire[3:0] T5321;
  wire[3:0] T5322;
  wire T5323;
  wire T5324;
  wire T5325;
  wire T5326;
  wire T5327;
  wire T5328;
  wire[3:0] T5329;
  wire[3:0] T5330;
  wire[3:0] T5331;
  wire[3:0] T5332;
  reg [3:0] counts_880;
  wire[3:0] T11225;
  wire[3:0] T5333;
  wire[3:0] T5334;
  wire T5335;
  wire T5336;
  reg [3:0] counts_881;
  wire[3:0] T11226;
  wire[3:0] T5337;
  wire[3:0] T5338;
  wire T5339;
  wire T5340;
  wire T5341;
  wire[3:0] T5342;
  reg [3:0] counts_882;
  wire[3:0] T11227;
  wire[3:0] T5343;
  wire[3:0] T5344;
  wire T5345;
  wire T5346;
  reg [3:0] counts_883;
  wire[3:0] T11228;
  wire[3:0] T5347;
  wire[3:0] T5348;
  wire T5349;
  wire T5350;
  wire T5351;
  wire T5352;
  wire[3:0] T5353;
  wire[3:0] T5354;
  reg [3:0] counts_884;
  wire[3:0] T11229;
  wire[3:0] T5355;
  wire[3:0] T5356;
  wire T5357;
  wire T5358;
  reg [3:0] counts_885;
  wire[3:0] T11230;
  wire[3:0] T5359;
  wire[3:0] T5360;
  wire T5361;
  wire T5362;
  wire T5363;
  wire[3:0] T5364;
  reg [3:0] counts_886;
  wire[3:0] T11231;
  wire[3:0] T5365;
  wire[3:0] T5366;
  wire T5367;
  wire T5368;
  reg [3:0] counts_887;
  wire[3:0] T11232;
  wire[3:0] T5369;
  wire[3:0] T5370;
  wire T5371;
  wire T5372;
  wire T5373;
  wire T5374;
  wire T5375;
  wire[3:0] T5376;
  wire[3:0] T5377;
  wire[3:0] T5378;
  reg [3:0] counts_888;
  wire[3:0] T11233;
  wire[3:0] T5379;
  wire[3:0] T5380;
  wire T5381;
  wire T5382;
  reg [3:0] counts_889;
  wire[3:0] T11234;
  wire[3:0] T5383;
  wire[3:0] T5384;
  wire T5385;
  wire T5386;
  wire T5387;
  wire[3:0] T5388;
  reg [3:0] counts_890;
  wire[3:0] T11235;
  wire[3:0] T5389;
  wire[3:0] T5390;
  wire T5391;
  wire T5392;
  reg [3:0] counts_891;
  wire[3:0] T11236;
  wire[3:0] T5393;
  wire[3:0] T5394;
  wire T5395;
  wire T5396;
  wire T5397;
  wire T5398;
  wire[3:0] T5399;
  wire[3:0] T5400;
  reg [3:0] counts_892;
  wire[3:0] T11237;
  wire[3:0] T5401;
  wire[3:0] T5402;
  wire T5403;
  wire T5404;
  reg [3:0] counts_893;
  wire[3:0] T11238;
  wire[3:0] T5405;
  wire[3:0] T5406;
  wire T5407;
  wire T5408;
  wire T5409;
  wire[3:0] T5410;
  reg [3:0] counts_894;
  wire[3:0] T11239;
  wire[3:0] T5411;
  wire[3:0] T5412;
  wire T5413;
  wire T5414;
  reg [3:0] counts_895;
  wire[3:0] T11240;
  wire[3:0] T5415;
  wire[3:0] T5416;
  wire T5417;
  wire T5418;
  wire T5419;
  wire T5420;
  wire T5421;
  wire T5422;
  wire T5423;
  wire T5424;
  wire T5425;
  wire[3:0] T5426;
  wire[3:0] T5427;
  wire[3:0] T5428;
  wire[3:0] T5429;
  wire[3:0] T5430;
  wire[3:0] T5431;
  wire[3:0] T5432;
  reg [3:0] counts_896;
  wire[3:0] T11241;
  wire[3:0] T5433;
  wire[3:0] T5434;
  wire T5435;
  wire T5436;
  reg [3:0] counts_897;
  wire[3:0] T11242;
  wire[3:0] T5437;
  wire[3:0] T5438;
  wire T5439;
  wire T5440;
  wire T5441;
  wire[3:0] T5442;
  reg [3:0] counts_898;
  wire[3:0] T11243;
  wire[3:0] T5443;
  wire[3:0] T5444;
  wire T5445;
  wire T5446;
  reg [3:0] counts_899;
  wire[3:0] T11244;
  wire[3:0] T5447;
  wire[3:0] T5448;
  wire T5449;
  wire T5450;
  wire T5451;
  wire T5452;
  wire[3:0] T5453;
  wire[3:0] T5454;
  reg [3:0] counts_900;
  wire[3:0] T11245;
  wire[3:0] T5455;
  wire[3:0] T5456;
  wire T5457;
  wire T5458;
  reg [3:0] counts_901;
  wire[3:0] T11246;
  wire[3:0] T5459;
  wire[3:0] T5460;
  wire T5461;
  wire T5462;
  wire T5463;
  wire[3:0] T5464;
  reg [3:0] counts_902;
  wire[3:0] T11247;
  wire[3:0] T5465;
  wire[3:0] T5466;
  wire T5467;
  wire T5468;
  reg [3:0] counts_903;
  wire[3:0] T11248;
  wire[3:0] T5469;
  wire[3:0] T5470;
  wire T5471;
  wire T5472;
  wire T5473;
  wire T5474;
  wire T5475;
  wire[3:0] T5476;
  wire[3:0] T5477;
  wire[3:0] T5478;
  reg [3:0] counts_904;
  wire[3:0] T11249;
  wire[3:0] T5479;
  wire[3:0] T5480;
  wire T5481;
  wire T5482;
  reg [3:0] counts_905;
  wire[3:0] T11250;
  wire[3:0] T5483;
  wire[3:0] T5484;
  wire T5485;
  wire T5486;
  wire T5487;
  wire[3:0] T5488;
  reg [3:0] counts_906;
  wire[3:0] T11251;
  wire[3:0] T5489;
  wire[3:0] T5490;
  wire T5491;
  wire T5492;
  reg [3:0] counts_907;
  wire[3:0] T11252;
  wire[3:0] T5493;
  wire[3:0] T5494;
  wire T5495;
  wire T5496;
  wire T5497;
  wire T5498;
  wire[3:0] T5499;
  wire[3:0] T5500;
  reg [3:0] counts_908;
  wire[3:0] T11253;
  wire[3:0] T5501;
  wire[3:0] T5502;
  wire T5503;
  wire T5504;
  reg [3:0] counts_909;
  wire[3:0] T11254;
  wire[3:0] T5505;
  wire[3:0] T5506;
  wire T5507;
  wire T5508;
  wire T5509;
  wire[3:0] T5510;
  reg [3:0] counts_910;
  wire[3:0] T11255;
  wire[3:0] T5511;
  wire[3:0] T5512;
  wire T5513;
  wire T5514;
  reg [3:0] counts_911;
  wire[3:0] T11256;
  wire[3:0] T5515;
  wire[3:0] T5516;
  wire T5517;
  wire T5518;
  wire T5519;
  wire T5520;
  wire T5521;
  wire T5522;
  wire[3:0] T5523;
  wire[3:0] T5524;
  wire[3:0] T5525;
  wire[3:0] T5526;
  reg [3:0] counts_912;
  wire[3:0] T11257;
  wire[3:0] T5527;
  wire[3:0] T5528;
  wire T5529;
  wire T5530;
  reg [3:0] counts_913;
  wire[3:0] T11258;
  wire[3:0] T5531;
  wire[3:0] T5532;
  wire T5533;
  wire T5534;
  wire T5535;
  wire[3:0] T5536;
  reg [3:0] counts_914;
  wire[3:0] T11259;
  wire[3:0] T5537;
  wire[3:0] T5538;
  wire T5539;
  wire T5540;
  reg [3:0] counts_915;
  wire[3:0] T11260;
  wire[3:0] T5541;
  wire[3:0] T5542;
  wire T5543;
  wire T5544;
  wire T5545;
  wire T5546;
  wire[3:0] T5547;
  wire[3:0] T5548;
  reg [3:0] counts_916;
  wire[3:0] T11261;
  wire[3:0] T5549;
  wire[3:0] T5550;
  wire T5551;
  wire T5552;
  reg [3:0] counts_917;
  wire[3:0] T11262;
  wire[3:0] T5553;
  wire[3:0] T5554;
  wire T5555;
  wire T5556;
  wire T5557;
  wire[3:0] T5558;
  reg [3:0] counts_918;
  wire[3:0] T11263;
  wire[3:0] T5559;
  wire[3:0] T5560;
  wire T5561;
  wire T5562;
  reg [3:0] counts_919;
  wire[3:0] T11264;
  wire[3:0] T5563;
  wire[3:0] T5564;
  wire T5565;
  wire T5566;
  wire T5567;
  wire T5568;
  wire T5569;
  wire[3:0] T5570;
  wire[3:0] T5571;
  wire[3:0] T5572;
  reg [3:0] counts_920;
  wire[3:0] T11265;
  wire[3:0] T5573;
  wire[3:0] T5574;
  wire T5575;
  wire T5576;
  reg [3:0] counts_921;
  wire[3:0] T11266;
  wire[3:0] T5577;
  wire[3:0] T5578;
  wire T5579;
  wire T5580;
  wire T5581;
  wire[3:0] T5582;
  reg [3:0] counts_922;
  wire[3:0] T11267;
  wire[3:0] T5583;
  wire[3:0] T5584;
  wire T5585;
  wire T5586;
  reg [3:0] counts_923;
  wire[3:0] T11268;
  wire[3:0] T5587;
  wire[3:0] T5588;
  wire T5589;
  wire T5590;
  wire T5591;
  wire T5592;
  wire[3:0] T5593;
  wire[3:0] T5594;
  reg [3:0] counts_924;
  wire[3:0] T11269;
  wire[3:0] T5595;
  wire[3:0] T5596;
  wire T5597;
  wire T5598;
  reg [3:0] counts_925;
  wire[3:0] T11270;
  wire[3:0] T5599;
  wire[3:0] T5600;
  wire T5601;
  wire T5602;
  wire T5603;
  wire[3:0] T5604;
  reg [3:0] counts_926;
  wire[3:0] T11271;
  wire[3:0] T5605;
  wire[3:0] T5606;
  wire T5607;
  wire T5608;
  reg [3:0] counts_927;
  wire[3:0] T11272;
  wire[3:0] T5609;
  wire[3:0] T5610;
  wire T5611;
  wire T5612;
  wire T5613;
  wire T5614;
  wire T5615;
  wire T5616;
  wire T5617;
  wire[3:0] T5618;
  wire[3:0] T5619;
  wire[3:0] T5620;
  wire[3:0] T5621;
  wire[3:0] T5622;
  reg [3:0] counts_928;
  wire[3:0] T11273;
  wire[3:0] T5623;
  wire[3:0] T5624;
  wire T5625;
  wire T5626;
  reg [3:0] counts_929;
  wire[3:0] T11274;
  wire[3:0] T5627;
  wire[3:0] T5628;
  wire T5629;
  wire T5630;
  wire T5631;
  wire[3:0] T5632;
  reg [3:0] counts_930;
  wire[3:0] T11275;
  wire[3:0] T5633;
  wire[3:0] T5634;
  wire T5635;
  wire T5636;
  reg [3:0] counts_931;
  wire[3:0] T11276;
  wire[3:0] T5637;
  wire[3:0] T5638;
  wire T5639;
  wire T5640;
  wire T5641;
  wire T5642;
  wire[3:0] T5643;
  wire[3:0] T5644;
  reg [3:0] counts_932;
  wire[3:0] T11277;
  wire[3:0] T5645;
  wire[3:0] T5646;
  wire T5647;
  wire T5648;
  reg [3:0] counts_933;
  wire[3:0] T11278;
  wire[3:0] T5649;
  wire[3:0] T5650;
  wire T5651;
  wire T5652;
  wire T5653;
  wire[3:0] T5654;
  reg [3:0] counts_934;
  wire[3:0] T11279;
  wire[3:0] T5655;
  wire[3:0] T5656;
  wire T5657;
  wire T5658;
  reg [3:0] counts_935;
  wire[3:0] T11280;
  wire[3:0] T5659;
  wire[3:0] T5660;
  wire T5661;
  wire T5662;
  wire T5663;
  wire T5664;
  wire T5665;
  wire[3:0] T5666;
  wire[3:0] T5667;
  wire[3:0] T5668;
  reg [3:0] counts_936;
  wire[3:0] T11281;
  wire[3:0] T5669;
  wire[3:0] T5670;
  wire T5671;
  wire T5672;
  reg [3:0] counts_937;
  wire[3:0] T11282;
  wire[3:0] T5673;
  wire[3:0] T5674;
  wire T5675;
  wire T5676;
  wire T5677;
  wire[3:0] T5678;
  reg [3:0] counts_938;
  wire[3:0] T11283;
  wire[3:0] T5679;
  wire[3:0] T5680;
  wire T5681;
  wire T5682;
  reg [3:0] counts_939;
  wire[3:0] T11284;
  wire[3:0] T5683;
  wire[3:0] T5684;
  wire T5685;
  wire T5686;
  wire T5687;
  wire T5688;
  wire[3:0] T5689;
  wire[3:0] T5690;
  reg [3:0] counts_940;
  wire[3:0] T11285;
  wire[3:0] T5691;
  wire[3:0] T5692;
  wire T5693;
  wire T5694;
  reg [3:0] counts_941;
  wire[3:0] T11286;
  wire[3:0] T5695;
  wire[3:0] T5696;
  wire T5697;
  wire T5698;
  wire T5699;
  wire[3:0] T5700;
  reg [3:0] counts_942;
  wire[3:0] T11287;
  wire[3:0] T5701;
  wire[3:0] T5702;
  wire T5703;
  wire T5704;
  reg [3:0] counts_943;
  wire[3:0] T11288;
  wire[3:0] T5705;
  wire[3:0] T5706;
  wire T5707;
  wire T5708;
  wire T5709;
  wire T5710;
  wire T5711;
  wire T5712;
  wire[3:0] T5713;
  wire[3:0] T5714;
  wire[3:0] T5715;
  wire[3:0] T5716;
  reg [3:0] counts_944;
  wire[3:0] T11289;
  wire[3:0] T5717;
  wire[3:0] T5718;
  wire T5719;
  wire T5720;
  reg [3:0] counts_945;
  wire[3:0] T11290;
  wire[3:0] T5721;
  wire[3:0] T5722;
  wire T5723;
  wire T5724;
  wire T5725;
  wire[3:0] T5726;
  reg [3:0] counts_946;
  wire[3:0] T11291;
  wire[3:0] T5727;
  wire[3:0] T5728;
  wire T5729;
  wire T5730;
  reg [3:0] counts_947;
  wire[3:0] T11292;
  wire[3:0] T5731;
  wire[3:0] T5732;
  wire T5733;
  wire T5734;
  wire T5735;
  wire T5736;
  wire[3:0] T5737;
  wire[3:0] T5738;
  reg [3:0] counts_948;
  wire[3:0] T11293;
  wire[3:0] T5739;
  wire[3:0] T5740;
  wire T5741;
  wire T5742;
  reg [3:0] counts_949;
  wire[3:0] T11294;
  wire[3:0] T5743;
  wire[3:0] T5744;
  wire T5745;
  wire T5746;
  wire T5747;
  wire[3:0] T5748;
  reg [3:0] counts_950;
  wire[3:0] T11295;
  wire[3:0] T5749;
  wire[3:0] T5750;
  wire T5751;
  wire T5752;
  reg [3:0] counts_951;
  wire[3:0] T11296;
  wire[3:0] T5753;
  wire[3:0] T5754;
  wire T5755;
  wire T5756;
  wire T5757;
  wire T5758;
  wire T5759;
  wire[3:0] T5760;
  wire[3:0] T5761;
  wire[3:0] T5762;
  reg [3:0] counts_952;
  wire[3:0] T11297;
  wire[3:0] T5763;
  wire[3:0] T5764;
  wire T5765;
  wire T5766;
  reg [3:0] counts_953;
  wire[3:0] T11298;
  wire[3:0] T5767;
  wire[3:0] T5768;
  wire T5769;
  wire T5770;
  wire T5771;
  wire[3:0] T5772;
  reg [3:0] counts_954;
  wire[3:0] T11299;
  wire[3:0] T5773;
  wire[3:0] T5774;
  wire T5775;
  wire T5776;
  reg [3:0] counts_955;
  wire[3:0] T11300;
  wire[3:0] T5777;
  wire[3:0] T5778;
  wire T5779;
  wire T5780;
  wire T5781;
  wire T5782;
  wire[3:0] T5783;
  wire[3:0] T5784;
  reg [3:0] counts_956;
  wire[3:0] T11301;
  wire[3:0] T5785;
  wire[3:0] T5786;
  wire T5787;
  wire T5788;
  reg [3:0] counts_957;
  wire[3:0] T11302;
  wire[3:0] T5789;
  wire[3:0] T5790;
  wire T5791;
  wire T5792;
  wire T5793;
  wire[3:0] T5794;
  reg [3:0] counts_958;
  wire[3:0] T11303;
  wire[3:0] T5795;
  wire[3:0] T5796;
  wire T5797;
  wire T5798;
  reg [3:0] counts_959;
  wire[3:0] T11304;
  wire[3:0] T5799;
  wire[3:0] T5800;
  wire T5801;
  wire T5802;
  wire T5803;
  wire T5804;
  wire T5805;
  wire T5806;
  wire T5807;
  wire T5808;
  wire[3:0] T5809;
  wire[3:0] T5810;
  wire[3:0] T5811;
  wire[3:0] T5812;
  wire[3:0] T5813;
  wire[3:0] T5814;
  reg [3:0] counts_960;
  wire[3:0] T11305;
  wire[3:0] T5815;
  wire[3:0] T5816;
  wire T5817;
  wire T5818;
  reg [3:0] counts_961;
  wire[3:0] T11306;
  wire[3:0] T5819;
  wire[3:0] T5820;
  wire T5821;
  wire T5822;
  wire T5823;
  wire[3:0] T5824;
  reg [3:0] counts_962;
  wire[3:0] T11307;
  wire[3:0] T5825;
  wire[3:0] T5826;
  wire T5827;
  wire T5828;
  reg [3:0] counts_963;
  wire[3:0] T11308;
  wire[3:0] T5829;
  wire[3:0] T5830;
  wire T5831;
  wire T5832;
  wire T5833;
  wire T5834;
  wire[3:0] T5835;
  wire[3:0] T5836;
  reg [3:0] counts_964;
  wire[3:0] T11309;
  wire[3:0] T5837;
  wire[3:0] T5838;
  wire T5839;
  wire T5840;
  reg [3:0] counts_965;
  wire[3:0] T11310;
  wire[3:0] T5841;
  wire[3:0] T5842;
  wire T5843;
  wire T5844;
  wire T5845;
  wire[3:0] T5846;
  reg [3:0] counts_966;
  wire[3:0] T11311;
  wire[3:0] T5847;
  wire[3:0] T5848;
  wire T5849;
  wire T5850;
  reg [3:0] counts_967;
  wire[3:0] T11312;
  wire[3:0] T5851;
  wire[3:0] T5852;
  wire T5853;
  wire T5854;
  wire T5855;
  wire T5856;
  wire T5857;
  wire[3:0] T5858;
  wire[3:0] T5859;
  wire[3:0] T5860;
  reg [3:0] counts_968;
  wire[3:0] T11313;
  wire[3:0] T5861;
  wire[3:0] T5862;
  wire T5863;
  wire T5864;
  reg [3:0] counts_969;
  wire[3:0] T11314;
  wire[3:0] T5865;
  wire[3:0] T5866;
  wire T5867;
  wire T5868;
  wire T5869;
  wire[3:0] T5870;
  reg [3:0] counts_970;
  wire[3:0] T11315;
  wire[3:0] T5871;
  wire[3:0] T5872;
  wire T5873;
  wire T5874;
  reg [3:0] counts_971;
  wire[3:0] T11316;
  wire[3:0] T5875;
  wire[3:0] T5876;
  wire T5877;
  wire T5878;
  wire T5879;
  wire T5880;
  wire[3:0] T5881;
  wire[3:0] T5882;
  reg [3:0] counts_972;
  wire[3:0] T11317;
  wire[3:0] T5883;
  wire[3:0] T5884;
  wire T5885;
  wire T5886;
  reg [3:0] counts_973;
  wire[3:0] T11318;
  wire[3:0] T5887;
  wire[3:0] T5888;
  wire T5889;
  wire T5890;
  wire T5891;
  wire[3:0] T5892;
  reg [3:0] counts_974;
  wire[3:0] T11319;
  wire[3:0] T5893;
  wire[3:0] T5894;
  wire T5895;
  wire T5896;
  reg [3:0] counts_975;
  wire[3:0] T11320;
  wire[3:0] T5897;
  wire[3:0] T5898;
  wire T5899;
  wire T5900;
  wire T5901;
  wire T5902;
  wire T5903;
  wire T5904;
  wire[3:0] T5905;
  wire[3:0] T5906;
  wire[3:0] T5907;
  wire[3:0] T5908;
  reg [3:0] counts_976;
  wire[3:0] T11321;
  wire[3:0] T5909;
  wire[3:0] T5910;
  wire T5911;
  wire T5912;
  reg [3:0] counts_977;
  wire[3:0] T11322;
  wire[3:0] T5913;
  wire[3:0] T5914;
  wire T5915;
  wire T5916;
  wire T5917;
  wire[3:0] T5918;
  reg [3:0] counts_978;
  wire[3:0] T11323;
  wire[3:0] T5919;
  wire[3:0] T5920;
  wire T5921;
  wire T5922;
  reg [3:0] counts_979;
  wire[3:0] T11324;
  wire[3:0] T5923;
  wire[3:0] T5924;
  wire T5925;
  wire T5926;
  wire T5927;
  wire T5928;
  wire[3:0] T5929;
  wire[3:0] T5930;
  reg [3:0] counts_980;
  wire[3:0] T11325;
  wire[3:0] T5931;
  wire[3:0] T5932;
  wire T5933;
  wire T5934;
  reg [3:0] counts_981;
  wire[3:0] T11326;
  wire[3:0] T5935;
  wire[3:0] T5936;
  wire T5937;
  wire T5938;
  wire T5939;
  wire[3:0] T5940;
  reg [3:0] counts_982;
  wire[3:0] T11327;
  wire[3:0] T5941;
  wire[3:0] T5942;
  wire T5943;
  wire T5944;
  reg [3:0] counts_983;
  wire[3:0] T11328;
  wire[3:0] T5945;
  wire[3:0] T5946;
  wire T5947;
  wire T5948;
  wire T5949;
  wire T5950;
  wire T5951;
  wire[3:0] T5952;
  wire[3:0] T5953;
  wire[3:0] T5954;
  reg [3:0] counts_984;
  wire[3:0] T11329;
  wire[3:0] T5955;
  wire[3:0] T5956;
  wire T5957;
  wire T5958;
  reg [3:0] counts_985;
  wire[3:0] T11330;
  wire[3:0] T5959;
  wire[3:0] T5960;
  wire T5961;
  wire T5962;
  wire T5963;
  wire[3:0] T5964;
  reg [3:0] counts_986;
  wire[3:0] T11331;
  wire[3:0] T5965;
  wire[3:0] T5966;
  wire T5967;
  wire T5968;
  reg [3:0] counts_987;
  wire[3:0] T11332;
  wire[3:0] T5969;
  wire[3:0] T5970;
  wire T5971;
  wire T5972;
  wire T5973;
  wire T5974;
  wire[3:0] T5975;
  wire[3:0] T5976;
  reg [3:0] counts_988;
  wire[3:0] T11333;
  wire[3:0] T5977;
  wire[3:0] T5978;
  wire T5979;
  wire T5980;
  reg [3:0] counts_989;
  wire[3:0] T11334;
  wire[3:0] T5981;
  wire[3:0] T5982;
  wire T5983;
  wire T5984;
  wire T5985;
  wire[3:0] T5986;
  reg [3:0] counts_990;
  wire[3:0] T11335;
  wire[3:0] T5987;
  wire[3:0] T5988;
  wire T5989;
  wire T5990;
  reg [3:0] counts_991;
  wire[3:0] T11336;
  wire[3:0] T5991;
  wire[3:0] T5992;
  wire T5993;
  wire T5994;
  wire T5995;
  wire T5996;
  wire T5997;
  wire T5998;
  wire T5999;
  wire[3:0] T6000;
  wire[3:0] T6001;
  wire[3:0] T6002;
  wire[3:0] T6003;
  wire[3:0] T6004;
  reg [3:0] counts_992;
  wire[3:0] T11337;
  wire[3:0] T6005;
  wire[3:0] T6006;
  wire T6007;
  wire T6008;
  reg [3:0] counts_993;
  wire[3:0] T11338;
  wire[3:0] T6009;
  wire[3:0] T6010;
  wire T6011;
  wire T6012;
  wire T6013;
  wire[3:0] T6014;
  reg [3:0] counts_994;
  wire[3:0] T11339;
  wire[3:0] T6015;
  wire[3:0] T6016;
  wire T6017;
  wire T6018;
  reg [3:0] counts_995;
  wire[3:0] T11340;
  wire[3:0] T6019;
  wire[3:0] T6020;
  wire T6021;
  wire T6022;
  wire T6023;
  wire T6024;
  wire[3:0] T6025;
  wire[3:0] T6026;
  reg [3:0] counts_996;
  wire[3:0] T11341;
  wire[3:0] T6027;
  wire[3:0] T6028;
  wire T6029;
  wire T6030;
  reg [3:0] counts_997;
  wire[3:0] T11342;
  wire[3:0] T6031;
  wire[3:0] T6032;
  wire T6033;
  wire T6034;
  wire T6035;
  wire[3:0] T6036;
  reg [3:0] counts_998;
  wire[3:0] T11343;
  wire[3:0] T6037;
  wire[3:0] T6038;
  wire T6039;
  wire T6040;
  reg [3:0] counts_999;
  wire[3:0] T11344;
  wire[3:0] T6041;
  wire[3:0] T6042;
  wire T6043;
  wire T6044;
  wire T6045;
  wire T6046;
  wire T6047;
  wire[3:0] T6048;
  wire[3:0] T6049;
  wire[3:0] T6050;
  reg [3:0] counts_1000;
  wire[3:0] T11345;
  wire[3:0] T6051;
  wire[3:0] T6052;
  wire T6053;
  wire T6054;
  reg [3:0] counts_1001;
  wire[3:0] T11346;
  wire[3:0] T6055;
  wire[3:0] T6056;
  wire T6057;
  wire T6058;
  wire T6059;
  wire[3:0] T6060;
  reg [3:0] counts_1002;
  wire[3:0] T11347;
  wire[3:0] T6061;
  wire[3:0] T6062;
  wire T6063;
  wire T6064;
  reg [3:0] counts_1003;
  wire[3:0] T11348;
  wire[3:0] T6065;
  wire[3:0] T6066;
  wire T6067;
  wire T6068;
  wire T6069;
  wire T6070;
  wire[3:0] T6071;
  wire[3:0] T6072;
  reg [3:0] counts_1004;
  wire[3:0] T11349;
  wire[3:0] T6073;
  wire[3:0] T6074;
  wire T6075;
  wire T6076;
  reg [3:0] counts_1005;
  wire[3:0] T11350;
  wire[3:0] T6077;
  wire[3:0] T6078;
  wire T6079;
  wire T6080;
  wire T6081;
  wire[3:0] T6082;
  reg [3:0] counts_1006;
  wire[3:0] T11351;
  wire[3:0] T6083;
  wire[3:0] T6084;
  wire T6085;
  wire T6086;
  reg [3:0] counts_1007;
  wire[3:0] T11352;
  wire[3:0] T6087;
  wire[3:0] T6088;
  wire T6089;
  wire T6090;
  wire T6091;
  wire T6092;
  wire T6093;
  wire T6094;
  wire[3:0] T6095;
  wire[3:0] T6096;
  wire[3:0] T6097;
  wire[3:0] T6098;
  reg [3:0] counts_1008;
  wire[3:0] T11353;
  wire[3:0] T6099;
  wire[3:0] T6100;
  wire T6101;
  wire T6102;
  reg [3:0] counts_1009;
  wire[3:0] T11354;
  wire[3:0] T6103;
  wire[3:0] T6104;
  wire T6105;
  wire T6106;
  wire T6107;
  wire[3:0] T6108;
  reg [3:0] counts_1010;
  wire[3:0] T11355;
  wire[3:0] T6109;
  wire[3:0] T6110;
  wire T6111;
  wire T6112;
  reg [3:0] counts_1011;
  wire[3:0] T11356;
  wire[3:0] T6113;
  wire[3:0] T6114;
  wire T6115;
  wire T6116;
  wire T6117;
  wire T6118;
  wire[3:0] T6119;
  wire[3:0] T6120;
  reg [3:0] counts_1012;
  wire[3:0] T11357;
  wire[3:0] T6121;
  wire[3:0] T6122;
  wire T6123;
  wire T6124;
  reg [3:0] counts_1013;
  wire[3:0] T11358;
  wire[3:0] T6125;
  wire[3:0] T6126;
  wire T6127;
  wire T6128;
  wire T6129;
  wire[3:0] T6130;
  reg [3:0] counts_1014;
  wire[3:0] T11359;
  wire[3:0] T6131;
  wire[3:0] T6132;
  wire T6133;
  wire T6134;
  reg [3:0] counts_1015;
  wire[3:0] T11360;
  wire[3:0] T6135;
  wire[3:0] T6136;
  wire T6137;
  wire T6138;
  wire T6139;
  wire T6140;
  wire T6141;
  wire[3:0] T6142;
  wire[3:0] T6143;
  wire[3:0] T6144;
  reg [3:0] counts_1016;
  wire[3:0] T11361;
  wire[3:0] T6145;
  wire[3:0] T6146;
  wire T6147;
  wire T6148;
  reg [3:0] counts_1017;
  wire[3:0] T11362;
  wire[3:0] T6149;
  wire[3:0] T6150;
  wire T6151;
  wire T6152;
  wire T6153;
  wire[3:0] T6154;
  reg [3:0] counts_1018;
  wire[3:0] T11363;
  wire[3:0] T6155;
  wire[3:0] T6156;
  wire T6157;
  wire T6158;
  reg [3:0] counts_1019;
  wire[3:0] T11364;
  wire[3:0] T6159;
  wire[3:0] T6160;
  wire T6161;
  wire T6162;
  wire T6163;
  wire T6164;
  wire[3:0] T6165;
  wire[3:0] T6166;
  reg [3:0] counts_1020;
  wire[3:0] T11365;
  wire[3:0] T6167;
  wire[3:0] T6168;
  wire T6169;
  wire T6170;
  reg [3:0] counts_1021;
  wire[3:0] T11366;
  wire[3:0] T6171;
  wire[3:0] T6172;
  wire T6173;
  wire T6174;
  wire T6175;
  wire[3:0] T6176;
  reg [3:0] counts_1022;
  wire[3:0] T11367;
  wire[3:0] T6177;
  wire[3:0] T6178;
  wire T6179;
  wire T6180;
  reg [3:0] counts_1023;
  wire[3:0] T11368;
  wire[3:0] T6181;
  wire[3:0] T6182;
  wire T6183;
  wire T6184;
  wire T6185;
  wire T6186;
  wire T6187;
  wire T6188;
  wire T6189;
  wire T6190;
  wire T6191;
  wire T6192;
  wire T6193;
  wire T6194;
  wire[3:0] T6195;
  wire T6196;
  wire T6197;
  reg [3:0] counts_1;
  wire[3:0] T11369;
  wire[3:0] T6198;
  wire[3:0] T6199;
  wire T6200;
  wire T6201;
  wire T6202;
  wire[9:0] T6203;
  wire[3:0] T6204;
  wire T6205;
  wire T6206;
  wire[3:0] T6207;
  wire[3:0] T6208;
  wire T6209;
  wire[3:0] T6210;
  wire T6211;
  wire T6212;
  wire T6213;
  wire[3:0] T6214;
  wire[3:0] T6215;
  wire[3:0] T6216;
  wire T6217;
  wire[3:0] T6218;
  wire T6219;
  wire T6220;
  wire[3:0] T6221;
  wire[3:0] T6222;
  wire T6223;
  wire[3:0] T6224;
  wire T6225;
  wire T6226;
  wire T6227;
  wire T6228;
  wire[3:0] T6229;
  wire[3:0] T6230;
  wire[3:0] T6231;
  wire[3:0] T6232;
  wire T6233;
  wire[3:0] T6234;
  wire T6235;
  wire T6236;
  wire[3:0] T6237;
  wire[3:0] T6238;
  wire T6239;
  wire[3:0] T6240;
  wire T6241;
  wire T6242;
  wire T6243;
  wire[3:0] T6244;
  wire[3:0] T6245;
  wire[3:0] T6246;
  wire T6247;
  wire[3:0] T6248;
  wire T6249;
  wire T6250;
  wire[3:0] T6251;
  wire[3:0] T6252;
  wire T6253;
  wire[3:0] T6254;
  wire T6255;
  wire T6256;
  wire T6257;
  wire T6258;
  wire T6259;
  wire[3:0] T6260;
  wire[3:0] T6261;
  wire[3:0] T6262;
  wire[3:0] T6263;
  wire[3:0] T6264;
  wire T6265;
  wire[3:0] T6266;
  wire T6267;
  wire T6268;
  wire[3:0] T6269;
  wire[3:0] T6270;
  wire T6271;
  wire[3:0] T6272;
  wire T6273;
  wire T6274;
  wire T6275;
  wire[3:0] T6276;
  wire[3:0] T6277;
  wire[3:0] T6278;
  wire T6279;
  wire[3:0] T6280;
  wire T6281;
  wire T6282;
  wire[3:0] T6283;
  wire[3:0] T6284;
  wire T6285;
  wire[3:0] T6286;
  wire T6287;
  wire T6288;
  wire T6289;
  wire T6290;
  wire[3:0] T6291;
  wire[3:0] T6292;
  wire[3:0] T6293;
  wire[3:0] T6294;
  wire T6295;
  wire[3:0] T6296;
  wire T6297;
  wire T6298;
  wire[3:0] T6299;
  wire[3:0] T6300;
  wire T6301;
  wire[3:0] T6302;
  wire T6303;
  wire T6304;
  wire T6305;
  wire[3:0] T6306;
  wire[3:0] T6307;
  wire[3:0] T6308;
  wire T6309;
  wire[3:0] T6310;
  wire T6311;
  wire T6312;
  wire[3:0] T6313;
  wire[3:0] T6314;
  wire T6315;
  wire[3:0] T6316;
  wire T6317;
  wire T6318;
  wire T6319;
  wire T6320;
  wire T6321;
  wire T6322;
  wire[3:0] T6323;
  wire[3:0] T6324;
  wire[3:0] T6325;
  wire[3:0] T6326;
  wire[3:0] T6327;
  wire[3:0] T6328;
  wire T6329;
  wire[3:0] T6330;
  wire T6331;
  wire T6332;
  wire[3:0] T6333;
  wire[3:0] T6334;
  wire T6335;
  wire[3:0] T6336;
  wire T6337;
  wire T6338;
  wire T6339;
  wire[3:0] T6340;
  wire[3:0] T6341;
  wire[3:0] T6342;
  wire T6343;
  wire[3:0] T6344;
  wire T6345;
  wire T6346;
  wire[3:0] T6347;
  wire[3:0] T6348;
  wire T6349;
  wire[3:0] T6350;
  wire T6351;
  wire T6352;
  wire T6353;
  wire T6354;
  wire[3:0] T6355;
  wire[3:0] T6356;
  wire[3:0] T6357;
  wire[3:0] T6358;
  wire T6359;
  wire[3:0] T6360;
  wire T6361;
  wire T6362;
  wire[3:0] T6363;
  wire[3:0] T6364;
  wire T6365;
  wire[3:0] T6366;
  wire T6367;
  wire T6368;
  wire T6369;
  wire[3:0] T6370;
  wire[3:0] T6371;
  wire[3:0] T6372;
  wire T6373;
  wire[3:0] T6374;
  wire T6375;
  wire T6376;
  wire[3:0] T6377;
  wire[3:0] T6378;
  wire T6379;
  wire[3:0] T6380;
  wire T6381;
  wire T6382;
  wire T6383;
  wire T6384;
  wire T6385;
  wire[3:0] T6386;
  wire[3:0] T6387;
  wire[3:0] T6388;
  wire[3:0] T6389;
  wire[3:0] T6390;
  wire T6391;
  wire[3:0] T6392;
  wire T6393;
  wire T6394;
  wire[3:0] T6395;
  wire[3:0] T6396;
  wire T6397;
  wire[3:0] T6398;
  wire T6399;
  wire T6400;
  wire T6401;
  wire[3:0] T6402;
  wire[3:0] T6403;
  wire[3:0] T6404;
  wire T6405;
  wire[3:0] T6406;
  wire T6407;
  wire T6408;
  wire[3:0] T6409;
  wire[3:0] T6410;
  wire T6411;
  wire[3:0] T6412;
  wire T6413;
  wire T6414;
  wire T6415;
  wire T6416;
  wire[3:0] T6417;
  wire[3:0] T6418;
  wire[3:0] T6419;
  wire[3:0] T6420;
  wire T6421;
  wire[3:0] T6422;
  wire T6423;
  wire T6424;
  wire[3:0] T6425;
  wire[3:0] T6426;
  wire T6427;
  wire[3:0] T6428;
  wire T6429;
  wire T6430;
  wire T6431;
  wire[3:0] T6432;
  wire[3:0] T6433;
  wire[3:0] T6434;
  wire T6435;
  wire[3:0] T6436;
  wire T6437;
  wire T6438;
  wire[3:0] T6439;
  wire[3:0] T6440;
  wire T6441;
  wire[3:0] T6442;
  wire T6443;
  wire T6444;
  wire T6445;
  wire T6446;
  wire T6447;
  wire T6448;
  wire T6449;
  wire[3:0] T6450;
  wire[3:0] T6451;
  wire[3:0] T6452;
  wire[3:0] T6453;
  wire[3:0] T6454;
  wire[3:0] T6455;
  wire[3:0] T6456;
  wire T6457;
  wire[3:0] T6458;
  wire T6459;
  wire T6460;
  wire[3:0] T6461;
  wire[3:0] T6462;
  wire T6463;
  wire[3:0] T6464;
  wire T6465;
  wire T6466;
  wire T6467;
  wire[3:0] T6468;
  wire[3:0] T6469;
  wire[3:0] T6470;
  wire T6471;
  wire[3:0] T6472;
  wire T6473;
  wire T6474;
  wire[3:0] T6475;
  wire[3:0] T6476;
  wire T6477;
  wire[3:0] T6478;
  wire T6479;
  wire T6480;
  wire T6481;
  wire T6482;
  wire[3:0] T6483;
  wire[3:0] T6484;
  wire[3:0] T6485;
  wire[3:0] T6486;
  wire T6487;
  wire[3:0] T6488;
  wire T6489;
  wire T6490;
  wire[3:0] T6491;
  wire[3:0] T6492;
  wire T6493;
  wire[3:0] T6494;
  wire T6495;
  wire T6496;
  wire T6497;
  wire[3:0] T6498;
  wire[3:0] T6499;
  wire[3:0] T6500;
  wire T6501;
  wire[3:0] T6502;
  wire T6503;
  wire T6504;
  wire[3:0] T6505;
  wire[3:0] T6506;
  wire T6507;
  wire[3:0] T6508;
  wire T6509;
  wire T6510;
  wire T6511;
  wire T6512;
  wire T6513;
  wire[3:0] T6514;
  wire[3:0] T6515;
  wire[3:0] T6516;
  wire[3:0] T6517;
  wire[3:0] T6518;
  wire T6519;
  wire[3:0] T6520;
  wire T6521;
  wire T6522;
  wire[3:0] T6523;
  wire[3:0] T6524;
  wire T6525;
  wire[3:0] T6526;
  wire T6527;
  wire T6528;
  wire T6529;
  wire[3:0] T6530;
  wire[3:0] T6531;
  wire[3:0] T6532;
  wire T6533;
  wire[3:0] T6534;
  wire T6535;
  wire T6536;
  wire[3:0] T6537;
  wire[3:0] T6538;
  wire T6539;
  wire[3:0] T6540;
  wire T6541;
  wire T6542;
  wire T6543;
  wire T6544;
  wire[3:0] T6545;
  wire[3:0] T6546;
  wire[3:0] T6547;
  wire[3:0] T6548;
  wire T6549;
  wire[3:0] T6550;
  wire T6551;
  wire T6552;
  wire[3:0] T6553;
  wire[3:0] T6554;
  wire T6555;
  wire[3:0] T6556;
  wire T6557;
  wire T6558;
  wire T6559;
  wire[3:0] T6560;
  wire[3:0] T6561;
  wire[3:0] T6562;
  wire T6563;
  wire[3:0] T6564;
  wire T6565;
  wire T6566;
  wire[3:0] T6567;
  wire[3:0] T6568;
  wire T6569;
  wire[3:0] T6570;
  wire T6571;
  wire T6572;
  wire T6573;
  wire T6574;
  wire T6575;
  wire T6576;
  wire[3:0] T6577;
  wire[3:0] T6578;
  wire[3:0] T6579;
  wire[3:0] T6580;
  wire[3:0] T6581;
  wire[3:0] T6582;
  wire T6583;
  wire[3:0] T6584;
  wire T6585;
  wire T6586;
  wire[3:0] T6587;
  wire[3:0] T6588;
  wire T6589;
  wire[3:0] T6590;
  wire T6591;
  wire T6592;
  wire T6593;
  wire[3:0] T6594;
  wire[3:0] T6595;
  wire[3:0] T6596;
  wire T6597;
  wire[3:0] T6598;
  wire T6599;
  wire T6600;
  wire[3:0] T6601;
  wire[3:0] T6602;
  wire T6603;
  wire[3:0] T6604;
  wire T6605;
  wire T6606;
  wire T6607;
  wire T6608;
  wire[3:0] T6609;
  wire[3:0] T6610;
  wire[3:0] T6611;
  wire[3:0] T6612;
  wire T6613;
  wire[3:0] T6614;
  wire T6615;
  wire T6616;
  wire[3:0] T6617;
  wire[3:0] T6618;
  wire T6619;
  wire[3:0] T6620;
  wire T6621;
  wire T6622;
  wire T6623;
  wire[3:0] T6624;
  wire[3:0] T6625;
  wire[3:0] T6626;
  wire T6627;
  wire[3:0] T6628;
  wire T6629;
  wire T6630;
  wire[3:0] T6631;
  wire[3:0] T6632;
  wire T6633;
  wire[3:0] T6634;
  wire T6635;
  wire T6636;
  wire T6637;
  wire T6638;
  wire T6639;
  wire[3:0] T6640;
  wire[3:0] T6641;
  wire[3:0] T6642;
  wire[3:0] T6643;
  wire[3:0] T6644;
  wire T6645;
  wire[3:0] T6646;
  wire T6647;
  wire T6648;
  wire[3:0] T6649;
  wire[3:0] T6650;
  wire T6651;
  wire[3:0] T6652;
  wire T6653;
  wire T6654;
  wire T6655;
  wire[3:0] T6656;
  wire[3:0] T6657;
  wire[3:0] T6658;
  wire T6659;
  wire[3:0] T6660;
  wire T6661;
  wire T6662;
  wire[3:0] T6663;
  wire[3:0] T6664;
  wire T6665;
  wire[3:0] T6666;
  wire T6667;
  wire T6668;
  wire T6669;
  wire T6670;
  wire[3:0] T6671;
  wire[3:0] T6672;
  wire[3:0] T6673;
  wire[3:0] T6674;
  wire T6675;
  wire[3:0] T6676;
  wire T6677;
  wire T6678;
  wire[3:0] T6679;
  wire[3:0] T6680;
  wire T6681;
  wire[3:0] T6682;
  wire T6683;
  wire T6684;
  wire T6685;
  wire[3:0] T6686;
  wire[3:0] T6687;
  wire[3:0] T6688;
  wire T6689;
  wire[3:0] T6690;
  wire T6691;
  wire T6692;
  wire[3:0] T6693;
  wire[3:0] T6694;
  wire T6695;
  wire[3:0] T6696;
  wire T6697;
  wire T6698;
  wire T6699;
  wire T6700;
  wire T6701;
  wire T6702;
  wire T6703;
  wire T6704;
  wire[3:0] T6705;
  wire[3:0] T6706;
  wire[3:0] T6707;
  wire[3:0] T6708;
  wire[3:0] T6709;
  wire[3:0] T6710;
  wire[3:0] T6711;
  wire[3:0] T6712;
  wire T6713;
  wire[3:0] T6714;
  wire T6715;
  wire T6716;
  wire[3:0] T6717;
  wire[3:0] T6718;
  wire T6719;
  wire[3:0] T6720;
  wire T6721;
  wire T6722;
  wire T6723;
  wire[3:0] T6724;
  wire[3:0] T6725;
  wire[3:0] T6726;
  wire T6727;
  wire[3:0] T6728;
  wire T6729;
  wire T6730;
  wire[3:0] T6731;
  wire[3:0] T6732;
  wire T6733;
  wire[3:0] T6734;
  wire T6735;
  wire T6736;
  wire T6737;
  wire T6738;
  wire[3:0] T6739;
  wire[3:0] T6740;
  wire[3:0] T6741;
  wire[3:0] T6742;
  wire T6743;
  wire[3:0] T6744;
  wire T6745;
  wire T6746;
  wire[3:0] T6747;
  wire[3:0] T6748;
  wire T6749;
  wire[3:0] T6750;
  wire T6751;
  wire T6752;
  wire T6753;
  wire[3:0] T6754;
  wire[3:0] T6755;
  wire[3:0] T6756;
  wire T6757;
  wire[3:0] T6758;
  wire T6759;
  wire T6760;
  wire[3:0] T6761;
  wire[3:0] T6762;
  wire T6763;
  wire[3:0] T6764;
  wire T6765;
  wire T6766;
  wire T6767;
  wire T6768;
  wire T6769;
  wire[3:0] T6770;
  wire[3:0] T6771;
  wire[3:0] T6772;
  wire[3:0] T6773;
  wire[3:0] T6774;
  wire T6775;
  wire[3:0] T6776;
  wire T6777;
  wire T6778;
  wire[3:0] T6779;
  wire[3:0] T6780;
  wire T6781;
  wire[3:0] T6782;
  wire T6783;
  wire T6784;
  wire T6785;
  wire[3:0] T6786;
  wire[3:0] T6787;
  wire[3:0] T6788;
  wire T6789;
  wire[3:0] T6790;
  wire T6791;
  wire T6792;
  wire[3:0] T6793;
  wire[3:0] T6794;
  wire T6795;
  wire[3:0] T6796;
  wire T6797;
  wire T6798;
  wire T6799;
  wire T6800;
  wire[3:0] T6801;
  wire[3:0] T6802;
  wire[3:0] T6803;
  wire[3:0] T6804;
  wire T6805;
  wire[3:0] T6806;
  wire T6807;
  wire T6808;
  wire[3:0] T6809;
  wire[3:0] T6810;
  wire T6811;
  wire[3:0] T6812;
  wire T6813;
  wire T6814;
  wire T6815;
  wire[3:0] T6816;
  wire[3:0] T6817;
  wire[3:0] T6818;
  wire T6819;
  wire[3:0] T6820;
  wire T6821;
  wire T6822;
  wire[3:0] T6823;
  wire[3:0] T6824;
  wire T6825;
  wire[3:0] T6826;
  wire T6827;
  wire T6828;
  wire T6829;
  wire T6830;
  wire T6831;
  wire T6832;
  wire[3:0] T6833;
  wire[3:0] T6834;
  wire[3:0] T6835;
  wire[3:0] T6836;
  wire[3:0] T6837;
  wire[3:0] T6838;
  wire T6839;
  wire[3:0] T6840;
  wire T6841;
  wire T6842;
  wire[3:0] T6843;
  wire[3:0] T6844;
  wire T6845;
  wire[3:0] T6846;
  wire T6847;
  wire T6848;
  wire T6849;
  wire[3:0] T6850;
  wire[3:0] T6851;
  wire[3:0] T6852;
  wire T6853;
  wire[3:0] T6854;
  wire T6855;
  wire T6856;
  wire[3:0] T6857;
  wire[3:0] T6858;
  wire T6859;
  wire[3:0] T6860;
  wire T6861;
  wire T6862;
  wire T6863;
  wire T6864;
  wire[3:0] T6865;
  wire[3:0] T6866;
  wire[3:0] T6867;
  wire[3:0] T6868;
  wire T6869;
  wire[3:0] T6870;
  wire T6871;
  wire T6872;
  wire[3:0] T6873;
  wire[3:0] T6874;
  wire T6875;
  wire[3:0] T6876;
  wire T6877;
  wire T6878;
  wire T6879;
  wire[3:0] T6880;
  wire[3:0] T6881;
  wire[3:0] T6882;
  wire T6883;
  wire[3:0] T6884;
  wire T6885;
  wire T6886;
  wire[3:0] T6887;
  wire[3:0] T6888;
  wire T6889;
  wire[3:0] T6890;
  wire T6891;
  wire T6892;
  wire T6893;
  wire T6894;
  wire T6895;
  wire[3:0] T6896;
  wire[3:0] T6897;
  wire[3:0] T6898;
  wire[3:0] T6899;
  wire[3:0] T6900;
  wire T6901;
  wire[3:0] T6902;
  wire T6903;
  wire T6904;
  wire[3:0] T6905;
  wire[3:0] T6906;
  wire T6907;
  wire[3:0] T6908;
  wire T6909;
  wire T6910;
  wire T6911;
  wire[3:0] T6912;
  wire[3:0] T6913;
  wire[3:0] T6914;
  wire T6915;
  wire[3:0] T6916;
  wire T6917;
  wire T6918;
  wire[3:0] T6919;
  wire[3:0] T6920;
  wire T6921;
  wire[3:0] T6922;
  wire T6923;
  wire T6924;
  wire T6925;
  wire T6926;
  wire[3:0] T6927;
  wire[3:0] T6928;
  wire[3:0] T6929;
  wire[3:0] T6930;
  wire T6931;
  wire[3:0] T6932;
  wire T6933;
  wire T6934;
  wire[3:0] T6935;
  wire[3:0] T6936;
  wire T6937;
  wire[3:0] T6938;
  wire T6939;
  wire T6940;
  wire T6941;
  wire[3:0] T6942;
  wire[3:0] T6943;
  wire[3:0] T6944;
  wire T6945;
  wire[3:0] T6946;
  wire T6947;
  wire T6948;
  wire[3:0] T6949;
  wire[3:0] T6950;
  wire T6951;
  wire[3:0] T6952;
  wire T6953;
  wire T6954;
  wire T6955;
  wire T6956;
  wire T6957;
  wire T6958;
  wire T6959;
  wire[3:0] T6960;
  wire[3:0] T6961;
  wire[3:0] T6962;
  wire[3:0] T6963;
  wire[3:0] T6964;
  wire[3:0] T6965;
  wire[3:0] T6966;
  wire T6967;
  wire[3:0] T6968;
  wire T6969;
  wire T6970;
  wire[3:0] T6971;
  wire[3:0] T6972;
  wire T6973;
  wire[3:0] T6974;
  wire T6975;
  wire T6976;
  wire T6977;
  wire[3:0] T6978;
  wire[3:0] T6979;
  wire[3:0] T6980;
  wire T6981;
  wire[3:0] T6982;
  wire T6983;
  wire T6984;
  wire[3:0] T6985;
  wire[3:0] T6986;
  wire T6987;
  wire[3:0] T6988;
  wire T6989;
  wire T6990;
  wire T6991;
  wire T6992;
  wire[3:0] T6993;
  wire[3:0] T6994;
  wire[3:0] T6995;
  wire[3:0] T6996;
  wire T6997;
  wire[3:0] T6998;
  wire T6999;
  wire T7000;
  wire[3:0] T7001;
  wire[3:0] T7002;
  wire T7003;
  wire[3:0] T7004;
  wire T7005;
  wire T7006;
  wire T7007;
  wire[3:0] T7008;
  wire[3:0] T7009;
  wire[3:0] T7010;
  wire T7011;
  wire[3:0] T7012;
  wire T7013;
  wire T7014;
  wire[3:0] T7015;
  wire[3:0] T7016;
  wire T7017;
  wire[3:0] T7018;
  wire T7019;
  wire T7020;
  wire T7021;
  wire T7022;
  wire T7023;
  wire[3:0] T7024;
  wire[3:0] T7025;
  wire[3:0] T7026;
  wire[3:0] T7027;
  wire[3:0] T7028;
  wire T7029;
  wire[3:0] T7030;
  wire T7031;
  wire T7032;
  wire[3:0] T7033;
  wire[3:0] T7034;
  wire T7035;
  wire[3:0] T7036;
  wire T7037;
  wire T7038;
  wire T7039;
  wire[3:0] T7040;
  wire[3:0] T7041;
  wire[3:0] T7042;
  wire T7043;
  wire[3:0] T7044;
  wire T7045;
  wire T7046;
  wire[3:0] T7047;
  wire[3:0] T7048;
  wire T7049;
  wire[3:0] T7050;
  wire T7051;
  wire T7052;
  wire T7053;
  wire T7054;
  wire[3:0] T7055;
  wire[3:0] T7056;
  wire[3:0] T7057;
  wire[3:0] T7058;
  wire T7059;
  wire[3:0] T7060;
  wire T7061;
  wire T7062;
  wire[3:0] T7063;
  wire[3:0] T7064;
  wire T7065;
  wire[3:0] T7066;
  wire T7067;
  wire T7068;
  wire T7069;
  wire[3:0] T7070;
  wire[3:0] T7071;
  wire[3:0] T7072;
  wire T7073;
  wire[3:0] T7074;
  wire T7075;
  wire T7076;
  wire[3:0] T7077;
  wire[3:0] T7078;
  wire T7079;
  wire[3:0] T7080;
  wire T7081;
  wire T7082;
  wire T7083;
  wire T7084;
  wire T7085;
  wire T7086;
  wire[3:0] T7087;
  wire[3:0] T7088;
  wire[3:0] T7089;
  wire[3:0] T7090;
  wire[3:0] T7091;
  wire[3:0] T7092;
  wire T7093;
  wire[3:0] T7094;
  wire T7095;
  wire T7096;
  wire[3:0] T7097;
  wire[3:0] T7098;
  wire T7099;
  wire[3:0] T7100;
  wire T7101;
  wire T7102;
  wire T7103;
  wire[3:0] T7104;
  wire[3:0] T7105;
  wire[3:0] T7106;
  wire T7107;
  wire[3:0] T7108;
  wire T7109;
  wire T7110;
  wire[3:0] T7111;
  wire[3:0] T7112;
  wire T7113;
  wire[3:0] T7114;
  wire T7115;
  wire T7116;
  wire T7117;
  wire T7118;
  wire[3:0] T7119;
  wire[3:0] T7120;
  wire[3:0] T7121;
  wire[3:0] T7122;
  wire T7123;
  wire[3:0] T7124;
  wire T7125;
  wire T7126;
  wire[3:0] T7127;
  wire[3:0] T7128;
  wire T7129;
  wire[3:0] T7130;
  wire T7131;
  wire T7132;
  wire T7133;
  wire[3:0] T7134;
  wire[3:0] T7135;
  wire[3:0] T7136;
  wire T7137;
  wire[3:0] T7138;
  wire T7139;
  wire T7140;
  wire[3:0] T7141;
  wire[3:0] T7142;
  wire T7143;
  wire[3:0] T7144;
  wire T7145;
  wire T7146;
  wire T7147;
  wire T7148;
  wire T7149;
  wire[3:0] T7150;
  wire[3:0] T7151;
  wire[3:0] T7152;
  wire[3:0] T7153;
  wire[3:0] T7154;
  wire T7155;
  wire[3:0] T7156;
  wire T7157;
  wire T7158;
  wire[3:0] T7159;
  wire[3:0] T7160;
  wire T7161;
  wire[3:0] T7162;
  wire T7163;
  wire T7164;
  wire T7165;
  wire[3:0] T7166;
  wire[3:0] T7167;
  wire[3:0] T7168;
  wire T7169;
  wire[3:0] T7170;
  wire T7171;
  wire T7172;
  wire[3:0] T7173;
  wire[3:0] T7174;
  wire T7175;
  wire[3:0] T7176;
  wire T7177;
  wire T7178;
  wire T7179;
  wire T7180;
  wire[3:0] T7181;
  wire[3:0] T7182;
  wire[3:0] T7183;
  wire[3:0] T7184;
  wire T7185;
  wire[3:0] T7186;
  wire T7187;
  wire T7188;
  wire[3:0] T7189;
  wire[3:0] T7190;
  wire T7191;
  wire[3:0] T7192;
  wire T7193;
  wire T7194;
  wire T7195;
  wire[3:0] T7196;
  wire[3:0] T7197;
  wire[3:0] T7198;
  wire T7199;
  wire[3:0] T7200;
  wire T7201;
  wire T7202;
  wire[3:0] T7203;
  wire[3:0] T7204;
  wire T7205;
  wire[3:0] T7206;
  wire T7207;
  wire T7208;
  wire T7209;
  wire T7210;
  wire T7211;
  wire T7212;
  wire T7213;
  wire T7214;
  wire T7215;
  wire[3:0] T7216;
  wire[3:0] T7217;
  wire[3:0] T7218;
  wire[3:0] T7219;
  wire[3:0] T7220;
  wire[3:0] T7221;
  wire[3:0] T7222;
  wire[3:0] T7223;
  wire[3:0] T7224;
  wire T7225;
  wire[3:0] T7226;
  wire T7227;
  wire T7228;
  wire[3:0] T7229;
  wire[3:0] T7230;
  wire T7231;
  wire[3:0] T7232;
  wire T7233;
  wire T7234;
  wire T7235;
  wire[3:0] T7236;
  wire[3:0] T7237;
  wire[3:0] T7238;
  wire T7239;
  wire[3:0] T7240;
  wire T7241;
  wire T7242;
  wire[3:0] T7243;
  wire[3:0] T7244;
  wire T7245;
  wire[3:0] T7246;
  wire T7247;
  wire T7248;
  wire T7249;
  wire T7250;
  wire[3:0] T7251;
  wire[3:0] T7252;
  wire[3:0] T7253;
  wire[3:0] T7254;
  wire T7255;
  wire[3:0] T7256;
  wire T7257;
  wire T7258;
  wire[3:0] T7259;
  wire[3:0] T7260;
  wire T7261;
  wire[3:0] T7262;
  wire T7263;
  wire T7264;
  wire T7265;
  wire[3:0] T7266;
  wire[3:0] T7267;
  wire[3:0] T7268;
  wire T7269;
  wire[3:0] T7270;
  wire T7271;
  wire T7272;
  wire[3:0] T7273;
  wire[3:0] T7274;
  wire T7275;
  wire[3:0] T7276;
  wire T7277;
  wire T7278;
  wire T7279;
  wire T7280;
  wire T7281;
  wire[3:0] T7282;
  wire[3:0] T7283;
  wire[3:0] T7284;
  wire[3:0] T7285;
  wire[3:0] T7286;
  wire T7287;
  wire[3:0] T7288;
  wire T7289;
  wire T7290;
  wire[3:0] T7291;
  wire[3:0] T7292;
  wire T7293;
  wire[3:0] T7294;
  wire T7295;
  wire T7296;
  wire T7297;
  wire[3:0] T7298;
  wire[3:0] T7299;
  wire[3:0] T7300;
  wire T7301;
  wire[3:0] T7302;
  wire T7303;
  wire T7304;
  wire[3:0] T7305;
  wire[3:0] T7306;
  wire T7307;
  wire[3:0] T7308;
  wire T7309;
  wire T7310;
  wire T7311;
  wire T7312;
  wire[3:0] T7313;
  wire[3:0] T7314;
  wire[3:0] T7315;
  wire[3:0] T7316;
  wire T7317;
  wire[3:0] T7318;
  wire T7319;
  wire T7320;
  wire[3:0] T7321;
  wire[3:0] T7322;
  wire T7323;
  wire[3:0] T7324;
  wire T7325;
  wire T7326;
  wire T7327;
  wire[3:0] T7328;
  wire[3:0] T7329;
  wire[3:0] T7330;
  wire T7331;
  wire[3:0] T7332;
  wire T7333;
  wire T7334;
  wire[3:0] T7335;
  wire[3:0] T7336;
  wire T7337;
  wire[3:0] T7338;
  wire T7339;
  wire T7340;
  wire T7341;
  wire T7342;
  wire T7343;
  wire T7344;
  wire[3:0] T7345;
  wire[3:0] T7346;
  wire[3:0] T7347;
  wire[3:0] T7348;
  wire[3:0] T7349;
  wire[3:0] T7350;
  wire T7351;
  wire[3:0] T7352;
  wire T7353;
  wire T7354;
  wire[3:0] T7355;
  wire[3:0] T7356;
  wire T7357;
  wire[3:0] T7358;
  wire T7359;
  wire T7360;
  wire T7361;
  wire[3:0] T7362;
  wire[3:0] T7363;
  wire[3:0] T7364;
  wire T7365;
  wire[3:0] T7366;
  wire T7367;
  wire T7368;
  wire[3:0] T7369;
  wire[3:0] T7370;
  wire T7371;
  wire[3:0] T7372;
  wire T7373;
  wire T7374;
  wire T7375;
  wire T7376;
  wire[3:0] T7377;
  wire[3:0] T7378;
  wire[3:0] T7379;
  wire[3:0] T7380;
  wire T7381;
  wire[3:0] T7382;
  wire T7383;
  wire T7384;
  wire[3:0] T7385;
  wire[3:0] T7386;
  wire T7387;
  wire[3:0] T7388;
  wire T7389;
  wire T7390;
  wire T7391;
  wire[3:0] T7392;
  wire[3:0] T7393;
  wire[3:0] T7394;
  wire T7395;
  wire[3:0] T7396;
  wire T7397;
  wire T7398;
  wire[3:0] T7399;
  wire[3:0] T7400;
  wire T7401;
  wire[3:0] T7402;
  wire T7403;
  wire T7404;
  wire T7405;
  wire T7406;
  wire T7407;
  wire[3:0] T7408;
  wire[3:0] T7409;
  wire[3:0] T7410;
  wire[3:0] T7411;
  wire[3:0] T7412;
  wire T7413;
  wire[3:0] T7414;
  wire T7415;
  wire T7416;
  wire[3:0] T7417;
  wire[3:0] T7418;
  wire T7419;
  wire[3:0] T7420;
  wire T7421;
  wire T7422;
  wire T7423;
  wire[3:0] T7424;
  wire[3:0] T7425;
  wire[3:0] T7426;
  wire T7427;
  wire[3:0] T7428;
  wire T7429;
  wire T7430;
  wire[3:0] T7431;
  wire[3:0] T7432;
  wire T7433;
  wire[3:0] T7434;
  wire T7435;
  wire T7436;
  wire T7437;
  wire T7438;
  wire[3:0] T7439;
  wire[3:0] T7440;
  wire[3:0] T7441;
  wire[3:0] T7442;
  wire T7443;
  wire[3:0] T7444;
  wire T7445;
  wire T7446;
  wire[3:0] T7447;
  wire[3:0] T7448;
  wire T7449;
  wire[3:0] T7450;
  wire T7451;
  wire T7452;
  wire T7453;
  wire[3:0] T7454;
  wire[3:0] T7455;
  wire[3:0] T7456;
  wire T7457;
  wire[3:0] T7458;
  wire T7459;
  wire T7460;
  wire[3:0] T7461;
  wire[3:0] T7462;
  wire T7463;
  wire[3:0] T7464;
  wire T7465;
  wire T7466;
  wire T7467;
  wire T7468;
  wire T7469;
  wire T7470;
  wire T7471;
  wire[3:0] T7472;
  wire[3:0] T7473;
  wire[3:0] T7474;
  wire[3:0] T7475;
  wire[3:0] T7476;
  wire[3:0] T7477;
  wire[3:0] T7478;
  wire T7479;
  wire[3:0] T7480;
  wire T7481;
  wire T7482;
  wire[3:0] T7483;
  wire[3:0] T7484;
  wire T7485;
  wire[3:0] T7486;
  wire T7487;
  wire T7488;
  wire T7489;
  wire[3:0] T7490;
  wire[3:0] T7491;
  wire[3:0] T7492;
  wire T7493;
  wire[3:0] T7494;
  wire T7495;
  wire T7496;
  wire[3:0] T7497;
  wire[3:0] T7498;
  wire T7499;
  wire[3:0] T7500;
  wire T7501;
  wire T7502;
  wire T7503;
  wire T7504;
  wire[3:0] T7505;
  wire[3:0] T7506;
  wire[3:0] T7507;
  wire[3:0] T7508;
  wire T7509;
  wire[3:0] T7510;
  wire T7511;
  wire T7512;
  wire[3:0] T7513;
  wire[3:0] T7514;
  wire T7515;
  wire[3:0] T7516;
  wire T7517;
  wire T7518;
  wire T7519;
  wire[3:0] T7520;
  wire[3:0] T7521;
  wire[3:0] T7522;
  wire T7523;
  wire[3:0] T7524;
  wire T7525;
  wire T7526;
  wire[3:0] T7527;
  wire[3:0] T7528;
  wire T7529;
  wire[3:0] T7530;
  wire T7531;
  wire T7532;
  wire T7533;
  wire T7534;
  wire T7535;
  wire[3:0] T7536;
  wire[3:0] T7537;
  wire[3:0] T7538;
  wire[3:0] T7539;
  wire[3:0] T7540;
  wire T7541;
  wire[3:0] T7542;
  wire T7543;
  wire T7544;
  wire[3:0] T7545;
  wire[3:0] T7546;
  wire T7547;
  wire[3:0] T7548;
  wire T7549;
  wire T7550;
  wire T7551;
  wire[3:0] T7552;
  wire[3:0] T7553;
  wire[3:0] T7554;
  wire T7555;
  wire[3:0] T7556;
  wire T7557;
  wire T7558;
  wire[3:0] T7559;
  wire[3:0] T7560;
  wire T7561;
  wire[3:0] T7562;
  wire T7563;
  wire T7564;
  wire T7565;
  wire T7566;
  wire[3:0] T7567;
  wire[3:0] T7568;
  wire[3:0] T7569;
  wire[3:0] T7570;
  wire T7571;
  wire[3:0] T7572;
  wire T7573;
  wire T7574;
  wire[3:0] T7575;
  wire[3:0] T7576;
  wire T7577;
  wire[3:0] T7578;
  wire T7579;
  wire T7580;
  wire T7581;
  wire[3:0] T7582;
  wire[3:0] T7583;
  wire[3:0] T7584;
  wire T7585;
  wire[3:0] T7586;
  wire T7587;
  wire T7588;
  wire[3:0] T7589;
  wire[3:0] T7590;
  wire T7591;
  wire[3:0] T7592;
  wire T7593;
  wire T7594;
  wire T7595;
  wire T7596;
  wire T7597;
  wire T7598;
  wire[3:0] T7599;
  wire[3:0] T7600;
  wire[3:0] T7601;
  wire[3:0] T7602;
  wire[3:0] T7603;
  wire[3:0] T7604;
  wire T7605;
  wire[3:0] T7606;
  wire T7607;
  wire T7608;
  wire[3:0] T7609;
  wire[3:0] T7610;
  wire T7611;
  wire[3:0] T7612;
  wire T7613;
  wire T7614;
  wire T7615;
  wire[3:0] T7616;
  wire[3:0] T7617;
  wire[3:0] T7618;
  wire T7619;
  wire[3:0] T7620;
  wire T7621;
  wire T7622;
  wire[3:0] T7623;
  wire[3:0] T7624;
  wire T7625;
  wire[3:0] T7626;
  wire T7627;
  wire T7628;
  wire T7629;
  wire T7630;
  wire[3:0] T7631;
  wire[3:0] T7632;
  wire[3:0] T7633;
  wire[3:0] T7634;
  wire T7635;
  wire[3:0] T7636;
  wire T7637;
  wire T7638;
  wire[3:0] T7639;
  wire[3:0] T7640;
  wire T7641;
  wire[3:0] T7642;
  wire T7643;
  wire T7644;
  wire T7645;
  wire[3:0] T7646;
  wire[3:0] T7647;
  wire[3:0] T7648;
  wire T7649;
  wire[3:0] T7650;
  wire T7651;
  wire T7652;
  wire[3:0] T7653;
  wire[3:0] T7654;
  wire T7655;
  wire[3:0] T7656;
  wire T7657;
  wire T7658;
  wire T7659;
  wire T7660;
  wire T7661;
  wire[3:0] T7662;
  wire[3:0] T7663;
  wire[3:0] T7664;
  wire[3:0] T7665;
  wire[3:0] T7666;
  wire T7667;
  wire[3:0] T7668;
  wire T7669;
  wire T7670;
  wire[3:0] T7671;
  wire[3:0] T7672;
  wire T7673;
  wire[3:0] T7674;
  wire T7675;
  wire T7676;
  wire T7677;
  wire[3:0] T7678;
  wire[3:0] T7679;
  wire[3:0] T7680;
  wire T7681;
  wire[3:0] T7682;
  wire T7683;
  wire T7684;
  wire[3:0] T7685;
  wire[3:0] T7686;
  wire T7687;
  wire[3:0] T7688;
  wire T7689;
  wire T7690;
  wire T7691;
  wire T7692;
  wire[3:0] T7693;
  wire[3:0] T7694;
  wire[3:0] T7695;
  wire[3:0] T7696;
  wire T7697;
  wire[3:0] T7698;
  wire T7699;
  wire T7700;
  wire[3:0] T7701;
  wire[3:0] T7702;
  wire T7703;
  wire[3:0] T7704;
  wire T7705;
  wire T7706;
  wire T7707;
  wire[3:0] T7708;
  wire[3:0] T7709;
  wire[3:0] T7710;
  wire T7711;
  wire[3:0] T7712;
  wire T7713;
  wire T7714;
  wire[3:0] T7715;
  wire[3:0] T7716;
  wire T7717;
  wire[3:0] T7718;
  wire T7719;
  wire T7720;
  wire T7721;
  wire T7722;
  wire T7723;
  wire T7724;
  wire T7725;
  wire T7726;
  wire[3:0] T7727;
  wire[3:0] T7728;
  wire[3:0] T7729;
  wire[3:0] T7730;
  wire[3:0] T7731;
  wire[3:0] T7732;
  wire[3:0] T7733;
  wire[3:0] T7734;
  wire T7735;
  wire[3:0] T7736;
  wire T7737;
  wire T7738;
  wire[3:0] T7739;
  wire[3:0] T7740;
  wire T7741;
  wire[3:0] T7742;
  wire T7743;
  wire T7744;
  wire T7745;
  wire[3:0] T7746;
  wire[3:0] T7747;
  wire[3:0] T7748;
  wire T7749;
  wire[3:0] T7750;
  wire T7751;
  wire T7752;
  wire[3:0] T7753;
  wire[3:0] T7754;
  wire T7755;
  wire[3:0] T7756;
  wire T7757;
  wire T7758;
  wire T7759;
  wire T7760;
  wire[3:0] T7761;
  wire[3:0] T7762;
  wire[3:0] T7763;
  wire[3:0] T7764;
  wire T7765;
  wire[3:0] T7766;
  wire T7767;
  wire T7768;
  wire[3:0] T7769;
  wire[3:0] T7770;
  wire T7771;
  wire[3:0] T7772;
  wire T7773;
  wire T7774;
  wire T7775;
  wire[3:0] T7776;
  wire[3:0] T7777;
  wire[3:0] T7778;
  wire T7779;
  wire[3:0] T7780;
  wire T7781;
  wire T7782;
  wire[3:0] T7783;
  wire[3:0] T7784;
  wire T7785;
  wire[3:0] T7786;
  wire T7787;
  wire T7788;
  wire T7789;
  wire T7790;
  wire T7791;
  wire[3:0] T7792;
  wire[3:0] T7793;
  wire[3:0] T7794;
  wire[3:0] T7795;
  wire[3:0] T7796;
  wire T7797;
  wire[3:0] T7798;
  wire T7799;
  wire T7800;
  wire[3:0] T7801;
  wire[3:0] T7802;
  wire T7803;
  wire[3:0] T7804;
  wire T7805;
  wire T7806;
  wire T7807;
  wire[3:0] T7808;
  wire[3:0] T7809;
  wire[3:0] T7810;
  wire T7811;
  wire[3:0] T7812;
  wire T7813;
  wire T7814;
  wire[3:0] T7815;
  wire[3:0] T7816;
  wire T7817;
  wire[3:0] T7818;
  wire T7819;
  wire T7820;
  wire T7821;
  wire T7822;
  wire[3:0] T7823;
  wire[3:0] T7824;
  wire[3:0] T7825;
  wire[3:0] T7826;
  wire T7827;
  wire[3:0] T7828;
  wire T7829;
  wire T7830;
  wire[3:0] T7831;
  wire[3:0] T7832;
  wire T7833;
  wire[3:0] T7834;
  wire T7835;
  wire T7836;
  wire T7837;
  wire[3:0] T7838;
  wire[3:0] T7839;
  wire[3:0] T7840;
  wire T7841;
  wire[3:0] T7842;
  wire T7843;
  wire T7844;
  wire[3:0] T7845;
  wire[3:0] T7846;
  wire T7847;
  wire[3:0] T7848;
  wire T7849;
  wire T7850;
  wire T7851;
  wire T7852;
  wire T7853;
  wire T7854;
  wire[3:0] T7855;
  wire[3:0] T7856;
  wire[3:0] T7857;
  wire[3:0] T7858;
  wire[3:0] T7859;
  wire[3:0] T7860;
  wire T7861;
  wire[3:0] T7862;
  wire T7863;
  wire T7864;
  wire[3:0] T7865;
  wire[3:0] T7866;
  wire T7867;
  wire[3:0] T7868;
  wire T7869;
  wire T7870;
  wire T7871;
  wire[3:0] T7872;
  wire[3:0] T7873;
  wire[3:0] T7874;
  wire T7875;
  wire[3:0] T7876;
  wire T7877;
  wire T7878;
  wire[3:0] T7879;
  wire[3:0] T7880;
  wire T7881;
  wire[3:0] T7882;
  wire T7883;
  wire T7884;
  wire T7885;
  wire T7886;
  wire[3:0] T7887;
  wire[3:0] T7888;
  wire[3:0] T7889;
  wire[3:0] T7890;
  wire T7891;
  wire[3:0] T7892;
  wire T7893;
  wire T7894;
  wire[3:0] T7895;
  wire[3:0] T7896;
  wire T7897;
  wire[3:0] T7898;
  wire T7899;
  wire T7900;
  wire T7901;
  wire[3:0] T7902;
  wire[3:0] T7903;
  wire[3:0] T7904;
  wire T7905;
  wire[3:0] T7906;
  wire T7907;
  wire T7908;
  wire[3:0] T7909;
  wire[3:0] T7910;
  wire T7911;
  wire[3:0] T7912;
  wire T7913;
  wire T7914;
  wire T7915;
  wire T7916;
  wire T7917;
  wire[3:0] T7918;
  wire[3:0] T7919;
  wire[3:0] T7920;
  wire[3:0] T7921;
  wire[3:0] T7922;
  wire T7923;
  wire[3:0] T7924;
  wire T7925;
  wire T7926;
  wire[3:0] T7927;
  wire[3:0] T7928;
  wire T7929;
  wire[3:0] T7930;
  wire T7931;
  wire T7932;
  wire T7933;
  wire[3:0] T7934;
  wire[3:0] T7935;
  wire[3:0] T7936;
  wire T7937;
  wire[3:0] T7938;
  wire T7939;
  wire T7940;
  wire[3:0] T7941;
  wire[3:0] T7942;
  wire T7943;
  wire[3:0] T7944;
  wire T7945;
  wire T7946;
  wire T7947;
  wire T7948;
  wire[3:0] T7949;
  wire[3:0] T7950;
  wire[3:0] T7951;
  wire[3:0] T7952;
  wire T7953;
  wire[3:0] T7954;
  wire T7955;
  wire T7956;
  wire[3:0] T7957;
  wire[3:0] T7958;
  wire T7959;
  wire[3:0] T7960;
  wire T7961;
  wire T7962;
  wire T7963;
  wire[3:0] T7964;
  wire[3:0] T7965;
  wire[3:0] T7966;
  wire T7967;
  wire[3:0] T7968;
  wire T7969;
  wire T7970;
  wire[3:0] T7971;
  wire[3:0] T7972;
  wire T7973;
  wire[3:0] T7974;
  wire T7975;
  wire T7976;
  wire T7977;
  wire T7978;
  wire T7979;
  wire T7980;
  wire T7981;
  wire[3:0] T7982;
  wire[3:0] T7983;
  wire[3:0] T7984;
  wire[3:0] T7985;
  wire[3:0] T7986;
  wire[3:0] T7987;
  wire[3:0] T7988;
  wire T7989;
  wire[3:0] T7990;
  wire T7991;
  wire T7992;
  wire[3:0] T7993;
  wire[3:0] T7994;
  wire T7995;
  wire[3:0] T7996;
  wire T7997;
  wire T7998;
  wire T7999;
  wire[3:0] T8000;
  wire[3:0] T8001;
  wire[3:0] T8002;
  wire T8003;
  wire[3:0] T8004;
  wire T8005;
  wire T8006;
  wire[3:0] T8007;
  wire[3:0] T8008;
  wire T8009;
  wire[3:0] T8010;
  wire T8011;
  wire T8012;
  wire T8013;
  wire T8014;
  wire[3:0] T8015;
  wire[3:0] T8016;
  wire[3:0] T8017;
  wire[3:0] T8018;
  wire T8019;
  wire[3:0] T8020;
  wire T8021;
  wire T8022;
  wire[3:0] T8023;
  wire[3:0] T8024;
  wire T8025;
  wire[3:0] T8026;
  wire T8027;
  wire T8028;
  wire T8029;
  wire[3:0] T8030;
  wire[3:0] T8031;
  wire[3:0] T8032;
  wire T8033;
  wire[3:0] T8034;
  wire T8035;
  wire T8036;
  wire[3:0] T8037;
  wire[3:0] T8038;
  wire T8039;
  wire[3:0] T8040;
  wire T8041;
  wire T8042;
  wire T8043;
  wire T8044;
  wire T8045;
  wire[3:0] T8046;
  wire[3:0] T8047;
  wire[3:0] T8048;
  wire[3:0] T8049;
  wire[3:0] T8050;
  wire T8051;
  wire[3:0] T8052;
  wire T8053;
  wire T8054;
  wire[3:0] T8055;
  wire[3:0] T8056;
  wire T8057;
  wire[3:0] T8058;
  wire T8059;
  wire T8060;
  wire T8061;
  wire[3:0] T8062;
  wire[3:0] T8063;
  wire[3:0] T8064;
  wire T8065;
  wire[3:0] T8066;
  wire T8067;
  wire T8068;
  wire[3:0] T8069;
  wire[3:0] T8070;
  wire T8071;
  wire[3:0] T8072;
  wire T8073;
  wire T8074;
  wire T8075;
  wire T8076;
  wire[3:0] T8077;
  wire[3:0] T8078;
  wire[3:0] T8079;
  wire[3:0] T8080;
  wire T8081;
  wire[3:0] T8082;
  wire T8083;
  wire T8084;
  wire[3:0] T8085;
  wire[3:0] T8086;
  wire T8087;
  wire[3:0] T8088;
  wire T8089;
  wire T8090;
  wire T8091;
  wire[3:0] T8092;
  wire[3:0] T8093;
  wire[3:0] T8094;
  wire T8095;
  wire[3:0] T8096;
  wire T8097;
  wire T8098;
  wire[3:0] T8099;
  wire[3:0] T8100;
  wire T8101;
  wire[3:0] T8102;
  wire T8103;
  wire T8104;
  wire T8105;
  wire T8106;
  wire T8107;
  wire T8108;
  wire[3:0] T8109;
  wire[3:0] T8110;
  wire[3:0] T8111;
  wire[3:0] T8112;
  wire[3:0] T8113;
  wire[3:0] T8114;
  wire T8115;
  wire[3:0] T8116;
  wire T8117;
  wire T8118;
  wire[3:0] T8119;
  wire[3:0] T8120;
  wire T8121;
  wire[3:0] T8122;
  wire T8123;
  wire T8124;
  wire T8125;
  wire[3:0] T8126;
  wire[3:0] T8127;
  wire[3:0] T8128;
  wire T8129;
  wire[3:0] T8130;
  wire T8131;
  wire T8132;
  wire[3:0] T8133;
  wire[3:0] T8134;
  wire T8135;
  wire[3:0] T8136;
  wire T8137;
  wire T8138;
  wire T8139;
  wire T8140;
  wire[3:0] T8141;
  wire[3:0] T8142;
  wire[3:0] T8143;
  wire[3:0] T8144;
  wire T8145;
  wire[3:0] T8146;
  wire T8147;
  wire T8148;
  wire[3:0] T8149;
  wire[3:0] T8150;
  wire T8151;
  wire[3:0] T8152;
  wire T8153;
  wire T8154;
  wire T8155;
  wire[3:0] T8156;
  wire[3:0] T8157;
  wire[3:0] T8158;
  wire T8159;
  wire[3:0] T8160;
  wire T8161;
  wire T8162;
  wire[3:0] T8163;
  wire[3:0] T8164;
  wire T8165;
  wire[3:0] T8166;
  wire T8167;
  wire T8168;
  wire T8169;
  wire T8170;
  wire T8171;
  wire[3:0] T8172;
  wire[3:0] T8173;
  wire[3:0] T8174;
  wire[3:0] T8175;
  wire[3:0] T8176;
  wire T8177;
  wire[3:0] T8178;
  wire T8179;
  wire T8180;
  wire[3:0] T8181;
  wire[3:0] T8182;
  wire T8183;
  wire[3:0] T8184;
  wire T8185;
  wire T8186;
  wire T8187;
  wire[3:0] T8188;
  wire[3:0] T8189;
  wire[3:0] T8190;
  wire T8191;
  wire[3:0] T8192;
  wire T8193;
  wire T8194;
  wire[3:0] T8195;
  wire[3:0] T8196;
  wire T8197;
  wire[3:0] T8198;
  wire T8199;
  wire T8200;
  wire T8201;
  wire T8202;
  wire[3:0] T8203;
  wire[3:0] T8204;
  wire[3:0] T8205;
  wire[3:0] T8206;
  wire T8207;
  wire[3:0] T8208;
  wire T8209;
  wire T8210;
  wire[3:0] T8211;
  wire[3:0] T8212;
  wire T8213;
  wire[3:0] T8214;
  wire T8215;
  wire T8216;
  wire T8217;
  wire[3:0] T8218;
  wire[3:0] T8219;
  wire[3:0] T8220;
  wire T8221;
  wire[3:0] T8222;
  wire T8223;
  wire T8224;
  wire[3:0] T8225;
  wire[3:0] T8226;
  wire T8227;
  wire[3:0] T8228;
  wire T8229;
  wire T8230;
  wire T8231;
  wire T8232;
  wire T8233;
  wire T8234;
  wire T8235;
  wire T8236;
  wire T8237;
  wire T8238;
  reg [3:0] hashCount1;
  wire[3:0] T11370;
  wire[3:0] T8239;
  wire[3:0] T8240;
  wire[3:0] T8241;
  wire[3:0] T8242;
  wire[3:0] T8243;
  wire[3:0] T8244;
  wire[3:0] T8245;
  wire[3:0] T8246;
  wire[3:0] T8247;
  wire[3:0] T8248;
  wire[3:0] T8249;
  wire T8250;
  wire[9:0] T8251;
  wire[3:0] T8252;
  wire T8253;
  wire T8254;
  wire[3:0] T8255;
  wire[3:0] T8256;
  wire T8257;
  wire[3:0] T8258;
  wire T8259;
  wire T8260;
  wire T8261;
  wire[3:0] T8262;
  wire[3:0] T8263;
  wire[3:0] T8264;
  wire T8265;
  wire[3:0] T8266;
  wire T8267;
  wire T8268;
  wire[3:0] T8269;
  wire[3:0] T8270;
  wire T8271;
  wire[3:0] T8272;
  wire T8273;
  wire T8274;
  wire T8275;
  wire T8276;
  wire[3:0] T8277;
  wire[3:0] T8278;
  wire[3:0] T8279;
  wire[3:0] T8280;
  wire T8281;
  wire[3:0] T8282;
  wire T8283;
  wire T8284;
  wire[3:0] T8285;
  wire[3:0] T8286;
  wire T8287;
  wire[3:0] T8288;
  wire T8289;
  wire T8290;
  wire T8291;
  wire[3:0] T8292;
  wire[3:0] T8293;
  wire[3:0] T8294;
  wire T8295;
  wire[3:0] T8296;
  wire T8297;
  wire T8298;
  wire[3:0] T8299;
  wire[3:0] T8300;
  wire T8301;
  wire[3:0] T8302;
  wire T8303;
  wire T8304;
  wire T8305;
  wire T8306;
  wire T8307;
  wire[3:0] T8308;
  wire[3:0] T8309;
  wire[3:0] T8310;
  wire[3:0] T8311;
  wire[3:0] T8312;
  wire T8313;
  wire[3:0] T8314;
  wire T8315;
  wire T8316;
  wire[3:0] T8317;
  wire[3:0] T8318;
  wire T8319;
  wire[3:0] T8320;
  wire T8321;
  wire T8322;
  wire T8323;
  wire[3:0] T8324;
  wire[3:0] T8325;
  wire[3:0] T8326;
  wire T8327;
  wire[3:0] T8328;
  wire T8329;
  wire T8330;
  wire[3:0] T8331;
  wire[3:0] T8332;
  wire T8333;
  wire[3:0] T8334;
  wire T8335;
  wire T8336;
  wire T8337;
  wire T8338;
  wire[3:0] T8339;
  wire[3:0] T8340;
  wire[3:0] T8341;
  wire[3:0] T8342;
  wire T8343;
  wire[3:0] T8344;
  wire T8345;
  wire T8346;
  wire[3:0] T8347;
  wire[3:0] T8348;
  wire T8349;
  wire[3:0] T8350;
  wire T8351;
  wire T8352;
  wire T8353;
  wire[3:0] T8354;
  wire[3:0] T8355;
  wire[3:0] T8356;
  wire T8357;
  wire[3:0] T8358;
  wire T8359;
  wire T8360;
  wire[3:0] T8361;
  wire[3:0] T8362;
  wire T8363;
  wire[3:0] T8364;
  wire T8365;
  wire T8366;
  wire T8367;
  wire T8368;
  wire T8369;
  wire T8370;
  wire[3:0] T8371;
  wire[3:0] T8372;
  wire[3:0] T8373;
  wire[3:0] T8374;
  wire[3:0] T8375;
  wire[3:0] T8376;
  wire T8377;
  wire[3:0] T8378;
  wire T8379;
  wire T8380;
  wire[3:0] T8381;
  wire[3:0] T8382;
  wire T8383;
  wire[3:0] T8384;
  wire T8385;
  wire T8386;
  wire T8387;
  wire[3:0] T8388;
  wire[3:0] T8389;
  wire[3:0] T8390;
  wire T8391;
  wire[3:0] T8392;
  wire T8393;
  wire T8394;
  wire[3:0] T8395;
  wire[3:0] T8396;
  wire T8397;
  wire[3:0] T8398;
  wire T8399;
  wire T8400;
  wire T8401;
  wire T8402;
  wire[3:0] T8403;
  wire[3:0] T8404;
  wire[3:0] T8405;
  wire[3:0] T8406;
  wire T8407;
  wire[3:0] T8408;
  wire T8409;
  wire T8410;
  wire[3:0] T8411;
  wire[3:0] T8412;
  wire T8413;
  wire[3:0] T8414;
  wire T8415;
  wire T8416;
  wire T8417;
  wire[3:0] T8418;
  wire[3:0] T8419;
  wire[3:0] T8420;
  wire T8421;
  wire[3:0] T8422;
  wire T8423;
  wire T8424;
  wire[3:0] T8425;
  wire[3:0] T8426;
  wire T8427;
  wire[3:0] T8428;
  wire T8429;
  wire T8430;
  wire T8431;
  wire T8432;
  wire T8433;
  wire[3:0] T8434;
  wire[3:0] T8435;
  wire[3:0] T8436;
  wire[3:0] T8437;
  wire[3:0] T8438;
  wire T8439;
  wire[3:0] T8440;
  wire T8441;
  wire T8442;
  wire[3:0] T8443;
  wire[3:0] T8444;
  wire T8445;
  wire[3:0] T8446;
  wire T8447;
  wire T8448;
  wire T8449;
  wire[3:0] T8450;
  wire[3:0] T8451;
  wire[3:0] T8452;
  wire T8453;
  wire[3:0] T8454;
  wire T8455;
  wire T8456;
  wire[3:0] T8457;
  wire[3:0] T8458;
  wire T8459;
  wire[3:0] T8460;
  wire T8461;
  wire T8462;
  wire T8463;
  wire T8464;
  wire[3:0] T8465;
  wire[3:0] T8466;
  wire[3:0] T8467;
  wire[3:0] T8468;
  wire T8469;
  wire[3:0] T8470;
  wire T8471;
  wire T8472;
  wire[3:0] T8473;
  wire[3:0] T8474;
  wire T8475;
  wire[3:0] T8476;
  wire T8477;
  wire T8478;
  wire T8479;
  wire[3:0] T8480;
  wire[3:0] T8481;
  wire[3:0] T8482;
  wire T8483;
  wire[3:0] T8484;
  wire T8485;
  wire T8486;
  wire[3:0] T8487;
  wire[3:0] T8488;
  wire T8489;
  wire[3:0] T8490;
  wire T8491;
  wire T8492;
  wire T8493;
  wire T8494;
  wire T8495;
  wire T8496;
  wire T8497;
  wire[3:0] T8498;
  wire[3:0] T8499;
  wire[3:0] T8500;
  wire[3:0] T8501;
  wire[3:0] T8502;
  wire[3:0] T8503;
  wire[3:0] T8504;
  wire T8505;
  wire[3:0] T8506;
  wire T8507;
  wire T8508;
  wire[3:0] T8509;
  wire[3:0] T8510;
  wire T8511;
  wire[3:0] T8512;
  wire T8513;
  wire T8514;
  wire T8515;
  wire[3:0] T8516;
  wire[3:0] T8517;
  wire[3:0] T8518;
  wire T8519;
  wire[3:0] T8520;
  wire T8521;
  wire T8522;
  wire[3:0] T8523;
  wire[3:0] T8524;
  wire T8525;
  wire[3:0] T8526;
  wire T8527;
  wire T8528;
  wire T8529;
  wire T8530;
  wire[3:0] T8531;
  wire[3:0] T8532;
  wire[3:0] T8533;
  wire[3:0] T8534;
  wire T8535;
  wire[3:0] T8536;
  wire T8537;
  wire T8538;
  wire[3:0] T8539;
  wire[3:0] T8540;
  wire T8541;
  wire[3:0] T8542;
  wire T8543;
  wire T8544;
  wire T8545;
  wire[3:0] T8546;
  wire[3:0] T8547;
  wire[3:0] T8548;
  wire T8549;
  wire[3:0] T8550;
  wire T8551;
  wire T8552;
  wire[3:0] T8553;
  wire[3:0] T8554;
  wire T8555;
  wire[3:0] T8556;
  wire T8557;
  wire T8558;
  wire T8559;
  wire T8560;
  wire T8561;
  wire[3:0] T8562;
  wire[3:0] T8563;
  wire[3:0] T8564;
  wire[3:0] T8565;
  wire[3:0] T8566;
  wire T8567;
  wire[3:0] T8568;
  wire T8569;
  wire T8570;
  wire[3:0] T8571;
  wire[3:0] T8572;
  wire T8573;
  wire[3:0] T8574;
  wire T8575;
  wire T8576;
  wire T8577;
  wire[3:0] T8578;
  wire[3:0] T8579;
  wire[3:0] T8580;
  wire T8581;
  wire[3:0] T8582;
  wire T8583;
  wire T8584;
  wire[3:0] T8585;
  wire[3:0] T8586;
  wire T8587;
  wire[3:0] T8588;
  wire T8589;
  wire T8590;
  wire T8591;
  wire T8592;
  wire[3:0] T8593;
  wire[3:0] T8594;
  wire[3:0] T8595;
  wire[3:0] T8596;
  wire T8597;
  wire[3:0] T8598;
  wire T8599;
  wire T8600;
  wire[3:0] T8601;
  wire[3:0] T8602;
  wire T8603;
  wire[3:0] T8604;
  wire T8605;
  wire T8606;
  wire T8607;
  wire[3:0] T8608;
  wire[3:0] T8609;
  wire[3:0] T8610;
  wire T8611;
  wire[3:0] T8612;
  wire T8613;
  wire T8614;
  wire[3:0] T8615;
  wire[3:0] T8616;
  wire T8617;
  wire[3:0] T8618;
  wire T8619;
  wire T8620;
  wire T8621;
  wire T8622;
  wire T8623;
  wire T8624;
  wire[3:0] T8625;
  wire[3:0] T8626;
  wire[3:0] T8627;
  wire[3:0] T8628;
  wire[3:0] T8629;
  wire[3:0] T8630;
  wire T8631;
  wire[3:0] T8632;
  wire T8633;
  wire T8634;
  wire[3:0] T8635;
  wire[3:0] T8636;
  wire T8637;
  wire[3:0] T8638;
  wire T8639;
  wire T8640;
  wire T8641;
  wire[3:0] T8642;
  wire[3:0] T8643;
  wire[3:0] T8644;
  wire T8645;
  wire[3:0] T8646;
  wire T8647;
  wire T8648;
  wire[3:0] T8649;
  wire[3:0] T8650;
  wire T8651;
  wire[3:0] T8652;
  wire T8653;
  wire T8654;
  wire T8655;
  wire T8656;
  wire[3:0] T8657;
  wire[3:0] T8658;
  wire[3:0] T8659;
  wire[3:0] T8660;
  wire T8661;
  wire[3:0] T8662;
  wire T8663;
  wire T8664;
  wire[3:0] T8665;
  wire[3:0] T8666;
  wire T8667;
  wire[3:0] T8668;
  wire T8669;
  wire T8670;
  wire T8671;
  wire[3:0] T8672;
  wire[3:0] T8673;
  wire[3:0] T8674;
  wire T8675;
  wire[3:0] T8676;
  wire T8677;
  wire T8678;
  wire[3:0] T8679;
  wire[3:0] T8680;
  wire T8681;
  wire[3:0] T8682;
  wire T8683;
  wire T8684;
  wire T8685;
  wire T8686;
  wire T8687;
  wire[3:0] T8688;
  wire[3:0] T8689;
  wire[3:0] T8690;
  wire[3:0] T8691;
  wire[3:0] T8692;
  wire T8693;
  wire[3:0] T8694;
  wire T8695;
  wire T8696;
  wire[3:0] T8697;
  wire[3:0] T8698;
  wire T8699;
  wire[3:0] T8700;
  wire T8701;
  wire T8702;
  wire T8703;
  wire[3:0] T8704;
  wire[3:0] T8705;
  wire[3:0] T8706;
  wire T8707;
  wire[3:0] T8708;
  wire T8709;
  wire T8710;
  wire[3:0] T8711;
  wire[3:0] T8712;
  wire T8713;
  wire[3:0] T8714;
  wire T8715;
  wire T8716;
  wire T8717;
  wire T8718;
  wire[3:0] T8719;
  wire[3:0] T8720;
  wire[3:0] T8721;
  wire[3:0] T8722;
  wire T8723;
  wire[3:0] T8724;
  wire T8725;
  wire T8726;
  wire[3:0] T8727;
  wire[3:0] T8728;
  wire T8729;
  wire[3:0] T8730;
  wire T8731;
  wire T8732;
  wire T8733;
  wire[3:0] T8734;
  wire[3:0] T8735;
  wire[3:0] T8736;
  wire T8737;
  wire[3:0] T8738;
  wire T8739;
  wire T8740;
  wire[3:0] T8741;
  wire[3:0] T8742;
  wire T8743;
  wire[3:0] T8744;
  wire T8745;
  wire T8746;
  wire T8747;
  wire T8748;
  wire T8749;
  wire T8750;
  wire T8751;
  wire T8752;
  wire[3:0] T8753;
  wire[3:0] T8754;
  wire[3:0] T8755;
  wire[3:0] T8756;
  wire[3:0] T8757;
  wire[3:0] T8758;
  wire[3:0] T8759;
  wire[3:0] T8760;
  wire T8761;
  wire[3:0] T8762;
  wire T8763;
  wire T8764;
  wire[3:0] T8765;
  wire[3:0] T8766;
  wire T8767;
  wire[3:0] T8768;
  wire T8769;
  wire T8770;
  wire T8771;
  wire[3:0] T8772;
  wire[3:0] T8773;
  wire[3:0] T8774;
  wire T8775;
  wire[3:0] T8776;
  wire T8777;
  wire T8778;
  wire[3:0] T8779;
  wire[3:0] T8780;
  wire T8781;
  wire[3:0] T8782;
  wire T8783;
  wire T8784;
  wire T8785;
  wire T8786;
  wire[3:0] T8787;
  wire[3:0] T8788;
  wire[3:0] T8789;
  wire[3:0] T8790;
  wire T8791;
  wire[3:0] T8792;
  wire T8793;
  wire T8794;
  wire[3:0] T8795;
  wire[3:0] T8796;
  wire T8797;
  wire[3:0] T8798;
  wire T8799;
  wire T8800;
  wire T8801;
  wire[3:0] T8802;
  wire[3:0] T8803;
  wire[3:0] T8804;
  wire T8805;
  wire[3:0] T8806;
  wire T8807;
  wire T8808;
  wire[3:0] T8809;
  wire[3:0] T8810;
  wire T8811;
  wire[3:0] T8812;
  wire T8813;
  wire T8814;
  wire T8815;
  wire T8816;
  wire T8817;
  wire[3:0] T8818;
  wire[3:0] T8819;
  wire[3:0] T8820;
  wire[3:0] T8821;
  wire[3:0] T8822;
  wire T8823;
  wire[3:0] T8824;
  wire T8825;
  wire T8826;
  wire[3:0] T8827;
  wire[3:0] T8828;
  wire T8829;
  wire[3:0] T8830;
  wire T8831;
  wire T8832;
  wire T8833;
  wire[3:0] T8834;
  wire[3:0] T8835;
  wire[3:0] T8836;
  wire T8837;
  wire[3:0] T8838;
  wire T8839;
  wire T8840;
  wire[3:0] T8841;
  wire[3:0] T8842;
  wire T8843;
  wire[3:0] T8844;
  wire T8845;
  wire T8846;
  wire T8847;
  wire T8848;
  wire[3:0] T8849;
  wire[3:0] T8850;
  wire[3:0] T8851;
  wire[3:0] T8852;
  wire T8853;
  wire[3:0] T8854;
  wire T8855;
  wire T8856;
  wire[3:0] T8857;
  wire[3:0] T8858;
  wire T8859;
  wire[3:0] T8860;
  wire T8861;
  wire T8862;
  wire T8863;
  wire[3:0] T8864;
  wire[3:0] T8865;
  wire[3:0] T8866;
  wire T8867;
  wire[3:0] T8868;
  wire T8869;
  wire T8870;
  wire[3:0] T8871;
  wire[3:0] T8872;
  wire T8873;
  wire[3:0] T8874;
  wire T8875;
  wire T8876;
  wire T8877;
  wire T8878;
  wire T8879;
  wire T8880;
  wire[3:0] T8881;
  wire[3:0] T8882;
  wire[3:0] T8883;
  wire[3:0] T8884;
  wire[3:0] T8885;
  wire[3:0] T8886;
  wire T8887;
  wire[3:0] T8888;
  wire T8889;
  wire T8890;
  wire[3:0] T8891;
  wire[3:0] T8892;
  wire T8893;
  wire[3:0] T8894;
  wire T8895;
  wire T8896;
  wire T8897;
  wire[3:0] T8898;
  wire[3:0] T8899;
  wire[3:0] T8900;
  wire T8901;
  wire[3:0] T8902;
  wire T8903;
  wire T8904;
  wire[3:0] T8905;
  wire[3:0] T8906;
  wire T8907;
  wire[3:0] T8908;
  wire T8909;
  wire T8910;
  wire T8911;
  wire T8912;
  wire[3:0] T8913;
  wire[3:0] T8914;
  wire[3:0] T8915;
  wire[3:0] T8916;
  wire T8917;
  wire[3:0] T8918;
  wire T8919;
  wire T8920;
  wire[3:0] T8921;
  wire[3:0] T8922;
  wire T8923;
  wire[3:0] T8924;
  wire T8925;
  wire T8926;
  wire T8927;
  wire[3:0] T8928;
  wire[3:0] T8929;
  wire[3:0] T8930;
  wire T8931;
  wire[3:0] T8932;
  wire T8933;
  wire T8934;
  wire[3:0] T8935;
  wire[3:0] T8936;
  wire T8937;
  wire[3:0] T8938;
  wire T8939;
  wire T8940;
  wire T8941;
  wire T8942;
  wire T8943;
  wire[3:0] T8944;
  wire[3:0] T8945;
  wire[3:0] T8946;
  wire[3:0] T8947;
  wire[3:0] T8948;
  wire T8949;
  wire[3:0] T8950;
  wire T8951;
  wire T8952;
  wire[3:0] T8953;
  wire[3:0] T8954;
  wire T8955;
  wire[3:0] T8956;
  wire T8957;
  wire T8958;
  wire T8959;
  wire[3:0] T8960;
  wire[3:0] T8961;
  wire[3:0] T8962;
  wire T8963;
  wire[3:0] T8964;
  wire T8965;
  wire T8966;
  wire[3:0] T8967;
  wire[3:0] T8968;
  wire T8969;
  wire[3:0] T8970;
  wire T8971;
  wire T8972;
  wire T8973;
  wire T8974;
  wire[3:0] T8975;
  wire[3:0] T8976;
  wire[3:0] T8977;
  wire[3:0] T8978;
  wire T8979;
  wire[3:0] T8980;
  wire T8981;
  wire T8982;
  wire[3:0] T8983;
  wire[3:0] T8984;
  wire T8985;
  wire[3:0] T8986;
  wire T8987;
  wire T8988;
  wire T8989;
  wire[3:0] T8990;
  wire[3:0] T8991;
  wire[3:0] T8992;
  wire T8993;
  wire[3:0] T8994;
  wire T8995;
  wire T8996;
  wire[3:0] T8997;
  wire[3:0] T8998;
  wire T8999;
  wire[3:0] T9000;
  wire T9001;
  wire T9002;
  wire T9003;
  wire T9004;
  wire T9005;
  wire T9006;
  wire T9007;
  wire[3:0] T9008;
  wire[3:0] T9009;
  wire[3:0] T9010;
  wire[3:0] T9011;
  wire[3:0] T9012;
  wire[3:0] T9013;
  wire[3:0] T9014;
  wire T9015;
  wire[3:0] T9016;
  wire T9017;
  wire T9018;
  wire[3:0] T9019;
  wire[3:0] T9020;
  wire T9021;
  wire[3:0] T9022;
  wire T9023;
  wire T9024;
  wire T9025;
  wire[3:0] T9026;
  wire[3:0] T9027;
  wire[3:0] T9028;
  wire T9029;
  wire[3:0] T9030;
  wire T9031;
  wire T9032;
  wire[3:0] T9033;
  wire[3:0] T9034;
  wire T9035;
  wire[3:0] T9036;
  wire T9037;
  wire T9038;
  wire T9039;
  wire T9040;
  wire[3:0] T9041;
  wire[3:0] T9042;
  wire[3:0] T9043;
  wire[3:0] T9044;
  wire T9045;
  wire[3:0] T9046;
  wire T9047;
  wire T9048;
  wire[3:0] T9049;
  wire[3:0] T9050;
  wire T9051;
  wire[3:0] T9052;
  wire T9053;
  wire T9054;
  wire T9055;
  wire[3:0] T9056;
  wire[3:0] T9057;
  wire[3:0] T9058;
  wire T9059;
  wire[3:0] T9060;
  wire T9061;
  wire T9062;
  wire[3:0] T9063;
  wire[3:0] T9064;
  wire T9065;
  wire[3:0] T9066;
  wire T9067;
  wire T9068;
  wire T9069;
  wire T9070;
  wire T9071;
  wire[3:0] T9072;
  wire[3:0] T9073;
  wire[3:0] T9074;
  wire[3:0] T9075;
  wire[3:0] T9076;
  wire T9077;
  wire[3:0] T9078;
  wire T9079;
  wire T9080;
  wire[3:0] T9081;
  wire[3:0] T9082;
  wire T9083;
  wire[3:0] T9084;
  wire T9085;
  wire T9086;
  wire T9087;
  wire[3:0] T9088;
  wire[3:0] T9089;
  wire[3:0] T9090;
  wire T9091;
  wire[3:0] T9092;
  wire T9093;
  wire T9094;
  wire[3:0] T9095;
  wire[3:0] T9096;
  wire T9097;
  wire[3:0] T9098;
  wire T9099;
  wire T9100;
  wire T9101;
  wire T9102;
  wire[3:0] T9103;
  wire[3:0] T9104;
  wire[3:0] T9105;
  wire[3:0] T9106;
  wire T9107;
  wire[3:0] T9108;
  wire T9109;
  wire T9110;
  wire[3:0] T9111;
  wire[3:0] T9112;
  wire T9113;
  wire[3:0] T9114;
  wire T9115;
  wire T9116;
  wire T9117;
  wire[3:0] T9118;
  wire[3:0] T9119;
  wire[3:0] T9120;
  wire T9121;
  wire[3:0] T9122;
  wire T9123;
  wire T9124;
  wire[3:0] T9125;
  wire[3:0] T9126;
  wire T9127;
  wire[3:0] T9128;
  wire T9129;
  wire T9130;
  wire T9131;
  wire T9132;
  wire T9133;
  wire T9134;
  wire[3:0] T9135;
  wire[3:0] T9136;
  wire[3:0] T9137;
  wire[3:0] T9138;
  wire[3:0] T9139;
  wire[3:0] T9140;
  wire T9141;
  wire[3:0] T9142;
  wire T9143;
  wire T9144;
  wire[3:0] T9145;
  wire[3:0] T9146;
  wire T9147;
  wire[3:0] T9148;
  wire T9149;
  wire T9150;
  wire T9151;
  wire[3:0] T9152;
  wire[3:0] T9153;
  wire[3:0] T9154;
  wire T9155;
  wire[3:0] T9156;
  wire T9157;
  wire T9158;
  wire[3:0] T9159;
  wire[3:0] T9160;
  wire T9161;
  wire[3:0] T9162;
  wire T9163;
  wire T9164;
  wire T9165;
  wire T9166;
  wire[3:0] T9167;
  wire[3:0] T9168;
  wire[3:0] T9169;
  wire[3:0] T9170;
  wire T9171;
  wire[3:0] T9172;
  wire T9173;
  wire T9174;
  wire[3:0] T9175;
  wire[3:0] T9176;
  wire T9177;
  wire[3:0] T9178;
  wire T9179;
  wire T9180;
  wire T9181;
  wire[3:0] T9182;
  wire[3:0] T9183;
  wire[3:0] T9184;
  wire T9185;
  wire[3:0] T9186;
  wire T9187;
  wire T9188;
  wire[3:0] T9189;
  wire[3:0] T9190;
  wire T9191;
  wire[3:0] T9192;
  wire T9193;
  wire T9194;
  wire T9195;
  wire T9196;
  wire T9197;
  wire[3:0] T9198;
  wire[3:0] T9199;
  wire[3:0] T9200;
  wire[3:0] T9201;
  wire[3:0] T9202;
  wire T9203;
  wire[3:0] T9204;
  wire T9205;
  wire T9206;
  wire[3:0] T9207;
  wire[3:0] T9208;
  wire T9209;
  wire[3:0] T9210;
  wire T9211;
  wire T9212;
  wire T9213;
  wire[3:0] T9214;
  wire[3:0] T9215;
  wire[3:0] T9216;
  wire T9217;
  wire[3:0] T9218;
  wire T9219;
  wire T9220;
  wire[3:0] T9221;
  wire[3:0] T9222;
  wire T9223;
  wire[3:0] T9224;
  wire T9225;
  wire T9226;
  wire T9227;
  wire T9228;
  wire[3:0] T9229;
  wire[3:0] T9230;
  wire[3:0] T9231;
  wire[3:0] T9232;
  wire T9233;
  wire[3:0] T9234;
  wire T9235;
  wire T9236;
  wire[3:0] T9237;
  wire[3:0] T9238;
  wire T9239;
  wire[3:0] T9240;
  wire T9241;
  wire T9242;
  wire T9243;
  wire[3:0] T9244;
  wire[3:0] T9245;
  wire[3:0] T9246;
  wire T9247;
  wire[3:0] T9248;
  wire T9249;
  wire T9250;
  wire[3:0] T9251;
  wire[3:0] T9252;
  wire T9253;
  wire[3:0] T9254;
  wire T9255;
  wire T9256;
  wire T9257;
  wire T9258;
  wire T9259;
  wire T9260;
  wire T9261;
  wire T9262;
  wire T9263;
  wire[3:0] T9264;
  wire[3:0] T9265;
  wire[3:0] T9266;
  wire[3:0] T9267;
  wire[3:0] T9268;
  wire[3:0] T9269;
  wire[3:0] T9270;
  wire[3:0] T9271;
  wire[3:0] T9272;
  wire T9273;
  wire[3:0] T9274;
  wire T9275;
  wire T9276;
  wire[3:0] T9277;
  wire[3:0] T9278;
  wire T9279;
  wire[3:0] T9280;
  wire T9281;
  wire T9282;
  wire T9283;
  wire[3:0] T9284;
  wire[3:0] T9285;
  wire[3:0] T9286;
  wire T9287;
  wire[3:0] T9288;
  wire T9289;
  wire T9290;
  wire[3:0] T9291;
  wire[3:0] T9292;
  wire T9293;
  wire[3:0] T9294;
  wire T9295;
  wire T9296;
  wire T9297;
  wire T9298;
  wire[3:0] T9299;
  wire[3:0] T9300;
  wire[3:0] T9301;
  wire[3:0] T9302;
  wire T9303;
  wire[3:0] T9304;
  wire T9305;
  wire T9306;
  wire[3:0] T9307;
  wire[3:0] T9308;
  wire T9309;
  wire[3:0] T9310;
  wire T9311;
  wire T9312;
  wire T9313;
  wire[3:0] T9314;
  wire[3:0] T9315;
  wire[3:0] T9316;
  wire T9317;
  wire[3:0] T9318;
  wire T9319;
  wire T9320;
  wire[3:0] T9321;
  wire[3:0] T9322;
  wire T9323;
  wire[3:0] T9324;
  wire T9325;
  wire T9326;
  wire T9327;
  wire T9328;
  wire T9329;
  wire[3:0] T9330;
  wire[3:0] T9331;
  wire[3:0] T9332;
  wire[3:0] T9333;
  wire[3:0] T9334;
  wire T9335;
  wire[3:0] T9336;
  wire T9337;
  wire T9338;
  wire[3:0] T9339;
  wire[3:0] T9340;
  wire T9341;
  wire[3:0] T9342;
  wire T9343;
  wire T9344;
  wire T9345;
  wire[3:0] T9346;
  wire[3:0] T9347;
  wire[3:0] T9348;
  wire T9349;
  wire[3:0] T9350;
  wire T9351;
  wire T9352;
  wire[3:0] T9353;
  wire[3:0] T9354;
  wire T9355;
  wire[3:0] T9356;
  wire T9357;
  wire T9358;
  wire T9359;
  wire T9360;
  wire[3:0] T9361;
  wire[3:0] T9362;
  wire[3:0] T9363;
  wire[3:0] T9364;
  wire T9365;
  wire[3:0] T9366;
  wire T9367;
  wire T9368;
  wire[3:0] T9369;
  wire[3:0] T9370;
  wire T9371;
  wire[3:0] T9372;
  wire T9373;
  wire T9374;
  wire T9375;
  wire[3:0] T9376;
  wire[3:0] T9377;
  wire[3:0] T9378;
  wire T9379;
  wire[3:0] T9380;
  wire T9381;
  wire T9382;
  wire[3:0] T9383;
  wire[3:0] T9384;
  wire T9385;
  wire[3:0] T9386;
  wire T9387;
  wire T9388;
  wire T9389;
  wire T9390;
  wire T9391;
  wire T9392;
  wire[3:0] T9393;
  wire[3:0] T9394;
  wire[3:0] T9395;
  wire[3:0] T9396;
  wire[3:0] T9397;
  wire[3:0] T9398;
  wire T9399;
  wire[3:0] T9400;
  wire T9401;
  wire T9402;
  wire[3:0] T9403;
  wire[3:0] T9404;
  wire T9405;
  wire[3:0] T9406;
  wire T9407;
  wire T9408;
  wire T9409;
  wire[3:0] T9410;
  wire[3:0] T9411;
  wire[3:0] T9412;
  wire T9413;
  wire[3:0] T9414;
  wire T9415;
  wire T9416;
  wire[3:0] T9417;
  wire[3:0] T9418;
  wire T9419;
  wire[3:0] T9420;
  wire T9421;
  wire T9422;
  wire T9423;
  wire T9424;
  wire[3:0] T9425;
  wire[3:0] T9426;
  wire[3:0] T9427;
  wire[3:0] T9428;
  wire T9429;
  wire[3:0] T9430;
  wire T9431;
  wire T9432;
  wire[3:0] T9433;
  wire[3:0] T9434;
  wire T9435;
  wire[3:0] T9436;
  wire T9437;
  wire T9438;
  wire T9439;
  wire[3:0] T9440;
  wire[3:0] T9441;
  wire[3:0] T9442;
  wire T9443;
  wire[3:0] T9444;
  wire T9445;
  wire T9446;
  wire[3:0] T9447;
  wire[3:0] T9448;
  wire T9449;
  wire[3:0] T9450;
  wire T9451;
  wire T9452;
  wire T9453;
  wire T9454;
  wire T9455;
  wire[3:0] T9456;
  wire[3:0] T9457;
  wire[3:0] T9458;
  wire[3:0] T9459;
  wire[3:0] T9460;
  wire T9461;
  wire[3:0] T9462;
  wire T9463;
  wire T9464;
  wire[3:0] T9465;
  wire[3:0] T9466;
  wire T9467;
  wire[3:0] T9468;
  wire T9469;
  wire T9470;
  wire T9471;
  wire[3:0] T9472;
  wire[3:0] T9473;
  wire[3:0] T9474;
  wire T9475;
  wire[3:0] T9476;
  wire T9477;
  wire T9478;
  wire[3:0] T9479;
  wire[3:0] T9480;
  wire T9481;
  wire[3:0] T9482;
  wire T9483;
  wire T9484;
  wire T9485;
  wire T9486;
  wire[3:0] T9487;
  wire[3:0] T9488;
  wire[3:0] T9489;
  wire[3:0] T9490;
  wire T9491;
  wire[3:0] T9492;
  wire T9493;
  wire T9494;
  wire[3:0] T9495;
  wire[3:0] T9496;
  wire T9497;
  wire[3:0] T9498;
  wire T9499;
  wire T9500;
  wire T9501;
  wire[3:0] T9502;
  wire[3:0] T9503;
  wire[3:0] T9504;
  wire T9505;
  wire[3:0] T9506;
  wire T9507;
  wire T9508;
  wire[3:0] T9509;
  wire[3:0] T9510;
  wire T9511;
  wire[3:0] T9512;
  wire T9513;
  wire T9514;
  wire T9515;
  wire T9516;
  wire T9517;
  wire T9518;
  wire T9519;
  wire[3:0] T9520;
  wire[3:0] T9521;
  wire[3:0] T9522;
  wire[3:0] T9523;
  wire[3:0] T9524;
  wire[3:0] T9525;
  wire[3:0] T9526;
  wire T9527;
  wire[3:0] T9528;
  wire T9529;
  wire T9530;
  wire[3:0] T9531;
  wire[3:0] T9532;
  wire T9533;
  wire[3:0] T9534;
  wire T9535;
  wire T9536;
  wire T9537;
  wire[3:0] T9538;
  wire[3:0] T9539;
  wire[3:0] T9540;
  wire T9541;
  wire[3:0] T9542;
  wire T9543;
  wire T9544;
  wire[3:0] T9545;
  wire[3:0] T9546;
  wire T9547;
  wire[3:0] T9548;
  wire T9549;
  wire T9550;
  wire T9551;
  wire T9552;
  wire[3:0] T9553;
  wire[3:0] T9554;
  wire[3:0] T9555;
  wire[3:0] T9556;
  wire T9557;
  wire[3:0] T9558;
  wire T9559;
  wire T9560;
  wire[3:0] T9561;
  wire[3:0] T9562;
  wire T9563;
  wire[3:0] T9564;
  wire T9565;
  wire T9566;
  wire T9567;
  wire[3:0] T9568;
  wire[3:0] T9569;
  wire[3:0] T9570;
  wire T9571;
  wire[3:0] T9572;
  wire T9573;
  wire T9574;
  wire[3:0] T9575;
  wire[3:0] T9576;
  wire T9577;
  wire[3:0] T9578;
  wire T9579;
  wire T9580;
  wire T9581;
  wire T9582;
  wire T9583;
  wire[3:0] T9584;
  wire[3:0] T9585;
  wire[3:0] T9586;
  wire[3:0] T9587;
  wire[3:0] T9588;
  wire T9589;
  wire[3:0] T9590;
  wire T9591;
  wire T9592;
  wire[3:0] T9593;
  wire[3:0] T9594;
  wire T9595;
  wire[3:0] T9596;
  wire T9597;
  wire T9598;
  wire T9599;
  wire[3:0] T9600;
  wire[3:0] T9601;
  wire[3:0] T9602;
  wire T9603;
  wire[3:0] T9604;
  wire T9605;
  wire T9606;
  wire[3:0] T9607;
  wire[3:0] T9608;
  wire T9609;
  wire[3:0] T9610;
  wire T9611;
  wire T9612;
  wire T9613;
  wire T9614;
  wire[3:0] T9615;
  wire[3:0] T9616;
  wire[3:0] T9617;
  wire[3:0] T9618;
  wire T9619;
  wire[3:0] T9620;
  wire T9621;
  wire T9622;
  wire[3:0] T9623;
  wire[3:0] T9624;
  wire T9625;
  wire[3:0] T9626;
  wire T9627;
  wire T9628;
  wire T9629;
  wire[3:0] T9630;
  wire[3:0] T9631;
  wire[3:0] T9632;
  wire T9633;
  wire[3:0] T9634;
  wire T9635;
  wire T9636;
  wire[3:0] T9637;
  wire[3:0] T9638;
  wire T9639;
  wire[3:0] T9640;
  wire T9641;
  wire T9642;
  wire T9643;
  wire T9644;
  wire T9645;
  wire T9646;
  wire[3:0] T9647;
  wire[3:0] T9648;
  wire[3:0] T9649;
  wire[3:0] T9650;
  wire[3:0] T9651;
  wire[3:0] T9652;
  wire T9653;
  wire[3:0] T9654;
  wire T9655;
  wire T9656;
  wire[3:0] T9657;
  wire[3:0] T9658;
  wire T9659;
  wire[3:0] T9660;
  wire T9661;
  wire T9662;
  wire T9663;
  wire[3:0] T9664;
  wire[3:0] T9665;
  wire[3:0] T9666;
  wire T9667;
  wire[3:0] T9668;
  wire T9669;
  wire T9670;
  wire[3:0] T9671;
  wire[3:0] T9672;
  wire T9673;
  wire[3:0] T9674;
  wire T9675;
  wire T9676;
  wire T9677;
  wire T9678;
  wire[3:0] T9679;
  wire[3:0] T9680;
  wire[3:0] T9681;
  wire[3:0] T9682;
  wire T9683;
  wire[3:0] T9684;
  wire T9685;
  wire T9686;
  wire[3:0] T9687;
  wire[3:0] T9688;
  wire T9689;
  wire[3:0] T9690;
  wire T9691;
  wire T9692;
  wire T9693;
  wire[3:0] T9694;
  wire[3:0] T9695;
  wire[3:0] T9696;
  wire T9697;
  wire[3:0] T9698;
  wire T9699;
  wire T9700;
  wire[3:0] T9701;
  wire[3:0] T9702;
  wire T9703;
  wire[3:0] T9704;
  wire T9705;
  wire T9706;
  wire T9707;
  wire T9708;
  wire T9709;
  wire[3:0] T9710;
  wire[3:0] T9711;
  wire[3:0] T9712;
  wire[3:0] T9713;
  wire[3:0] T9714;
  wire T9715;
  wire[3:0] T9716;
  wire T9717;
  wire T9718;
  wire[3:0] T9719;
  wire[3:0] T9720;
  wire T9721;
  wire[3:0] T9722;
  wire T9723;
  wire T9724;
  wire T9725;
  wire[3:0] T9726;
  wire[3:0] T9727;
  wire[3:0] T9728;
  wire T9729;
  wire[3:0] T9730;
  wire T9731;
  wire T9732;
  wire[3:0] T9733;
  wire[3:0] T9734;
  wire T9735;
  wire[3:0] T9736;
  wire T9737;
  wire T9738;
  wire T9739;
  wire T9740;
  wire[3:0] T9741;
  wire[3:0] T9742;
  wire[3:0] T9743;
  wire[3:0] T9744;
  wire T9745;
  wire[3:0] T9746;
  wire T9747;
  wire T9748;
  wire[3:0] T9749;
  wire[3:0] T9750;
  wire T9751;
  wire[3:0] T9752;
  wire T9753;
  wire T9754;
  wire T9755;
  wire[3:0] T9756;
  wire[3:0] T9757;
  wire[3:0] T9758;
  wire T9759;
  wire[3:0] T9760;
  wire T9761;
  wire T9762;
  wire[3:0] T9763;
  wire[3:0] T9764;
  wire T9765;
  wire[3:0] T9766;
  wire T9767;
  wire T9768;
  wire T9769;
  wire T9770;
  wire T9771;
  wire T9772;
  wire T9773;
  wire T9774;
  wire[3:0] T9775;
  wire[3:0] T9776;
  wire[3:0] T9777;
  wire[3:0] T9778;
  wire[3:0] T9779;
  wire[3:0] T9780;
  wire[3:0] T9781;
  wire[3:0] T9782;
  wire T9783;
  wire[3:0] T9784;
  wire T9785;
  wire T9786;
  wire[3:0] T9787;
  wire[3:0] T9788;
  wire T9789;
  wire[3:0] T9790;
  wire T9791;
  wire T9792;
  wire T9793;
  wire[3:0] T9794;
  wire[3:0] T9795;
  wire[3:0] T9796;
  wire T9797;
  wire[3:0] T9798;
  wire T9799;
  wire T9800;
  wire[3:0] T9801;
  wire[3:0] T9802;
  wire T9803;
  wire[3:0] T9804;
  wire T9805;
  wire T9806;
  wire T9807;
  wire T9808;
  wire[3:0] T9809;
  wire[3:0] T9810;
  wire[3:0] T9811;
  wire[3:0] T9812;
  wire T9813;
  wire[3:0] T9814;
  wire T9815;
  wire T9816;
  wire[3:0] T9817;
  wire[3:0] T9818;
  wire T9819;
  wire[3:0] T9820;
  wire T9821;
  wire T9822;
  wire T9823;
  wire[3:0] T9824;
  wire[3:0] T9825;
  wire[3:0] T9826;
  wire T9827;
  wire[3:0] T9828;
  wire T9829;
  wire T9830;
  wire[3:0] T9831;
  wire[3:0] T9832;
  wire T9833;
  wire[3:0] T9834;
  wire T9835;
  wire T9836;
  wire T9837;
  wire T9838;
  wire T9839;
  wire[3:0] T9840;
  wire[3:0] T9841;
  wire[3:0] T9842;
  wire[3:0] T9843;
  wire[3:0] T9844;
  wire T9845;
  wire[3:0] T9846;
  wire T9847;
  wire T9848;
  wire[3:0] T9849;
  wire[3:0] T9850;
  wire T9851;
  wire[3:0] T9852;
  wire T9853;
  wire T9854;
  wire T9855;
  wire[3:0] T9856;
  wire[3:0] T9857;
  wire[3:0] T9858;
  wire T9859;
  wire[3:0] T9860;
  wire T9861;
  wire T9862;
  wire[3:0] T9863;
  wire[3:0] T9864;
  wire T9865;
  wire[3:0] T9866;
  wire T9867;
  wire T9868;
  wire T9869;
  wire T9870;
  wire[3:0] T9871;
  wire[3:0] T9872;
  wire[3:0] T9873;
  wire[3:0] T9874;
  wire T9875;
  wire[3:0] T9876;
  wire T9877;
  wire T9878;
  wire[3:0] T9879;
  wire[3:0] T9880;
  wire T9881;
  wire[3:0] T9882;
  wire T9883;
  wire T9884;
  wire T9885;
  wire[3:0] T9886;
  wire[3:0] T9887;
  wire[3:0] T9888;
  wire T9889;
  wire[3:0] T9890;
  wire T9891;
  wire T9892;
  wire[3:0] T9893;
  wire[3:0] T9894;
  wire T9895;
  wire[3:0] T9896;
  wire T9897;
  wire T9898;
  wire T9899;
  wire T9900;
  wire T9901;
  wire T9902;
  wire[3:0] T9903;
  wire[3:0] T9904;
  wire[3:0] T9905;
  wire[3:0] T9906;
  wire[3:0] T9907;
  wire[3:0] T9908;
  wire T9909;
  wire[3:0] T9910;
  wire T9911;
  wire T9912;
  wire[3:0] T9913;
  wire[3:0] T9914;
  wire T9915;
  wire[3:0] T9916;
  wire T9917;
  wire T9918;
  wire T9919;
  wire[3:0] T9920;
  wire[3:0] T9921;
  wire[3:0] T9922;
  wire T9923;
  wire[3:0] T9924;
  wire T9925;
  wire T9926;
  wire[3:0] T9927;
  wire[3:0] T9928;
  wire T9929;
  wire[3:0] T9930;
  wire T9931;
  wire T9932;
  wire T9933;
  wire T9934;
  wire[3:0] T9935;
  wire[3:0] T9936;
  wire[3:0] T9937;
  wire[3:0] T9938;
  wire T9939;
  wire[3:0] T9940;
  wire T9941;
  wire T9942;
  wire[3:0] T9943;
  wire[3:0] T9944;
  wire T9945;
  wire[3:0] T9946;
  wire T9947;
  wire T9948;
  wire T9949;
  wire[3:0] T9950;
  wire[3:0] T9951;
  wire[3:0] T9952;
  wire T9953;
  wire[3:0] T9954;
  wire T9955;
  wire T9956;
  wire[3:0] T9957;
  wire[3:0] T9958;
  wire T9959;
  wire[3:0] T9960;
  wire T9961;
  wire T9962;
  wire T9963;
  wire T9964;
  wire T9965;
  wire[3:0] T9966;
  wire[3:0] T9967;
  wire[3:0] T9968;
  wire[3:0] T9969;
  wire[3:0] T9970;
  wire T9971;
  wire[3:0] T9972;
  wire T9973;
  wire T9974;
  wire[3:0] T9975;
  wire[3:0] T9976;
  wire T9977;
  wire[3:0] T9978;
  wire T9979;
  wire T9980;
  wire T9981;
  wire[3:0] T9982;
  wire[3:0] T9983;
  wire[3:0] T9984;
  wire T9985;
  wire[3:0] T9986;
  wire T9987;
  wire T9988;
  wire[3:0] T9989;
  wire[3:0] T9990;
  wire T9991;
  wire[3:0] T9992;
  wire T9993;
  wire T9994;
  wire T9995;
  wire T9996;
  wire[3:0] T9997;
  wire[3:0] T9998;
  wire[3:0] T9999;
  wire[3:0] T10000;
  wire T10001;
  wire[3:0] T10002;
  wire T10003;
  wire T10004;
  wire[3:0] T10005;
  wire[3:0] T10006;
  wire T10007;
  wire[3:0] T10008;
  wire T10009;
  wire T10010;
  wire T10011;
  wire[3:0] T10012;
  wire[3:0] T10013;
  wire[3:0] T10014;
  wire T10015;
  wire[3:0] T10016;
  wire T10017;
  wire T10018;
  wire[3:0] T10019;
  wire[3:0] T10020;
  wire T10021;
  wire[3:0] T10022;
  wire T10023;
  wire T10024;
  wire T10025;
  wire T10026;
  wire T10027;
  wire T10028;
  wire T10029;
  wire[3:0] T10030;
  wire[3:0] T10031;
  wire[3:0] T10032;
  wire[3:0] T10033;
  wire[3:0] T10034;
  wire[3:0] T10035;
  wire[3:0] T10036;
  wire T10037;
  wire[3:0] T10038;
  wire T10039;
  wire T10040;
  wire[3:0] T10041;
  wire[3:0] T10042;
  wire T10043;
  wire[3:0] T10044;
  wire T10045;
  wire T10046;
  wire T10047;
  wire[3:0] T10048;
  wire[3:0] T10049;
  wire[3:0] T10050;
  wire T10051;
  wire[3:0] T10052;
  wire T10053;
  wire T10054;
  wire[3:0] T10055;
  wire[3:0] T10056;
  wire T10057;
  wire[3:0] T10058;
  wire T10059;
  wire T10060;
  wire T10061;
  wire T10062;
  wire[3:0] T10063;
  wire[3:0] T10064;
  wire[3:0] T10065;
  wire[3:0] T10066;
  wire T10067;
  wire[3:0] T10068;
  wire T10069;
  wire T10070;
  wire[3:0] T10071;
  wire[3:0] T10072;
  wire T10073;
  wire[3:0] T10074;
  wire T10075;
  wire T10076;
  wire T10077;
  wire[3:0] T10078;
  wire[3:0] T10079;
  wire[3:0] T10080;
  wire T10081;
  wire[3:0] T10082;
  wire T10083;
  wire T10084;
  wire[3:0] T10085;
  wire[3:0] T10086;
  wire T10087;
  wire[3:0] T10088;
  wire T10089;
  wire T10090;
  wire T10091;
  wire T10092;
  wire T10093;
  wire[3:0] T10094;
  wire[3:0] T10095;
  wire[3:0] T10096;
  wire[3:0] T10097;
  wire[3:0] T10098;
  wire T10099;
  wire[3:0] T10100;
  wire T10101;
  wire T10102;
  wire[3:0] T10103;
  wire[3:0] T10104;
  wire T10105;
  wire[3:0] T10106;
  wire T10107;
  wire T10108;
  wire T10109;
  wire[3:0] T10110;
  wire[3:0] T10111;
  wire[3:0] T10112;
  wire T10113;
  wire[3:0] T10114;
  wire T10115;
  wire T10116;
  wire[3:0] T10117;
  wire[3:0] T10118;
  wire T10119;
  wire[3:0] T10120;
  wire T10121;
  wire T10122;
  wire T10123;
  wire T10124;
  wire[3:0] T10125;
  wire[3:0] T10126;
  wire[3:0] T10127;
  wire[3:0] T10128;
  wire T10129;
  wire[3:0] T10130;
  wire T10131;
  wire T10132;
  wire[3:0] T10133;
  wire[3:0] T10134;
  wire T10135;
  wire[3:0] T10136;
  wire T10137;
  wire T10138;
  wire T10139;
  wire[3:0] T10140;
  wire[3:0] T10141;
  wire[3:0] T10142;
  wire T10143;
  wire[3:0] T10144;
  wire T10145;
  wire T10146;
  wire[3:0] T10147;
  wire[3:0] T10148;
  wire T10149;
  wire[3:0] T10150;
  wire T10151;
  wire T10152;
  wire T10153;
  wire T10154;
  wire T10155;
  wire T10156;
  wire[3:0] T10157;
  wire[3:0] T10158;
  wire[3:0] T10159;
  wire[3:0] T10160;
  wire[3:0] T10161;
  wire[3:0] T10162;
  wire T10163;
  wire[3:0] T10164;
  wire T10165;
  wire T10166;
  wire[3:0] T10167;
  wire[3:0] T10168;
  wire T10169;
  wire[3:0] T10170;
  wire T10171;
  wire T10172;
  wire T10173;
  wire[3:0] T10174;
  wire[3:0] T10175;
  wire[3:0] T10176;
  wire T10177;
  wire[3:0] T10178;
  wire T10179;
  wire T10180;
  wire[3:0] T10181;
  wire[3:0] T10182;
  wire T10183;
  wire[3:0] T10184;
  wire T10185;
  wire T10186;
  wire T10187;
  wire T10188;
  wire[3:0] T10189;
  wire[3:0] T10190;
  wire[3:0] T10191;
  wire[3:0] T10192;
  wire T10193;
  wire[3:0] T10194;
  wire T10195;
  wire T10196;
  wire[3:0] T10197;
  wire[3:0] T10198;
  wire T10199;
  wire[3:0] T10200;
  wire T10201;
  wire T10202;
  wire T10203;
  wire[3:0] T10204;
  wire[3:0] T10205;
  wire[3:0] T10206;
  wire T10207;
  wire[3:0] T10208;
  wire T10209;
  wire T10210;
  wire[3:0] T10211;
  wire[3:0] T10212;
  wire T10213;
  wire[3:0] T10214;
  wire T10215;
  wire T10216;
  wire T10217;
  wire T10218;
  wire T10219;
  wire[3:0] T10220;
  wire[3:0] T10221;
  wire[3:0] T10222;
  wire[3:0] T10223;
  wire[3:0] T10224;
  wire T10225;
  wire[3:0] T10226;
  wire T10227;
  wire T10228;
  wire[3:0] T10229;
  wire[3:0] T10230;
  wire T10231;
  wire[3:0] T10232;
  wire T10233;
  wire T10234;
  wire T10235;
  wire[3:0] T10236;
  wire[3:0] T10237;
  wire[3:0] T10238;
  wire T10239;
  wire[3:0] T10240;
  wire T10241;
  wire T10242;
  wire[3:0] T10243;
  wire[3:0] T10244;
  wire T10245;
  wire[3:0] T10246;
  wire T10247;
  wire T10248;
  wire T10249;
  wire T10250;
  wire[3:0] T10251;
  wire[3:0] T10252;
  wire[3:0] T10253;
  wire[3:0] T10254;
  wire T10255;
  wire[3:0] T10256;
  wire T10257;
  wire T10258;
  wire[3:0] T10259;
  wire[3:0] T10260;
  wire T10261;
  wire[3:0] T10262;
  wire T10263;
  wire T10264;
  wire T10265;
  wire[3:0] T10266;
  wire[3:0] T10267;
  wire[3:0] T10268;
  wire T10269;
  wire[3:0] T10270;
  wire T10271;
  wire T10272;
  wire[3:0] T10273;
  wire[3:0] T10274;
  wire T10275;
  wire[3:0] T10276;
  wire T10277;
  wire T10278;
  wire T10279;
  wire T10280;
  wire T10281;
  wire T10282;
  wire T10283;
  wire T10284;
  wire T10285;
  wire T10286;
  wire T10287;
  wire T10288;
  wire T10289;
  wire T10290;
  wire T10291;
  wire T10292;
  wire T10293;
  wire T10294;
  wire T10295;
  wire T10296;
  wire T10297;
  wire T10298;
  wire T10299;
  reg  delayCount;
  wire T10300;
  wire T10301;
  wire T10302;
  wire T10303;
  wire T10304;
  wire T10305;
  wire T10306;
  wire T10307;
  wire T10308;
  wire T10309;
  wire T10310;
  wire T10311;
  wire T10312;
  wire T10313;
  wire T10314;
  wire T10315;
  wire T10316;
  wire T10317;
  wire T10318;
  wire T10319;
  wire T10320;
  wire T10321;
  wire reachedEnd;
  wire T10322;
  wire[5:0] wordLen;
  reg [5:0] delayedIndex;
  reg [5:0] R10323;
  reg [5:0] index;
  wire[5:0] T10324;
  wire[5:0] T10325;
  wire[5:0] T10326;
  wire[5:0] T10327;
  wire[5:0] T10328;
  wire T10329;
  wire T10330;
  wire T10331;
  wire T10332;
  wire[5:0] T10333;
  wire T10334;
  wire[1:0] T10335;
  wire T10336;
  wire T10337;
  reg [3:0] curInfo_tag;
  wire[3:0] T10338;
  wire[3:0] curCount;
  wire T10339;
  wire T10340;
  wire T10341;
  wire[15:0] T10342;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    hashFound = {1{$random}};
    state = {1{$random}};
    curInfo_len = {1{$random}};
    checkFirst = {1{$random}};
    hashCount2 = {1{$random}};
    counts_0 = {1{$random}};
    curInfo_hash2 = {1{$random}};
    curInfo_hash1 = {1{$random}};
    counts_2 = {1{$random}};
    counts_3 = {1{$random}};
    counts_4 = {1{$random}};
    counts_5 = {1{$random}};
    counts_6 = {1{$random}};
    counts_7 = {1{$random}};
    counts_8 = {1{$random}};
    counts_9 = {1{$random}};
    counts_10 = {1{$random}};
    counts_11 = {1{$random}};
    counts_12 = {1{$random}};
    counts_13 = {1{$random}};
    counts_14 = {1{$random}};
    counts_15 = {1{$random}};
    counts_16 = {1{$random}};
    counts_17 = {1{$random}};
    counts_18 = {1{$random}};
    counts_19 = {1{$random}};
    counts_20 = {1{$random}};
    counts_21 = {1{$random}};
    counts_22 = {1{$random}};
    counts_23 = {1{$random}};
    counts_24 = {1{$random}};
    counts_25 = {1{$random}};
    counts_26 = {1{$random}};
    counts_27 = {1{$random}};
    counts_28 = {1{$random}};
    counts_29 = {1{$random}};
    counts_30 = {1{$random}};
    counts_31 = {1{$random}};
    counts_32 = {1{$random}};
    counts_33 = {1{$random}};
    counts_34 = {1{$random}};
    counts_35 = {1{$random}};
    counts_36 = {1{$random}};
    counts_37 = {1{$random}};
    counts_38 = {1{$random}};
    counts_39 = {1{$random}};
    counts_40 = {1{$random}};
    counts_41 = {1{$random}};
    counts_42 = {1{$random}};
    counts_43 = {1{$random}};
    counts_44 = {1{$random}};
    counts_45 = {1{$random}};
    counts_46 = {1{$random}};
    counts_47 = {1{$random}};
    counts_48 = {1{$random}};
    counts_49 = {1{$random}};
    counts_50 = {1{$random}};
    counts_51 = {1{$random}};
    counts_52 = {1{$random}};
    counts_53 = {1{$random}};
    counts_54 = {1{$random}};
    counts_55 = {1{$random}};
    counts_56 = {1{$random}};
    counts_57 = {1{$random}};
    counts_58 = {1{$random}};
    counts_59 = {1{$random}};
    counts_60 = {1{$random}};
    counts_61 = {1{$random}};
    counts_62 = {1{$random}};
    counts_63 = {1{$random}};
    counts_64 = {1{$random}};
    counts_65 = {1{$random}};
    counts_66 = {1{$random}};
    counts_67 = {1{$random}};
    counts_68 = {1{$random}};
    counts_69 = {1{$random}};
    counts_70 = {1{$random}};
    counts_71 = {1{$random}};
    counts_72 = {1{$random}};
    counts_73 = {1{$random}};
    counts_74 = {1{$random}};
    counts_75 = {1{$random}};
    counts_76 = {1{$random}};
    counts_77 = {1{$random}};
    counts_78 = {1{$random}};
    counts_79 = {1{$random}};
    counts_80 = {1{$random}};
    counts_81 = {1{$random}};
    counts_82 = {1{$random}};
    counts_83 = {1{$random}};
    counts_84 = {1{$random}};
    counts_85 = {1{$random}};
    counts_86 = {1{$random}};
    counts_87 = {1{$random}};
    counts_88 = {1{$random}};
    counts_89 = {1{$random}};
    counts_90 = {1{$random}};
    counts_91 = {1{$random}};
    counts_92 = {1{$random}};
    counts_93 = {1{$random}};
    counts_94 = {1{$random}};
    counts_95 = {1{$random}};
    counts_96 = {1{$random}};
    counts_97 = {1{$random}};
    counts_98 = {1{$random}};
    counts_99 = {1{$random}};
    counts_100 = {1{$random}};
    counts_101 = {1{$random}};
    counts_102 = {1{$random}};
    counts_103 = {1{$random}};
    counts_104 = {1{$random}};
    counts_105 = {1{$random}};
    counts_106 = {1{$random}};
    counts_107 = {1{$random}};
    counts_108 = {1{$random}};
    counts_109 = {1{$random}};
    counts_110 = {1{$random}};
    counts_111 = {1{$random}};
    counts_112 = {1{$random}};
    counts_113 = {1{$random}};
    counts_114 = {1{$random}};
    counts_115 = {1{$random}};
    counts_116 = {1{$random}};
    counts_117 = {1{$random}};
    counts_118 = {1{$random}};
    counts_119 = {1{$random}};
    counts_120 = {1{$random}};
    counts_121 = {1{$random}};
    counts_122 = {1{$random}};
    counts_123 = {1{$random}};
    counts_124 = {1{$random}};
    counts_125 = {1{$random}};
    counts_126 = {1{$random}};
    counts_127 = {1{$random}};
    counts_128 = {1{$random}};
    counts_129 = {1{$random}};
    counts_130 = {1{$random}};
    counts_131 = {1{$random}};
    counts_132 = {1{$random}};
    counts_133 = {1{$random}};
    counts_134 = {1{$random}};
    counts_135 = {1{$random}};
    counts_136 = {1{$random}};
    counts_137 = {1{$random}};
    counts_138 = {1{$random}};
    counts_139 = {1{$random}};
    counts_140 = {1{$random}};
    counts_141 = {1{$random}};
    counts_142 = {1{$random}};
    counts_143 = {1{$random}};
    counts_144 = {1{$random}};
    counts_145 = {1{$random}};
    counts_146 = {1{$random}};
    counts_147 = {1{$random}};
    counts_148 = {1{$random}};
    counts_149 = {1{$random}};
    counts_150 = {1{$random}};
    counts_151 = {1{$random}};
    counts_152 = {1{$random}};
    counts_153 = {1{$random}};
    counts_154 = {1{$random}};
    counts_155 = {1{$random}};
    counts_156 = {1{$random}};
    counts_157 = {1{$random}};
    counts_158 = {1{$random}};
    counts_159 = {1{$random}};
    counts_160 = {1{$random}};
    counts_161 = {1{$random}};
    counts_162 = {1{$random}};
    counts_163 = {1{$random}};
    counts_164 = {1{$random}};
    counts_165 = {1{$random}};
    counts_166 = {1{$random}};
    counts_167 = {1{$random}};
    counts_168 = {1{$random}};
    counts_169 = {1{$random}};
    counts_170 = {1{$random}};
    counts_171 = {1{$random}};
    counts_172 = {1{$random}};
    counts_173 = {1{$random}};
    counts_174 = {1{$random}};
    counts_175 = {1{$random}};
    counts_176 = {1{$random}};
    counts_177 = {1{$random}};
    counts_178 = {1{$random}};
    counts_179 = {1{$random}};
    counts_180 = {1{$random}};
    counts_181 = {1{$random}};
    counts_182 = {1{$random}};
    counts_183 = {1{$random}};
    counts_184 = {1{$random}};
    counts_185 = {1{$random}};
    counts_186 = {1{$random}};
    counts_187 = {1{$random}};
    counts_188 = {1{$random}};
    counts_189 = {1{$random}};
    counts_190 = {1{$random}};
    counts_191 = {1{$random}};
    counts_192 = {1{$random}};
    counts_193 = {1{$random}};
    counts_194 = {1{$random}};
    counts_195 = {1{$random}};
    counts_196 = {1{$random}};
    counts_197 = {1{$random}};
    counts_198 = {1{$random}};
    counts_199 = {1{$random}};
    counts_200 = {1{$random}};
    counts_201 = {1{$random}};
    counts_202 = {1{$random}};
    counts_203 = {1{$random}};
    counts_204 = {1{$random}};
    counts_205 = {1{$random}};
    counts_206 = {1{$random}};
    counts_207 = {1{$random}};
    counts_208 = {1{$random}};
    counts_209 = {1{$random}};
    counts_210 = {1{$random}};
    counts_211 = {1{$random}};
    counts_212 = {1{$random}};
    counts_213 = {1{$random}};
    counts_214 = {1{$random}};
    counts_215 = {1{$random}};
    counts_216 = {1{$random}};
    counts_217 = {1{$random}};
    counts_218 = {1{$random}};
    counts_219 = {1{$random}};
    counts_220 = {1{$random}};
    counts_221 = {1{$random}};
    counts_222 = {1{$random}};
    counts_223 = {1{$random}};
    counts_224 = {1{$random}};
    counts_225 = {1{$random}};
    counts_226 = {1{$random}};
    counts_227 = {1{$random}};
    counts_228 = {1{$random}};
    counts_229 = {1{$random}};
    counts_230 = {1{$random}};
    counts_231 = {1{$random}};
    counts_232 = {1{$random}};
    counts_233 = {1{$random}};
    counts_234 = {1{$random}};
    counts_235 = {1{$random}};
    counts_236 = {1{$random}};
    counts_237 = {1{$random}};
    counts_238 = {1{$random}};
    counts_239 = {1{$random}};
    counts_240 = {1{$random}};
    counts_241 = {1{$random}};
    counts_242 = {1{$random}};
    counts_243 = {1{$random}};
    counts_244 = {1{$random}};
    counts_245 = {1{$random}};
    counts_246 = {1{$random}};
    counts_247 = {1{$random}};
    counts_248 = {1{$random}};
    counts_249 = {1{$random}};
    counts_250 = {1{$random}};
    counts_251 = {1{$random}};
    counts_252 = {1{$random}};
    counts_253 = {1{$random}};
    counts_254 = {1{$random}};
    counts_255 = {1{$random}};
    counts_256 = {1{$random}};
    counts_257 = {1{$random}};
    counts_258 = {1{$random}};
    counts_259 = {1{$random}};
    counts_260 = {1{$random}};
    counts_261 = {1{$random}};
    counts_262 = {1{$random}};
    counts_263 = {1{$random}};
    counts_264 = {1{$random}};
    counts_265 = {1{$random}};
    counts_266 = {1{$random}};
    counts_267 = {1{$random}};
    counts_268 = {1{$random}};
    counts_269 = {1{$random}};
    counts_270 = {1{$random}};
    counts_271 = {1{$random}};
    counts_272 = {1{$random}};
    counts_273 = {1{$random}};
    counts_274 = {1{$random}};
    counts_275 = {1{$random}};
    counts_276 = {1{$random}};
    counts_277 = {1{$random}};
    counts_278 = {1{$random}};
    counts_279 = {1{$random}};
    counts_280 = {1{$random}};
    counts_281 = {1{$random}};
    counts_282 = {1{$random}};
    counts_283 = {1{$random}};
    counts_284 = {1{$random}};
    counts_285 = {1{$random}};
    counts_286 = {1{$random}};
    counts_287 = {1{$random}};
    counts_288 = {1{$random}};
    counts_289 = {1{$random}};
    counts_290 = {1{$random}};
    counts_291 = {1{$random}};
    counts_292 = {1{$random}};
    counts_293 = {1{$random}};
    counts_294 = {1{$random}};
    counts_295 = {1{$random}};
    counts_296 = {1{$random}};
    counts_297 = {1{$random}};
    counts_298 = {1{$random}};
    counts_299 = {1{$random}};
    counts_300 = {1{$random}};
    counts_301 = {1{$random}};
    counts_302 = {1{$random}};
    counts_303 = {1{$random}};
    counts_304 = {1{$random}};
    counts_305 = {1{$random}};
    counts_306 = {1{$random}};
    counts_307 = {1{$random}};
    counts_308 = {1{$random}};
    counts_309 = {1{$random}};
    counts_310 = {1{$random}};
    counts_311 = {1{$random}};
    counts_312 = {1{$random}};
    counts_313 = {1{$random}};
    counts_314 = {1{$random}};
    counts_315 = {1{$random}};
    counts_316 = {1{$random}};
    counts_317 = {1{$random}};
    counts_318 = {1{$random}};
    counts_319 = {1{$random}};
    counts_320 = {1{$random}};
    counts_321 = {1{$random}};
    counts_322 = {1{$random}};
    counts_323 = {1{$random}};
    counts_324 = {1{$random}};
    counts_325 = {1{$random}};
    counts_326 = {1{$random}};
    counts_327 = {1{$random}};
    counts_328 = {1{$random}};
    counts_329 = {1{$random}};
    counts_330 = {1{$random}};
    counts_331 = {1{$random}};
    counts_332 = {1{$random}};
    counts_333 = {1{$random}};
    counts_334 = {1{$random}};
    counts_335 = {1{$random}};
    counts_336 = {1{$random}};
    counts_337 = {1{$random}};
    counts_338 = {1{$random}};
    counts_339 = {1{$random}};
    counts_340 = {1{$random}};
    counts_341 = {1{$random}};
    counts_342 = {1{$random}};
    counts_343 = {1{$random}};
    counts_344 = {1{$random}};
    counts_345 = {1{$random}};
    counts_346 = {1{$random}};
    counts_347 = {1{$random}};
    counts_348 = {1{$random}};
    counts_349 = {1{$random}};
    counts_350 = {1{$random}};
    counts_351 = {1{$random}};
    counts_352 = {1{$random}};
    counts_353 = {1{$random}};
    counts_354 = {1{$random}};
    counts_355 = {1{$random}};
    counts_356 = {1{$random}};
    counts_357 = {1{$random}};
    counts_358 = {1{$random}};
    counts_359 = {1{$random}};
    counts_360 = {1{$random}};
    counts_361 = {1{$random}};
    counts_362 = {1{$random}};
    counts_363 = {1{$random}};
    counts_364 = {1{$random}};
    counts_365 = {1{$random}};
    counts_366 = {1{$random}};
    counts_367 = {1{$random}};
    counts_368 = {1{$random}};
    counts_369 = {1{$random}};
    counts_370 = {1{$random}};
    counts_371 = {1{$random}};
    counts_372 = {1{$random}};
    counts_373 = {1{$random}};
    counts_374 = {1{$random}};
    counts_375 = {1{$random}};
    counts_376 = {1{$random}};
    counts_377 = {1{$random}};
    counts_378 = {1{$random}};
    counts_379 = {1{$random}};
    counts_380 = {1{$random}};
    counts_381 = {1{$random}};
    counts_382 = {1{$random}};
    counts_383 = {1{$random}};
    counts_384 = {1{$random}};
    counts_385 = {1{$random}};
    counts_386 = {1{$random}};
    counts_387 = {1{$random}};
    counts_388 = {1{$random}};
    counts_389 = {1{$random}};
    counts_390 = {1{$random}};
    counts_391 = {1{$random}};
    counts_392 = {1{$random}};
    counts_393 = {1{$random}};
    counts_394 = {1{$random}};
    counts_395 = {1{$random}};
    counts_396 = {1{$random}};
    counts_397 = {1{$random}};
    counts_398 = {1{$random}};
    counts_399 = {1{$random}};
    counts_400 = {1{$random}};
    counts_401 = {1{$random}};
    counts_402 = {1{$random}};
    counts_403 = {1{$random}};
    counts_404 = {1{$random}};
    counts_405 = {1{$random}};
    counts_406 = {1{$random}};
    counts_407 = {1{$random}};
    counts_408 = {1{$random}};
    counts_409 = {1{$random}};
    counts_410 = {1{$random}};
    counts_411 = {1{$random}};
    counts_412 = {1{$random}};
    counts_413 = {1{$random}};
    counts_414 = {1{$random}};
    counts_415 = {1{$random}};
    counts_416 = {1{$random}};
    counts_417 = {1{$random}};
    counts_418 = {1{$random}};
    counts_419 = {1{$random}};
    counts_420 = {1{$random}};
    counts_421 = {1{$random}};
    counts_422 = {1{$random}};
    counts_423 = {1{$random}};
    counts_424 = {1{$random}};
    counts_425 = {1{$random}};
    counts_426 = {1{$random}};
    counts_427 = {1{$random}};
    counts_428 = {1{$random}};
    counts_429 = {1{$random}};
    counts_430 = {1{$random}};
    counts_431 = {1{$random}};
    counts_432 = {1{$random}};
    counts_433 = {1{$random}};
    counts_434 = {1{$random}};
    counts_435 = {1{$random}};
    counts_436 = {1{$random}};
    counts_437 = {1{$random}};
    counts_438 = {1{$random}};
    counts_439 = {1{$random}};
    counts_440 = {1{$random}};
    counts_441 = {1{$random}};
    counts_442 = {1{$random}};
    counts_443 = {1{$random}};
    counts_444 = {1{$random}};
    counts_445 = {1{$random}};
    counts_446 = {1{$random}};
    counts_447 = {1{$random}};
    counts_448 = {1{$random}};
    counts_449 = {1{$random}};
    counts_450 = {1{$random}};
    counts_451 = {1{$random}};
    counts_452 = {1{$random}};
    counts_453 = {1{$random}};
    counts_454 = {1{$random}};
    counts_455 = {1{$random}};
    counts_456 = {1{$random}};
    counts_457 = {1{$random}};
    counts_458 = {1{$random}};
    counts_459 = {1{$random}};
    counts_460 = {1{$random}};
    counts_461 = {1{$random}};
    counts_462 = {1{$random}};
    counts_463 = {1{$random}};
    counts_464 = {1{$random}};
    counts_465 = {1{$random}};
    counts_466 = {1{$random}};
    counts_467 = {1{$random}};
    counts_468 = {1{$random}};
    counts_469 = {1{$random}};
    counts_470 = {1{$random}};
    counts_471 = {1{$random}};
    counts_472 = {1{$random}};
    counts_473 = {1{$random}};
    counts_474 = {1{$random}};
    counts_475 = {1{$random}};
    counts_476 = {1{$random}};
    counts_477 = {1{$random}};
    counts_478 = {1{$random}};
    counts_479 = {1{$random}};
    counts_480 = {1{$random}};
    counts_481 = {1{$random}};
    counts_482 = {1{$random}};
    counts_483 = {1{$random}};
    counts_484 = {1{$random}};
    counts_485 = {1{$random}};
    counts_486 = {1{$random}};
    counts_487 = {1{$random}};
    counts_488 = {1{$random}};
    counts_489 = {1{$random}};
    counts_490 = {1{$random}};
    counts_491 = {1{$random}};
    counts_492 = {1{$random}};
    counts_493 = {1{$random}};
    counts_494 = {1{$random}};
    counts_495 = {1{$random}};
    counts_496 = {1{$random}};
    counts_497 = {1{$random}};
    counts_498 = {1{$random}};
    counts_499 = {1{$random}};
    counts_500 = {1{$random}};
    counts_501 = {1{$random}};
    counts_502 = {1{$random}};
    counts_503 = {1{$random}};
    counts_504 = {1{$random}};
    counts_505 = {1{$random}};
    counts_506 = {1{$random}};
    counts_507 = {1{$random}};
    counts_508 = {1{$random}};
    counts_509 = {1{$random}};
    counts_510 = {1{$random}};
    counts_511 = {1{$random}};
    counts_512 = {1{$random}};
    counts_513 = {1{$random}};
    counts_514 = {1{$random}};
    counts_515 = {1{$random}};
    counts_516 = {1{$random}};
    counts_517 = {1{$random}};
    counts_518 = {1{$random}};
    counts_519 = {1{$random}};
    counts_520 = {1{$random}};
    counts_521 = {1{$random}};
    counts_522 = {1{$random}};
    counts_523 = {1{$random}};
    counts_524 = {1{$random}};
    counts_525 = {1{$random}};
    counts_526 = {1{$random}};
    counts_527 = {1{$random}};
    counts_528 = {1{$random}};
    counts_529 = {1{$random}};
    counts_530 = {1{$random}};
    counts_531 = {1{$random}};
    counts_532 = {1{$random}};
    counts_533 = {1{$random}};
    counts_534 = {1{$random}};
    counts_535 = {1{$random}};
    counts_536 = {1{$random}};
    counts_537 = {1{$random}};
    counts_538 = {1{$random}};
    counts_539 = {1{$random}};
    counts_540 = {1{$random}};
    counts_541 = {1{$random}};
    counts_542 = {1{$random}};
    counts_543 = {1{$random}};
    counts_544 = {1{$random}};
    counts_545 = {1{$random}};
    counts_546 = {1{$random}};
    counts_547 = {1{$random}};
    counts_548 = {1{$random}};
    counts_549 = {1{$random}};
    counts_550 = {1{$random}};
    counts_551 = {1{$random}};
    counts_552 = {1{$random}};
    counts_553 = {1{$random}};
    counts_554 = {1{$random}};
    counts_555 = {1{$random}};
    counts_556 = {1{$random}};
    counts_557 = {1{$random}};
    counts_558 = {1{$random}};
    counts_559 = {1{$random}};
    counts_560 = {1{$random}};
    counts_561 = {1{$random}};
    counts_562 = {1{$random}};
    counts_563 = {1{$random}};
    counts_564 = {1{$random}};
    counts_565 = {1{$random}};
    counts_566 = {1{$random}};
    counts_567 = {1{$random}};
    counts_568 = {1{$random}};
    counts_569 = {1{$random}};
    counts_570 = {1{$random}};
    counts_571 = {1{$random}};
    counts_572 = {1{$random}};
    counts_573 = {1{$random}};
    counts_574 = {1{$random}};
    counts_575 = {1{$random}};
    counts_576 = {1{$random}};
    counts_577 = {1{$random}};
    counts_578 = {1{$random}};
    counts_579 = {1{$random}};
    counts_580 = {1{$random}};
    counts_581 = {1{$random}};
    counts_582 = {1{$random}};
    counts_583 = {1{$random}};
    counts_584 = {1{$random}};
    counts_585 = {1{$random}};
    counts_586 = {1{$random}};
    counts_587 = {1{$random}};
    counts_588 = {1{$random}};
    counts_589 = {1{$random}};
    counts_590 = {1{$random}};
    counts_591 = {1{$random}};
    counts_592 = {1{$random}};
    counts_593 = {1{$random}};
    counts_594 = {1{$random}};
    counts_595 = {1{$random}};
    counts_596 = {1{$random}};
    counts_597 = {1{$random}};
    counts_598 = {1{$random}};
    counts_599 = {1{$random}};
    counts_600 = {1{$random}};
    counts_601 = {1{$random}};
    counts_602 = {1{$random}};
    counts_603 = {1{$random}};
    counts_604 = {1{$random}};
    counts_605 = {1{$random}};
    counts_606 = {1{$random}};
    counts_607 = {1{$random}};
    counts_608 = {1{$random}};
    counts_609 = {1{$random}};
    counts_610 = {1{$random}};
    counts_611 = {1{$random}};
    counts_612 = {1{$random}};
    counts_613 = {1{$random}};
    counts_614 = {1{$random}};
    counts_615 = {1{$random}};
    counts_616 = {1{$random}};
    counts_617 = {1{$random}};
    counts_618 = {1{$random}};
    counts_619 = {1{$random}};
    counts_620 = {1{$random}};
    counts_621 = {1{$random}};
    counts_622 = {1{$random}};
    counts_623 = {1{$random}};
    counts_624 = {1{$random}};
    counts_625 = {1{$random}};
    counts_626 = {1{$random}};
    counts_627 = {1{$random}};
    counts_628 = {1{$random}};
    counts_629 = {1{$random}};
    counts_630 = {1{$random}};
    counts_631 = {1{$random}};
    counts_632 = {1{$random}};
    counts_633 = {1{$random}};
    counts_634 = {1{$random}};
    counts_635 = {1{$random}};
    counts_636 = {1{$random}};
    counts_637 = {1{$random}};
    counts_638 = {1{$random}};
    counts_639 = {1{$random}};
    counts_640 = {1{$random}};
    counts_641 = {1{$random}};
    counts_642 = {1{$random}};
    counts_643 = {1{$random}};
    counts_644 = {1{$random}};
    counts_645 = {1{$random}};
    counts_646 = {1{$random}};
    counts_647 = {1{$random}};
    counts_648 = {1{$random}};
    counts_649 = {1{$random}};
    counts_650 = {1{$random}};
    counts_651 = {1{$random}};
    counts_652 = {1{$random}};
    counts_653 = {1{$random}};
    counts_654 = {1{$random}};
    counts_655 = {1{$random}};
    counts_656 = {1{$random}};
    counts_657 = {1{$random}};
    counts_658 = {1{$random}};
    counts_659 = {1{$random}};
    counts_660 = {1{$random}};
    counts_661 = {1{$random}};
    counts_662 = {1{$random}};
    counts_663 = {1{$random}};
    counts_664 = {1{$random}};
    counts_665 = {1{$random}};
    counts_666 = {1{$random}};
    counts_667 = {1{$random}};
    counts_668 = {1{$random}};
    counts_669 = {1{$random}};
    counts_670 = {1{$random}};
    counts_671 = {1{$random}};
    counts_672 = {1{$random}};
    counts_673 = {1{$random}};
    counts_674 = {1{$random}};
    counts_675 = {1{$random}};
    counts_676 = {1{$random}};
    counts_677 = {1{$random}};
    counts_678 = {1{$random}};
    counts_679 = {1{$random}};
    counts_680 = {1{$random}};
    counts_681 = {1{$random}};
    counts_682 = {1{$random}};
    counts_683 = {1{$random}};
    counts_684 = {1{$random}};
    counts_685 = {1{$random}};
    counts_686 = {1{$random}};
    counts_687 = {1{$random}};
    counts_688 = {1{$random}};
    counts_689 = {1{$random}};
    counts_690 = {1{$random}};
    counts_691 = {1{$random}};
    counts_692 = {1{$random}};
    counts_693 = {1{$random}};
    counts_694 = {1{$random}};
    counts_695 = {1{$random}};
    counts_696 = {1{$random}};
    counts_697 = {1{$random}};
    counts_698 = {1{$random}};
    counts_699 = {1{$random}};
    counts_700 = {1{$random}};
    counts_701 = {1{$random}};
    counts_702 = {1{$random}};
    counts_703 = {1{$random}};
    counts_704 = {1{$random}};
    counts_705 = {1{$random}};
    counts_706 = {1{$random}};
    counts_707 = {1{$random}};
    counts_708 = {1{$random}};
    counts_709 = {1{$random}};
    counts_710 = {1{$random}};
    counts_711 = {1{$random}};
    counts_712 = {1{$random}};
    counts_713 = {1{$random}};
    counts_714 = {1{$random}};
    counts_715 = {1{$random}};
    counts_716 = {1{$random}};
    counts_717 = {1{$random}};
    counts_718 = {1{$random}};
    counts_719 = {1{$random}};
    counts_720 = {1{$random}};
    counts_721 = {1{$random}};
    counts_722 = {1{$random}};
    counts_723 = {1{$random}};
    counts_724 = {1{$random}};
    counts_725 = {1{$random}};
    counts_726 = {1{$random}};
    counts_727 = {1{$random}};
    counts_728 = {1{$random}};
    counts_729 = {1{$random}};
    counts_730 = {1{$random}};
    counts_731 = {1{$random}};
    counts_732 = {1{$random}};
    counts_733 = {1{$random}};
    counts_734 = {1{$random}};
    counts_735 = {1{$random}};
    counts_736 = {1{$random}};
    counts_737 = {1{$random}};
    counts_738 = {1{$random}};
    counts_739 = {1{$random}};
    counts_740 = {1{$random}};
    counts_741 = {1{$random}};
    counts_742 = {1{$random}};
    counts_743 = {1{$random}};
    counts_744 = {1{$random}};
    counts_745 = {1{$random}};
    counts_746 = {1{$random}};
    counts_747 = {1{$random}};
    counts_748 = {1{$random}};
    counts_749 = {1{$random}};
    counts_750 = {1{$random}};
    counts_751 = {1{$random}};
    counts_752 = {1{$random}};
    counts_753 = {1{$random}};
    counts_754 = {1{$random}};
    counts_755 = {1{$random}};
    counts_756 = {1{$random}};
    counts_757 = {1{$random}};
    counts_758 = {1{$random}};
    counts_759 = {1{$random}};
    counts_760 = {1{$random}};
    counts_761 = {1{$random}};
    counts_762 = {1{$random}};
    counts_763 = {1{$random}};
    counts_764 = {1{$random}};
    counts_765 = {1{$random}};
    counts_766 = {1{$random}};
    counts_767 = {1{$random}};
    counts_768 = {1{$random}};
    counts_769 = {1{$random}};
    counts_770 = {1{$random}};
    counts_771 = {1{$random}};
    counts_772 = {1{$random}};
    counts_773 = {1{$random}};
    counts_774 = {1{$random}};
    counts_775 = {1{$random}};
    counts_776 = {1{$random}};
    counts_777 = {1{$random}};
    counts_778 = {1{$random}};
    counts_779 = {1{$random}};
    counts_780 = {1{$random}};
    counts_781 = {1{$random}};
    counts_782 = {1{$random}};
    counts_783 = {1{$random}};
    counts_784 = {1{$random}};
    counts_785 = {1{$random}};
    counts_786 = {1{$random}};
    counts_787 = {1{$random}};
    counts_788 = {1{$random}};
    counts_789 = {1{$random}};
    counts_790 = {1{$random}};
    counts_791 = {1{$random}};
    counts_792 = {1{$random}};
    counts_793 = {1{$random}};
    counts_794 = {1{$random}};
    counts_795 = {1{$random}};
    counts_796 = {1{$random}};
    counts_797 = {1{$random}};
    counts_798 = {1{$random}};
    counts_799 = {1{$random}};
    counts_800 = {1{$random}};
    counts_801 = {1{$random}};
    counts_802 = {1{$random}};
    counts_803 = {1{$random}};
    counts_804 = {1{$random}};
    counts_805 = {1{$random}};
    counts_806 = {1{$random}};
    counts_807 = {1{$random}};
    counts_808 = {1{$random}};
    counts_809 = {1{$random}};
    counts_810 = {1{$random}};
    counts_811 = {1{$random}};
    counts_812 = {1{$random}};
    counts_813 = {1{$random}};
    counts_814 = {1{$random}};
    counts_815 = {1{$random}};
    counts_816 = {1{$random}};
    counts_817 = {1{$random}};
    counts_818 = {1{$random}};
    counts_819 = {1{$random}};
    counts_820 = {1{$random}};
    counts_821 = {1{$random}};
    counts_822 = {1{$random}};
    counts_823 = {1{$random}};
    counts_824 = {1{$random}};
    counts_825 = {1{$random}};
    counts_826 = {1{$random}};
    counts_827 = {1{$random}};
    counts_828 = {1{$random}};
    counts_829 = {1{$random}};
    counts_830 = {1{$random}};
    counts_831 = {1{$random}};
    counts_832 = {1{$random}};
    counts_833 = {1{$random}};
    counts_834 = {1{$random}};
    counts_835 = {1{$random}};
    counts_836 = {1{$random}};
    counts_837 = {1{$random}};
    counts_838 = {1{$random}};
    counts_839 = {1{$random}};
    counts_840 = {1{$random}};
    counts_841 = {1{$random}};
    counts_842 = {1{$random}};
    counts_843 = {1{$random}};
    counts_844 = {1{$random}};
    counts_845 = {1{$random}};
    counts_846 = {1{$random}};
    counts_847 = {1{$random}};
    counts_848 = {1{$random}};
    counts_849 = {1{$random}};
    counts_850 = {1{$random}};
    counts_851 = {1{$random}};
    counts_852 = {1{$random}};
    counts_853 = {1{$random}};
    counts_854 = {1{$random}};
    counts_855 = {1{$random}};
    counts_856 = {1{$random}};
    counts_857 = {1{$random}};
    counts_858 = {1{$random}};
    counts_859 = {1{$random}};
    counts_860 = {1{$random}};
    counts_861 = {1{$random}};
    counts_862 = {1{$random}};
    counts_863 = {1{$random}};
    counts_864 = {1{$random}};
    counts_865 = {1{$random}};
    counts_866 = {1{$random}};
    counts_867 = {1{$random}};
    counts_868 = {1{$random}};
    counts_869 = {1{$random}};
    counts_870 = {1{$random}};
    counts_871 = {1{$random}};
    counts_872 = {1{$random}};
    counts_873 = {1{$random}};
    counts_874 = {1{$random}};
    counts_875 = {1{$random}};
    counts_876 = {1{$random}};
    counts_877 = {1{$random}};
    counts_878 = {1{$random}};
    counts_879 = {1{$random}};
    counts_880 = {1{$random}};
    counts_881 = {1{$random}};
    counts_882 = {1{$random}};
    counts_883 = {1{$random}};
    counts_884 = {1{$random}};
    counts_885 = {1{$random}};
    counts_886 = {1{$random}};
    counts_887 = {1{$random}};
    counts_888 = {1{$random}};
    counts_889 = {1{$random}};
    counts_890 = {1{$random}};
    counts_891 = {1{$random}};
    counts_892 = {1{$random}};
    counts_893 = {1{$random}};
    counts_894 = {1{$random}};
    counts_895 = {1{$random}};
    counts_896 = {1{$random}};
    counts_897 = {1{$random}};
    counts_898 = {1{$random}};
    counts_899 = {1{$random}};
    counts_900 = {1{$random}};
    counts_901 = {1{$random}};
    counts_902 = {1{$random}};
    counts_903 = {1{$random}};
    counts_904 = {1{$random}};
    counts_905 = {1{$random}};
    counts_906 = {1{$random}};
    counts_907 = {1{$random}};
    counts_908 = {1{$random}};
    counts_909 = {1{$random}};
    counts_910 = {1{$random}};
    counts_911 = {1{$random}};
    counts_912 = {1{$random}};
    counts_913 = {1{$random}};
    counts_914 = {1{$random}};
    counts_915 = {1{$random}};
    counts_916 = {1{$random}};
    counts_917 = {1{$random}};
    counts_918 = {1{$random}};
    counts_919 = {1{$random}};
    counts_920 = {1{$random}};
    counts_921 = {1{$random}};
    counts_922 = {1{$random}};
    counts_923 = {1{$random}};
    counts_924 = {1{$random}};
    counts_925 = {1{$random}};
    counts_926 = {1{$random}};
    counts_927 = {1{$random}};
    counts_928 = {1{$random}};
    counts_929 = {1{$random}};
    counts_930 = {1{$random}};
    counts_931 = {1{$random}};
    counts_932 = {1{$random}};
    counts_933 = {1{$random}};
    counts_934 = {1{$random}};
    counts_935 = {1{$random}};
    counts_936 = {1{$random}};
    counts_937 = {1{$random}};
    counts_938 = {1{$random}};
    counts_939 = {1{$random}};
    counts_940 = {1{$random}};
    counts_941 = {1{$random}};
    counts_942 = {1{$random}};
    counts_943 = {1{$random}};
    counts_944 = {1{$random}};
    counts_945 = {1{$random}};
    counts_946 = {1{$random}};
    counts_947 = {1{$random}};
    counts_948 = {1{$random}};
    counts_949 = {1{$random}};
    counts_950 = {1{$random}};
    counts_951 = {1{$random}};
    counts_952 = {1{$random}};
    counts_953 = {1{$random}};
    counts_954 = {1{$random}};
    counts_955 = {1{$random}};
    counts_956 = {1{$random}};
    counts_957 = {1{$random}};
    counts_958 = {1{$random}};
    counts_959 = {1{$random}};
    counts_960 = {1{$random}};
    counts_961 = {1{$random}};
    counts_962 = {1{$random}};
    counts_963 = {1{$random}};
    counts_964 = {1{$random}};
    counts_965 = {1{$random}};
    counts_966 = {1{$random}};
    counts_967 = {1{$random}};
    counts_968 = {1{$random}};
    counts_969 = {1{$random}};
    counts_970 = {1{$random}};
    counts_971 = {1{$random}};
    counts_972 = {1{$random}};
    counts_973 = {1{$random}};
    counts_974 = {1{$random}};
    counts_975 = {1{$random}};
    counts_976 = {1{$random}};
    counts_977 = {1{$random}};
    counts_978 = {1{$random}};
    counts_979 = {1{$random}};
    counts_980 = {1{$random}};
    counts_981 = {1{$random}};
    counts_982 = {1{$random}};
    counts_983 = {1{$random}};
    counts_984 = {1{$random}};
    counts_985 = {1{$random}};
    counts_986 = {1{$random}};
    counts_987 = {1{$random}};
    counts_988 = {1{$random}};
    counts_989 = {1{$random}};
    counts_990 = {1{$random}};
    counts_991 = {1{$random}};
    counts_992 = {1{$random}};
    counts_993 = {1{$random}};
    counts_994 = {1{$random}};
    counts_995 = {1{$random}};
    counts_996 = {1{$random}};
    counts_997 = {1{$random}};
    counts_998 = {1{$random}};
    counts_999 = {1{$random}};
    counts_1000 = {1{$random}};
    counts_1001 = {1{$random}};
    counts_1002 = {1{$random}};
    counts_1003 = {1{$random}};
    counts_1004 = {1{$random}};
    counts_1005 = {1{$random}};
    counts_1006 = {1{$random}};
    counts_1007 = {1{$random}};
    counts_1008 = {1{$random}};
    counts_1009 = {1{$random}};
    counts_1010 = {1{$random}};
    counts_1011 = {1{$random}};
    counts_1012 = {1{$random}};
    counts_1013 = {1{$random}};
    counts_1014 = {1{$random}};
    counts_1015 = {1{$random}};
    counts_1016 = {1{$random}};
    counts_1017 = {1{$random}};
    counts_1018 = {1{$random}};
    counts_1019 = {1{$random}};
    counts_1020 = {1{$random}};
    counts_1021 = {1{$random}};
    counts_1022 = {1{$random}};
    counts_1023 = {1{$random}};
    counts_1 = {1{$random}};
    hashCount1 = {1{$random}};
    delayCount = {1{$random}};
    delayedIndex = {1{$random}};
    R10323 = {1{$random}};
    index = {1{$random}};
    curInfo_tag = {1{$random}};
  end
`endif

  assign io_hashOut_bits_found = hashFound;
  assign T0 = T10339 ? T10337 : T1;
  assign T1 = T10320 ? 1'h1 : T2;
  assign T2 = T10319 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : hashFound;
  assign T4 = 3'h0 == state;
  assign T10343 = reset ? 3'h0 : T5;
  assign T5 = T10317 ? 3'h0 : T6;
  assign T6 = T10339 ? 3'h7 : T7;
  assign T7 = T10316 ? 3'h6 : T8;
  assign T8 = T10320 ? 3'h7 : T9;
  assign T9 = T10313 ? 3'h7 : T10;
  assign T10 = T10310 ? 3'h5 : T11;
  assign T11 = T10306 ? 3'h1 : T12;
  assign T12 = T10298 ? 3'h4 : T13;
  assign T13 = T10295 ? 3'h7 : T14;
  assign T14 = T10291 ? 3'h5 : T15;
  assign T15 = T30 ? 3'h1 : T16;
  assign T16 = T22 ? 3'h3 : T17;
  assign T17 = T10319 ? 3'h7 : T18;
  assign T18 = T21 ? 3'h2 : T19;
  assign T19 = T20 ? 3'h1 : state;
  assign T20 = T4 & io_hashIn_valid;
  assign T21 = 3'h1 == state;
  assign T22 = T29 & T23;
  assign T23 = T26 & T24;
  assign T24 = io_lenData == curInfo_len;
  assign T25 = T20 ? io_hashIn_bits_len : curInfo_len;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_findAvailable & T28;
  assign T28 = io_lenData == 8'h0;
  assign T29 = 3'h2 == state;
  assign T30 = T29 & T31;
  assign T31 = T10289 & checkFirst;
  assign T32 = T10287 ? 1'h0 : T33;
  assign T33 = T37 ? 1'h1 : T34;
  assign T34 = T10306 ? 1'h0 : T35;
  assign T35 = T30 ? 1'h0 : T36;
  assign T36 = T4 ? 1'h1 : checkFirst;
  assign T37 = T10316 & T38;
  assign T38 = hashCount1 < hashCount2;
  assign T10344 = reset ? 4'h0 : T39;
  assign T39 = T21 ? T40 : hashCount2;
  assign T40 = T8238 ? T7216 : T41;
  assign T41 = T7215 ? T6705 : T42;
  assign T42 = T6704 ? T6450 : T43;
  assign T43 = T6449 ? T6323 : T44;
  assign T44 = T6322 ? T6260 : T45;
  assign T45 = T6259 ? T6229 : T46;
  assign T46 = T6228 ? T6214 : T47;
  assign T47 = T6213 ? T6207 : T48;
  assign T48 = T6206 ? T6204 : T49;
  assign T49 = T6202 ? counts_1 : counts_0;
  assign T10345 = reset ? 4'h0 : T50;
  assign T50 = T6196 ? T52 : T51;
  assign T51 = io_resetCounts ? 4'h0 : counts_0;
  assign T52 = T6195 ^ T53;
  assign T53 = 4'h0 - T10346;
  assign T10346 = {3'h0, T54};
  assign T54 = T55[3'h4:3'h4];
  assign T55 = T56 + 5'h1;
  assign T56 = {1'h0, T57};
  assign T57 = T6194 ? T3124 : T58;
  assign T58 = T3123 ? T1589 : T59;
  assign T59 = T1588 ? T822 : T60;
  assign T60 = T821 ? T439 : T61;
  assign T61 = T438 ? T248 : T62;
  assign T62 = T247 ? T153 : T63;
  assign T63 = T152 ? T106 : T64;
  assign T64 = T105 ? T83 : T65;
  assign T65 = T82 ? T71 : T66;
  assign T66 = T67 ? counts_1 : counts_0;
  assign T67 = T68[1'h0:1'h0];
  assign T68 = curHash;
  assign curHash = checkFirst ? curInfo_hash1 : curInfo_hash2;
  assign T69 = T20 ? io_hashIn_bits_hash2 : curInfo_hash2;
  assign T70 = T20 ? io_hashIn_bits_hash1 : curInfo_hash1;
  assign T71 = T81 ? counts_3 : counts_2;
  assign T10347 = reset ? 4'h0 : T72;
  assign T72 = T74 ? T52 : T73;
  assign T73 = io_resetCounts ? 4'h0 : counts_2;
  assign T74 = T10320 & T75;
  assign T75 = T76[2'h2:2'h2];
  assign T76 = 1'h1 << T68;
  assign T10348 = reset ? 4'h0 : T77;
  assign T77 = T79 ? T52 : T78;
  assign T78 = io_resetCounts ? 4'h0 : counts_3;
  assign T79 = T10320 & T80;
  assign T80 = T76[2'h3:2'h3];
  assign T81 = T68[1'h0:1'h0];
  assign T82 = T68[1'h1:1'h1];
  assign T83 = T104 ? T94 : T84;
  assign T84 = T93 ? counts_5 : counts_4;
  assign T10349 = reset ? 4'h0 : T85;
  assign T85 = T87 ? T52 : T86;
  assign T86 = io_resetCounts ? 4'h0 : counts_4;
  assign T87 = T10320 & T88;
  assign T88 = T76[3'h4:3'h4];
  assign T10350 = reset ? 4'h0 : T89;
  assign T89 = T91 ? T52 : T90;
  assign T90 = io_resetCounts ? 4'h0 : counts_5;
  assign T91 = T10320 & T92;
  assign T92 = T76[3'h5:3'h5];
  assign T93 = T68[1'h0:1'h0];
  assign T94 = T103 ? counts_7 : counts_6;
  assign T10351 = reset ? 4'h0 : T95;
  assign T95 = T97 ? T52 : T96;
  assign T96 = io_resetCounts ? 4'h0 : counts_6;
  assign T97 = T10320 & T98;
  assign T98 = T76[3'h6:3'h6];
  assign T10352 = reset ? 4'h0 : T99;
  assign T99 = T101 ? T52 : T100;
  assign T100 = io_resetCounts ? 4'h0 : counts_7;
  assign T101 = T10320 & T102;
  assign T102 = T76[3'h7:3'h7];
  assign T103 = T68[1'h0:1'h0];
  assign T104 = T68[1'h1:1'h1];
  assign T105 = T68[2'h2:2'h2];
  assign T106 = T151 ? T129 : T107;
  assign T107 = T128 ? T118 : T108;
  assign T108 = T117 ? counts_9 : counts_8;
  assign T10353 = reset ? 4'h0 : T109;
  assign T109 = T111 ? T52 : T110;
  assign T110 = io_resetCounts ? 4'h0 : counts_8;
  assign T111 = T10320 & T112;
  assign T112 = T76[4'h8:4'h8];
  assign T10354 = reset ? 4'h0 : T113;
  assign T113 = T115 ? T52 : T114;
  assign T114 = io_resetCounts ? 4'h0 : counts_9;
  assign T115 = T10320 & T116;
  assign T116 = T76[4'h9:4'h9];
  assign T117 = T68[1'h0:1'h0];
  assign T118 = T127 ? counts_11 : counts_10;
  assign T10355 = reset ? 4'h0 : T119;
  assign T119 = T121 ? T52 : T120;
  assign T120 = io_resetCounts ? 4'h0 : counts_10;
  assign T121 = T10320 & T122;
  assign T122 = T76[4'ha:4'ha];
  assign T10356 = reset ? 4'h0 : T123;
  assign T123 = T125 ? T52 : T124;
  assign T124 = io_resetCounts ? 4'h0 : counts_11;
  assign T125 = T10320 & T126;
  assign T126 = T76[4'hb:4'hb];
  assign T127 = T68[1'h0:1'h0];
  assign T128 = T68[1'h1:1'h1];
  assign T129 = T150 ? T140 : T130;
  assign T130 = T139 ? counts_13 : counts_12;
  assign T10357 = reset ? 4'h0 : T131;
  assign T131 = T133 ? T52 : T132;
  assign T132 = io_resetCounts ? 4'h0 : counts_12;
  assign T133 = T10320 & T134;
  assign T134 = T76[4'hc:4'hc];
  assign T10358 = reset ? 4'h0 : T135;
  assign T135 = T137 ? T52 : T136;
  assign T136 = io_resetCounts ? 4'h0 : counts_13;
  assign T137 = T10320 & T138;
  assign T138 = T76[4'hd:4'hd];
  assign T139 = T68[1'h0:1'h0];
  assign T140 = T149 ? counts_15 : counts_14;
  assign T10359 = reset ? 4'h0 : T141;
  assign T141 = T143 ? T52 : T142;
  assign T142 = io_resetCounts ? 4'h0 : counts_14;
  assign T143 = T10320 & T144;
  assign T144 = T76[4'he:4'he];
  assign T10360 = reset ? 4'h0 : T145;
  assign T145 = T147 ? T52 : T146;
  assign T146 = io_resetCounts ? 4'h0 : counts_15;
  assign T147 = T10320 & T148;
  assign T148 = T76[4'hf:4'hf];
  assign T149 = T68[1'h0:1'h0];
  assign T150 = T68[1'h1:1'h1];
  assign T151 = T68[2'h2:2'h2];
  assign T152 = T68[2'h3:2'h3];
  assign T153 = T246 ? T200 : T154;
  assign T154 = T199 ? T177 : T155;
  assign T155 = T176 ? T166 : T156;
  assign T156 = T165 ? counts_17 : counts_16;
  assign T10361 = reset ? 4'h0 : T157;
  assign T157 = T159 ? T52 : T158;
  assign T158 = io_resetCounts ? 4'h0 : counts_16;
  assign T159 = T10320 & T160;
  assign T160 = T76[5'h10:5'h10];
  assign T10362 = reset ? 4'h0 : T161;
  assign T161 = T163 ? T52 : T162;
  assign T162 = io_resetCounts ? 4'h0 : counts_17;
  assign T163 = T10320 & T164;
  assign T164 = T76[5'h11:5'h11];
  assign T165 = T68[1'h0:1'h0];
  assign T166 = T175 ? counts_19 : counts_18;
  assign T10363 = reset ? 4'h0 : T167;
  assign T167 = T169 ? T52 : T168;
  assign T168 = io_resetCounts ? 4'h0 : counts_18;
  assign T169 = T10320 & T170;
  assign T170 = T76[5'h12:5'h12];
  assign T10364 = reset ? 4'h0 : T171;
  assign T171 = T173 ? T52 : T172;
  assign T172 = io_resetCounts ? 4'h0 : counts_19;
  assign T173 = T10320 & T174;
  assign T174 = T76[5'h13:5'h13];
  assign T175 = T68[1'h0:1'h0];
  assign T176 = T68[1'h1:1'h1];
  assign T177 = T198 ? T188 : T178;
  assign T178 = T187 ? counts_21 : counts_20;
  assign T10365 = reset ? 4'h0 : T179;
  assign T179 = T181 ? T52 : T180;
  assign T180 = io_resetCounts ? 4'h0 : counts_20;
  assign T181 = T10320 & T182;
  assign T182 = T76[5'h14:5'h14];
  assign T10366 = reset ? 4'h0 : T183;
  assign T183 = T185 ? T52 : T184;
  assign T184 = io_resetCounts ? 4'h0 : counts_21;
  assign T185 = T10320 & T186;
  assign T186 = T76[5'h15:5'h15];
  assign T187 = T68[1'h0:1'h0];
  assign T188 = T197 ? counts_23 : counts_22;
  assign T10367 = reset ? 4'h0 : T189;
  assign T189 = T191 ? T52 : T190;
  assign T190 = io_resetCounts ? 4'h0 : counts_22;
  assign T191 = T10320 & T192;
  assign T192 = T76[5'h16:5'h16];
  assign T10368 = reset ? 4'h0 : T193;
  assign T193 = T195 ? T52 : T194;
  assign T194 = io_resetCounts ? 4'h0 : counts_23;
  assign T195 = T10320 & T196;
  assign T196 = T76[5'h17:5'h17];
  assign T197 = T68[1'h0:1'h0];
  assign T198 = T68[1'h1:1'h1];
  assign T199 = T68[2'h2:2'h2];
  assign T200 = T245 ? T223 : T201;
  assign T201 = T222 ? T212 : T202;
  assign T202 = T211 ? counts_25 : counts_24;
  assign T10369 = reset ? 4'h0 : T203;
  assign T203 = T205 ? T52 : T204;
  assign T204 = io_resetCounts ? 4'h0 : counts_24;
  assign T205 = T10320 & T206;
  assign T206 = T76[5'h18:5'h18];
  assign T10370 = reset ? 4'h0 : T207;
  assign T207 = T209 ? T52 : T208;
  assign T208 = io_resetCounts ? 4'h0 : counts_25;
  assign T209 = T10320 & T210;
  assign T210 = T76[5'h19:5'h19];
  assign T211 = T68[1'h0:1'h0];
  assign T212 = T221 ? counts_27 : counts_26;
  assign T10371 = reset ? 4'h0 : T213;
  assign T213 = T215 ? T52 : T214;
  assign T214 = io_resetCounts ? 4'h0 : counts_26;
  assign T215 = T10320 & T216;
  assign T216 = T76[5'h1a:5'h1a];
  assign T10372 = reset ? 4'h0 : T217;
  assign T217 = T219 ? T52 : T218;
  assign T218 = io_resetCounts ? 4'h0 : counts_27;
  assign T219 = T10320 & T220;
  assign T220 = T76[5'h1b:5'h1b];
  assign T221 = T68[1'h0:1'h0];
  assign T222 = T68[1'h1:1'h1];
  assign T223 = T244 ? T234 : T224;
  assign T224 = T233 ? counts_29 : counts_28;
  assign T10373 = reset ? 4'h0 : T225;
  assign T225 = T227 ? T52 : T226;
  assign T226 = io_resetCounts ? 4'h0 : counts_28;
  assign T227 = T10320 & T228;
  assign T228 = T76[5'h1c:5'h1c];
  assign T10374 = reset ? 4'h0 : T229;
  assign T229 = T231 ? T52 : T230;
  assign T230 = io_resetCounts ? 4'h0 : counts_29;
  assign T231 = T10320 & T232;
  assign T232 = T76[5'h1d:5'h1d];
  assign T233 = T68[1'h0:1'h0];
  assign T234 = T243 ? counts_31 : counts_30;
  assign T10375 = reset ? 4'h0 : T235;
  assign T235 = T237 ? T52 : T236;
  assign T236 = io_resetCounts ? 4'h0 : counts_30;
  assign T237 = T10320 & T238;
  assign T238 = T76[5'h1e:5'h1e];
  assign T10376 = reset ? 4'h0 : T239;
  assign T239 = T241 ? T52 : T240;
  assign T240 = io_resetCounts ? 4'h0 : counts_31;
  assign T241 = T10320 & T242;
  assign T242 = T76[5'h1f:5'h1f];
  assign T243 = T68[1'h0:1'h0];
  assign T244 = T68[1'h1:1'h1];
  assign T245 = T68[2'h2:2'h2];
  assign T246 = T68[2'h3:2'h3];
  assign T247 = T68[3'h4:3'h4];
  assign T248 = T437 ? T343 : T249;
  assign T249 = T342 ? T296 : T250;
  assign T250 = T295 ? T273 : T251;
  assign T251 = T272 ? T262 : T252;
  assign T252 = T261 ? counts_33 : counts_32;
  assign T10377 = reset ? 4'h0 : T253;
  assign T253 = T255 ? T52 : T254;
  assign T254 = io_resetCounts ? 4'h0 : counts_32;
  assign T255 = T10320 & T256;
  assign T256 = T76[6'h20:6'h20];
  assign T10378 = reset ? 4'h0 : T257;
  assign T257 = T259 ? T52 : T258;
  assign T258 = io_resetCounts ? 4'h0 : counts_33;
  assign T259 = T10320 & T260;
  assign T260 = T76[6'h21:6'h21];
  assign T261 = T68[1'h0:1'h0];
  assign T262 = T271 ? counts_35 : counts_34;
  assign T10379 = reset ? 4'h0 : T263;
  assign T263 = T265 ? T52 : T264;
  assign T264 = io_resetCounts ? 4'h0 : counts_34;
  assign T265 = T10320 & T266;
  assign T266 = T76[6'h22:6'h22];
  assign T10380 = reset ? 4'h0 : T267;
  assign T267 = T269 ? T52 : T268;
  assign T268 = io_resetCounts ? 4'h0 : counts_35;
  assign T269 = T10320 & T270;
  assign T270 = T76[6'h23:6'h23];
  assign T271 = T68[1'h0:1'h0];
  assign T272 = T68[1'h1:1'h1];
  assign T273 = T294 ? T284 : T274;
  assign T274 = T283 ? counts_37 : counts_36;
  assign T10381 = reset ? 4'h0 : T275;
  assign T275 = T277 ? T52 : T276;
  assign T276 = io_resetCounts ? 4'h0 : counts_36;
  assign T277 = T10320 & T278;
  assign T278 = T76[6'h24:6'h24];
  assign T10382 = reset ? 4'h0 : T279;
  assign T279 = T281 ? T52 : T280;
  assign T280 = io_resetCounts ? 4'h0 : counts_37;
  assign T281 = T10320 & T282;
  assign T282 = T76[6'h25:6'h25];
  assign T283 = T68[1'h0:1'h0];
  assign T284 = T293 ? counts_39 : counts_38;
  assign T10383 = reset ? 4'h0 : T285;
  assign T285 = T287 ? T52 : T286;
  assign T286 = io_resetCounts ? 4'h0 : counts_38;
  assign T287 = T10320 & T288;
  assign T288 = T76[6'h26:6'h26];
  assign T10384 = reset ? 4'h0 : T289;
  assign T289 = T291 ? T52 : T290;
  assign T290 = io_resetCounts ? 4'h0 : counts_39;
  assign T291 = T10320 & T292;
  assign T292 = T76[6'h27:6'h27];
  assign T293 = T68[1'h0:1'h0];
  assign T294 = T68[1'h1:1'h1];
  assign T295 = T68[2'h2:2'h2];
  assign T296 = T341 ? T319 : T297;
  assign T297 = T318 ? T308 : T298;
  assign T298 = T307 ? counts_41 : counts_40;
  assign T10385 = reset ? 4'h0 : T299;
  assign T299 = T301 ? T52 : T300;
  assign T300 = io_resetCounts ? 4'h0 : counts_40;
  assign T301 = T10320 & T302;
  assign T302 = T76[6'h28:6'h28];
  assign T10386 = reset ? 4'h0 : T303;
  assign T303 = T305 ? T52 : T304;
  assign T304 = io_resetCounts ? 4'h0 : counts_41;
  assign T305 = T10320 & T306;
  assign T306 = T76[6'h29:6'h29];
  assign T307 = T68[1'h0:1'h0];
  assign T308 = T317 ? counts_43 : counts_42;
  assign T10387 = reset ? 4'h0 : T309;
  assign T309 = T311 ? T52 : T310;
  assign T310 = io_resetCounts ? 4'h0 : counts_42;
  assign T311 = T10320 & T312;
  assign T312 = T76[6'h2a:6'h2a];
  assign T10388 = reset ? 4'h0 : T313;
  assign T313 = T315 ? T52 : T314;
  assign T314 = io_resetCounts ? 4'h0 : counts_43;
  assign T315 = T10320 & T316;
  assign T316 = T76[6'h2b:6'h2b];
  assign T317 = T68[1'h0:1'h0];
  assign T318 = T68[1'h1:1'h1];
  assign T319 = T340 ? T330 : T320;
  assign T320 = T329 ? counts_45 : counts_44;
  assign T10389 = reset ? 4'h0 : T321;
  assign T321 = T323 ? T52 : T322;
  assign T322 = io_resetCounts ? 4'h0 : counts_44;
  assign T323 = T10320 & T324;
  assign T324 = T76[6'h2c:6'h2c];
  assign T10390 = reset ? 4'h0 : T325;
  assign T325 = T327 ? T52 : T326;
  assign T326 = io_resetCounts ? 4'h0 : counts_45;
  assign T327 = T10320 & T328;
  assign T328 = T76[6'h2d:6'h2d];
  assign T329 = T68[1'h0:1'h0];
  assign T330 = T339 ? counts_47 : counts_46;
  assign T10391 = reset ? 4'h0 : T331;
  assign T331 = T333 ? T52 : T332;
  assign T332 = io_resetCounts ? 4'h0 : counts_46;
  assign T333 = T10320 & T334;
  assign T334 = T76[6'h2e:6'h2e];
  assign T10392 = reset ? 4'h0 : T335;
  assign T335 = T337 ? T52 : T336;
  assign T336 = io_resetCounts ? 4'h0 : counts_47;
  assign T337 = T10320 & T338;
  assign T338 = T76[6'h2f:6'h2f];
  assign T339 = T68[1'h0:1'h0];
  assign T340 = T68[1'h1:1'h1];
  assign T341 = T68[2'h2:2'h2];
  assign T342 = T68[2'h3:2'h3];
  assign T343 = T436 ? T390 : T344;
  assign T344 = T389 ? T367 : T345;
  assign T345 = T366 ? T356 : T346;
  assign T346 = T355 ? counts_49 : counts_48;
  assign T10393 = reset ? 4'h0 : T347;
  assign T347 = T349 ? T52 : T348;
  assign T348 = io_resetCounts ? 4'h0 : counts_48;
  assign T349 = T10320 & T350;
  assign T350 = T76[6'h30:6'h30];
  assign T10394 = reset ? 4'h0 : T351;
  assign T351 = T353 ? T52 : T352;
  assign T352 = io_resetCounts ? 4'h0 : counts_49;
  assign T353 = T10320 & T354;
  assign T354 = T76[6'h31:6'h31];
  assign T355 = T68[1'h0:1'h0];
  assign T356 = T365 ? counts_51 : counts_50;
  assign T10395 = reset ? 4'h0 : T357;
  assign T357 = T359 ? T52 : T358;
  assign T358 = io_resetCounts ? 4'h0 : counts_50;
  assign T359 = T10320 & T360;
  assign T360 = T76[6'h32:6'h32];
  assign T10396 = reset ? 4'h0 : T361;
  assign T361 = T363 ? T52 : T362;
  assign T362 = io_resetCounts ? 4'h0 : counts_51;
  assign T363 = T10320 & T364;
  assign T364 = T76[6'h33:6'h33];
  assign T365 = T68[1'h0:1'h0];
  assign T366 = T68[1'h1:1'h1];
  assign T367 = T388 ? T378 : T368;
  assign T368 = T377 ? counts_53 : counts_52;
  assign T10397 = reset ? 4'h0 : T369;
  assign T369 = T371 ? T52 : T370;
  assign T370 = io_resetCounts ? 4'h0 : counts_52;
  assign T371 = T10320 & T372;
  assign T372 = T76[6'h34:6'h34];
  assign T10398 = reset ? 4'h0 : T373;
  assign T373 = T375 ? T52 : T374;
  assign T374 = io_resetCounts ? 4'h0 : counts_53;
  assign T375 = T10320 & T376;
  assign T376 = T76[6'h35:6'h35];
  assign T377 = T68[1'h0:1'h0];
  assign T378 = T387 ? counts_55 : counts_54;
  assign T10399 = reset ? 4'h0 : T379;
  assign T379 = T381 ? T52 : T380;
  assign T380 = io_resetCounts ? 4'h0 : counts_54;
  assign T381 = T10320 & T382;
  assign T382 = T76[6'h36:6'h36];
  assign T10400 = reset ? 4'h0 : T383;
  assign T383 = T385 ? T52 : T384;
  assign T384 = io_resetCounts ? 4'h0 : counts_55;
  assign T385 = T10320 & T386;
  assign T386 = T76[6'h37:6'h37];
  assign T387 = T68[1'h0:1'h0];
  assign T388 = T68[1'h1:1'h1];
  assign T389 = T68[2'h2:2'h2];
  assign T390 = T435 ? T413 : T391;
  assign T391 = T412 ? T402 : T392;
  assign T392 = T401 ? counts_57 : counts_56;
  assign T10401 = reset ? 4'h0 : T393;
  assign T393 = T395 ? T52 : T394;
  assign T394 = io_resetCounts ? 4'h0 : counts_56;
  assign T395 = T10320 & T396;
  assign T396 = T76[6'h38:6'h38];
  assign T10402 = reset ? 4'h0 : T397;
  assign T397 = T399 ? T52 : T398;
  assign T398 = io_resetCounts ? 4'h0 : counts_57;
  assign T399 = T10320 & T400;
  assign T400 = T76[6'h39:6'h39];
  assign T401 = T68[1'h0:1'h0];
  assign T402 = T411 ? counts_59 : counts_58;
  assign T10403 = reset ? 4'h0 : T403;
  assign T403 = T405 ? T52 : T404;
  assign T404 = io_resetCounts ? 4'h0 : counts_58;
  assign T405 = T10320 & T406;
  assign T406 = T76[6'h3a:6'h3a];
  assign T10404 = reset ? 4'h0 : T407;
  assign T407 = T409 ? T52 : T408;
  assign T408 = io_resetCounts ? 4'h0 : counts_59;
  assign T409 = T10320 & T410;
  assign T410 = T76[6'h3b:6'h3b];
  assign T411 = T68[1'h0:1'h0];
  assign T412 = T68[1'h1:1'h1];
  assign T413 = T434 ? T424 : T414;
  assign T414 = T423 ? counts_61 : counts_60;
  assign T10405 = reset ? 4'h0 : T415;
  assign T415 = T417 ? T52 : T416;
  assign T416 = io_resetCounts ? 4'h0 : counts_60;
  assign T417 = T10320 & T418;
  assign T418 = T76[6'h3c:6'h3c];
  assign T10406 = reset ? 4'h0 : T419;
  assign T419 = T421 ? T52 : T420;
  assign T420 = io_resetCounts ? 4'h0 : counts_61;
  assign T421 = T10320 & T422;
  assign T422 = T76[6'h3d:6'h3d];
  assign T423 = T68[1'h0:1'h0];
  assign T424 = T433 ? counts_63 : counts_62;
  assign T10407 = reset ? 4'h0 : T425;
  assign T425 = T427 ? T52 : T426;
  assign T426 = io_resetCounts ? 4'h0 : counts_62;
  assign T427 = T10320 & T428;
  assign T428 = T76[6'h3e:6'h3e];
  assign T10408 = reset ? 4'h0 : T429;
  assign T429 = T431 ? T52 : T430;
  assign T430 = io_resetCounts ? 4'h0 : counts_63;
  assign T431 = T10320 & T432;
  assign T432 = T76[6'h3f:6'h3f];
  assign T433 = T68[1'h0:1'h0];
  assign T434 = T68[1'h1:1'h1];
  assign T435 = T68[2'h2:2'h2];
  assign T436 = T68[2'h3:2'h3];
  assign T437 = T68[3'h4:3'h4];
  assign T438 = T68[3'h5:3'h5];
  assign T439 = T820 ? T630 : T440;
  assign T440 = T629 ? T535 : T441;
  assign T441 = T534 ? T488 : T442;
  assign T442 = T487 ? T465 : T443;
  assign T443 = T464 ? T454 : T444;
  assign T444 = T453 ? counts_65 : counts_64;
  assign T10409 = reset ? 4'h0 : T445;
  assign T445 = T447 ? T52 : T446;
  assign T446 = io_resetCounts ? 4'h0 : counts_64;
  assign T447 = T10320 & T448;
  assign T448 = T76[7'h40:7'h40];
  assign T10410 = reset ? 4'h0 : T449;
  assign T449 = T451 ? T52 : T450;
  assign T450 = io_resetCounts ? 4'h0 : counts_65;
  assign T451 = T10320 & T452;
  assign T452 = T76[7'h41:7'h41];
  assign T453 = T68[1'h0:1'h0];
  assign T454 = T463 ? counts_67 : counts_66;
  assign T10411 = reset ? 4'h0 : T455;
  assign T455 = T457 ? T52 : T456;
  assign T456 = io_resetCounts ? 4'h0 : counts_66;
  assign T457 = T10320 & T458;
  assign T458 = T76[7'h42:7'h42];
  assign T10412 = reset ? 4'h0 : T459;
  assign T459 = T461 ? T52 : T460;
  assign T460 = io_resetCounts ? 4'h0 : counts_67;
  assign T461 = T10320 & T462;
  assign T462 = T76[7'h43:7'h43];
  assign T463 = T68[1'h0:1'h0];
  assign T464 = T68[1'h1:1'h1];
  assign T465 = T486 ? T476 : T466;
  assign T466 = T475 ? counts_69 : counts_68;
  assign T10413 = reset ? 4'h0 : T467;
  assign T467 = T469 ? T52 : T468;
  assign T468 = io_resetCounts ? 4'h0 : counts_68;
  assign T469 = T10320 & T470;
  assign T470 = T76[7'h44:7'h44];
  assign T10414 = reset ? 4'h0 : T471;
  assign T471 = T473 ? T52 : T472;
  assign T472 = io_resetCounts ? 4'h0 : counts_69;
  assign T473 = T10320 & T474;
  assign T474 = T76[7'h45:7'h45];
  assign T475 = T68[1'h0:1'h0];
  assign T476 = T485 ? counts_71 : counts_70;
  assign T10415 = reset ? 4'h0 : T477;
  assign T477 = T479 ? T52 : T478;
  assign T478 = io_resetCounts ? 4'h0 : counts_70;
  assign T479 = T10320 & T480;
  assign T480 = T76[7'h46:7'h46];
  assign T10416 = reset ? 4'h0 : T481;
  assign T481 = T483 ? T52 : T482;
  assign T482 = io_resetCounts ? 4'h0 : counts_71;
  assign T483 = T10320 & T484;
  assign T484 = T76[7'h47:7'h47];
  assign T485 = T68[1'h0:1'h0];
  assign T486 = T68[1'h1:1'h1];
  assign T487 = T68[2'h2:2'h2];
  assign T488 = T533 ? T511 : T489;
  assign T489 = T510 ? T500 : T490;
  assign T490 = T499 ? counts_73 : counts_72;
  assign T10417 = reset ? 4'h0 : T491;
  assign T491 = T493 ? T52 : T492;
  assign T492 = io_resetCounts ? 4'h0 : counts_72;
  assign T493 = T10320 & T494;
  assign T494 = T76[7'h48:7'h48];
  assign T10418 = reset ? 4'h0 : T495;
  assign T495 = T497 ? T52 : T496;
  assign T496 = io_resetCounts ? 4'h0 : counts_73;
  assign T497 = T10320 & T498;
  assign T498 = T76[7'h49:7'h49];
  assign T499 = T68[1'h0:1'h0];
  assign T500 = T509 ? counts_75 : counts_74;
  assign T10419 = reset ? 4'h0 : T501;
  assign T501 = T503 ? T52 : T502;
  assign T502 = io_resetCounts ? 4'h0 : counts_74;
  assign T503 = T10320 & T504;
  assign T504 = T76[7'h4a:7'h4a];
  assign T10420 = reset ? 4'h0 : T505;
  assign T505 = T507 ? T52 : T506;
  assign T506 = io_resetCounts ? 4'h0 : counts_75;
  assign T507 = T10320 & T508;
  assign T508 = T76[7'h4b:7'h4b];
  assign T509 = T68[1'h0:1'h0];
  assign T510 = T68[1'h1:1'h1];
  assign T511 = T532 ? T522 : T512;
  assign T512 = T521 ? counts_77 : counts_76;
  assign T10421 = reset ? 4'h0 : T513;
  assign T513 = T515 ? T52 : T514;
  assign T514 = io_resetCounts ? 4'h0 : counts_76;
  assign T515 = T10320 & T516;
  assign T516 = T76[7'h4c:7'h4c];
  assign T10422 = reset ? 4'h0 : T517;
  assign T517 = T519 ? T52 : T518;
  assign T518 = io_resetCounts ? 4'h0 : counts_77;
  assign T519 = T10320 & T520;
  assign T520 = T76[7'h4d:7'h4d];
  assign T521 = T68[1'h0:1'h0];
  assign T522 = T531 ? counts_79 : counts_78;
  assign T10423 = reset ? 4'h0 : T523;
  assign T523 = T525 ? T52 : T524;
  assign T524 = io_resetCounts ? 4'h0 : counts_78;
  assign T525 = T10320 & T526;
  assign T526 = T76[7'h4e:7'h4e];
  assign T10424 = reset ? 4'h0 : T527;
  assign T527 = T529 ? T52 : T528;
  assign T528 = io_resetCounts ? 4'h0 : counts_79;
  assign T529 = T10320 & T530;
  assign T530 = T76[7'h4f:7'h4f];
  assign T531 = T68[1'h0:1'h0];
  assign T532 = T68[1'h1:1'h1];
  assign T533 = T68[2'h2:2'h2];
  assign T534 = T68[2'h3:2'h3];
  assign T535 = T628 ? T582 : T536;
  assign T536 = T581 ? T559 : T537;
  assign T537 = T558 ? T548 : T538;
  assign T538 = T547 ? counts_81 : counts_80;
  assign T10425 = reset ? 4'h0 : T539;
  assign T539 = T541 ? T52 : T540;
  assign T540 = io_resetCounts ? 4'h0 : counts_80;
  assign T541 = T10320 & T542;
  assign T542 = T76[7'h50:7'h50];
  assign T10426 = reset ? 4'h0 : T543;
  assign T543 = T545 ? T52 : T544;
  assign T544 = io_resetCounts ? 4'h0 : counts_81;
  assign T545 = T10320 & T546;
  assign T546 = T76[7'h51:7'h51];
  assign T547 = T68[1'h0:1'h0];
  assign T548 = T557 ? counts_83 : counts_82;
  assign T10427 = reset ? 4'h0 : T549;
  assign T549 = T551 ? T52 : T550;
  assign T550 = io_resetCounts ? 4'h0 : counts_82;
  assign T551 = T10320 & T552;
  assign T552 = T76[7'h52:7'h52];
  assign T10428 = reset ? 4'h0 : T553;
  assign T553 = T555 ? T52 : T554;
  assign T554 = io_resetCounts ? 4'h0 : counts_83;
  assign T555 = T10320 & T556;
  assign T556 = T76[7'h53:7'h53];
  assign T557 = T68[1'h0:1'h0];
  assign T558 = T68[1'h1:1'h1];
  assign T559 = T580 ? T570 : T560;
  assign T560 = T569 ? counts_85 : counts_84;
  assign T10429 = reset ? 4'h0 : T561;
  assign T561 = T563 ? T52 : T562;
  assign T562 = io_resetCounts ? 4'h0 : counts_84;
  assign T563 = T10320 & T564;
  assign T564 = T76[7'h54:7'h54];
  assign T10430 = reset ? 4'h0 : T565;
  assign T565 = T567 ? T52 : T566;
  assign T566 = io_resetCounts ? 4'h0 : counts_85;
  assign T567 = T10320 & T568;
  assign T568 = T76[7'h55:7'h55];
  assign T569 = T68[1'h0:1'h0];
  assign T570 = T579 ? counts_87 : counts_86;
  assign T10431 = reset ? 4'h0 : T571;
  assign T571 = T573 ? T52 : T572;
  assign T572 = io_resetCounts ? 4'h0 : counts_86;
  assign T573 = T10320 & T574;
  assign T574 = T76[7'h56:7'h56];
  assign T10432 = reset ? 4'h0 : T575;
  assign T575 = T577 ? T52 : T576;
  assign T576 = io_resetCounts ? 4'h0 : counts_87;
  assign T577 = T10320 & T578;
  assign T578 = T76[7'h57:7'h57];
  assign T579 = T68[1'h0:1'h0];
  assign T580 = T68[1'h1:1'h1];
  assign T581 = T68[2'h2:2'h2];
  assign T582 = T627 ? T605 : T583;
  assign T583 = T604 ? T594 : T584;
  assign T584 = T593 ? counts_89 : counts_88;
  assign T10433 = reset ? 4'h0 : T585;
  assign T585 = T587 ? T52 : T586;
  assign T586 = io_resetCounts ? 4'h0 : counts_88;
  assign T587 = T10320 & T588;
  assign T588 = T76[7'h58:7'h58];
  assign T10434 = reset ? 4'h0 : T589;
  assign T589 = T591 ? T52 : T590;
  assign T590 = io_resetCounts ? 4'h0 : counts_89;
  assign T591 = T10320 & T592;
  assign T592 = T76[7'h59:7'h59];
  assign T593 = T68[1'h0:1'h0];
  assign T594 = T603 ? counts_91 : counts_90;
  assign T10435 = reset ? 4'h0 : T595;
  assign T595 = T597 ? T52 : T596;
  assign T596 = io_resetCounts ? 4'h0 : counts_90;
  assign T597 = T10320 & T598;
  assign T598 = T76[7'h5a:7'h5a];
  assign T10436 = reset ? 4'h0 : T599;
  assign T599 = T601 ? T52 : T600;
  assign T600 = io_resetCounts ? 4'h0 : counts_91;
  assign T601 = T10320 & T602;
  assign T602 = T76[7'h5b:7'h5b];
  assign T603 = T68[1'h0:1'h0];
  assign T604 = T68[1'h1:1'h1];
  assign T605 = T626 ? T616 : T606;
  assign T606 = T615 ? counts_93 : counts_92;
  assign T10437 = reset ? 4'h0 : T607;
  assign T607 = T609 ? T52 : T608;
  assign T608 = io_resetCounts ? 4'h0 : counts_92;
  assign T609 = T10320 & T610;
  assign T610 = T76[7'h5c:7'h5c];
  assign T10438 = reset ? 4'h0 : T611;
  assign T611 = T613 ? T52 : T612;
  assign T612 = io_resetCounts ? 4'h0 : counts_93;
  assign T613 = T10320 & T614;
  assign T614 = T76[7'h5d:7'h5d];
  assign T615 = T68[1'h0:1'h0];
  assign T616 = T625 ? counts_95 : counts_94;
  assign T10439 = reset ? 4'h0 : T617;
  assign T617 = T619 ? T52 : T618;
  assign T618 = io_resetCounts ? 4'h0 : counts_94;
  assign T619 = T10320 & T620;
  assign T620 = T76[7'h5e:7'h5e];
  assign T10440 = reset ? 4'h0 : T621;
  assign T621 = T623 ? T52 : T622;
  assign T622 = io_resetCounts ? 4'h0 : counts_95;
  assign T623 = T10320 & T624;
  assign T624 = T76[7'h5f:7'h5f];
  assign T625 = T68[1'h0:1'h0];
  assign T626 = T68[1'h1:1'h1];
  assign T627 = T68[2'h2:2'h2];
  assign T628 = T68[2'h3:2'h3];
  assign T629 = T68[3'h4:3'h4];
  assign T630 = T819 ? T725 : T631;
  assign T631 = T724 ? T678 : T632;
  assign T632 = T677 ? T655 : T633;
  assign T633 = T654 ? T644 : T634;
  assign T634 = T643 ? counts_97 : counts_96;
  assign T10441 = reset ? 4'h0 : T635;
  assign T635 = T637 ? T52 : T636;
  assign T636 = io_resetCounts ? 4'h0 : counts_96;
  assign T637 = T10320 & T638;
  assign T638 = T76[7'h60:7'h60];
  assign T10442 = reset ? 4'h0 : T639;
  assign T639 = T641 ? T52 : T640;
  assign T640 = io_resetCounts ? 4'h0 : counts_97;
  assign T641 = T10320 & T642;
  assign T642 = T76[7'h61:7'h61];
  assign T643 = T68[1'h0:1'h0];
  assign T644 = T653 ? counts_99 : counts_98;
  assign T10443 = reset ? 4'h0 : T645;
  assign T645 = T647 ? T52 : T646;
  assign T646 = io_resetCounts ? 4'h0 : counts_98;
  assign T647 = T10320 & T648;
  assign T648 = T76[7'h62:7'h62];
  assign T10444 = reset ? 4'h0 : T649;
  assign T649 = T651 ? T52 : T650;
  assign T650 = io_resetCounts ? 4'h0 : counts_99;
  assign T651 = T10320 & T652;
  assign T652 = T76[7'h63:7'h63];
  assign T653 = T68[1'h0:1'h0];
  assign T654 = T68[1'h1:1'h1];
  assign T655 = T676 ? T666 : T656;
  assign T656 = T665 ? counts_101 : counts_100;
  assign T10445 = reset ? 4'h0 : T657;
  assign T657 = T659 ? T52 : T658;
  assign T658 = io_resetCounts ? 4'h0 : counts_100;
  assign T659 = T10320 & T660;
  assign T660 = T76[7'h64:7'h64];
  assign T10446 = reset ? 4'h0 : T661;
  assign T661 = T663 ? T52 : T662;
  assign T662 = io_resetCounts ? 4'h0 : counts_101;
  assign T663 = T10320 & T664;
  assign T664 = T76[7'h65:7'h65];
  assign T665 = T68[1'h0:1'h0];
  assign T666 = T675 ? counts_103 : counts_102;
  assign T10447 = reset ? 4'h0 : T667;
  assign T667 = T669 ? T52 : T668;
  assign T668 = io_resetCounts ? 4'h0 : counts_102;
  assign T669 = T10320 & T670;
  assign T670 = T76[7'h66:7'h66];
  assign T10448 = reset ? 4'h0 : T671;
  assign T671 = T673 ? T52 : T672;
  assign T672 = io_resetCounts ? 4'h0 : counts_103;
  assign T673 = T10320 & T674;
  assign T674 = T76[7'h67:7'h67];
  assign T675 = T68[1'h0:1'h0];
  assign T676 = T68[1'h1:1'h1];
  assign T677 = T68[2'h2:2'h2];
  assign T678 = T723 ? T701 : T679;
  assign T679 = T700 ? T690 : T680;
  assign T680 = T689 ? counts_105 : counts_104;
  assign T10449 = reset ? 4'h0 : T681;
  assign T681 = T683 ? T52 : T682;
  assign T682 = io_resetCounts ? 4'h0 : counts_104;
  assign T683 = T10320 & T684;
  assign T684 = T76[7'h68:7'h68];
  assign T10450 = reset ? 4'h0 : T685;
  assign T685 = T687 ? T52 : T686;
  assign T686 = io_resetCounts ? 4'h0 : counts_105;
  assign T687 = T10320 & T688;
  assign T688 = T76[7'h69:7'h69];
  assign T689 = T68[1'h0:1'h0];
  assign T690 = T699 ? counts_107 : counts_106;
  assign T10451 = reset ? 4'h0 : T691;
  assign T691 = T693 ? T52 : T692;
  assign T692 = io_resetCounts ? 4'h0 : counts_106;
  assign T693 = T10320 & T694;
  assign T694 = T76[7'h6a:7'h6a];
  assign T10452 = reset ? 4'h0 : T695;
  assign T695 = T697 ? T52 : T696;
  assign T696 = io_resetCounts ? 4'h0 : counts_107;
  assign T697 = T10320 & T698;
  assign T698 = T76[7'h6b:7'h6b];
  assign T699 = T68[1'h0:1'h0];
  assign T700 = T68[1'h1:1'h1];
  assign T701 = T722 ? T712 : T702;
  assign T702 = T711 ? counts_109 : counts_108;
  assign T10453 = reset ? 4'h0 : T703;
  assign T703 = T705 ? T52 : T704;
  assign T704 = io_resetCounts ? 4'h0 : counts_108;
  assign T705 = T10320 & T706;
  assign T706 = T76[7'h6c:7'h6c];
  assign T10454 = reset ? 4'h0 : T707;
  assign T707 = T709 ? T52 : T708;
  assign T708 = io_resetCounts ? 4'h0 : counts_109;
  assign T709 = T10320 & T710;
  assign T710 = T76[7'h6d:7'h6d];
  assign T711 = T68[1'h0:1'h0];
  assign T712 = T721 ? counts_111 : counts_110;
  assign T10455 = reset ? 4'h0 : T713;
  assign T713 = T715 ? T52 : T714;
  assign T714 = io_resetCounts ? 4'h0 : counts_110;
  assign T715 = T10320 & T716;
  assign T716 = T76[7'h6e:7'h6e];
  assign T10456 = reset ? 4'h0 : T717;
  assign T717 = T719 ? T52 : T718;
  assign T718 = io_resetCounts ? 4'h0 : counts_111;
  assign T719 = T10320 & T720;
  assign T720 = T76[7'h6f:7'h6f];
  assign T721 = T68[1'h0:1'h0];
  assign T722 = T68[1'h1:1'h1];
  assign T723 = T68[2'h2:2'h2];
  assign T724 = T68[2'h3:2'h3];
  assign T725 = T818 ? T772 : T726;
  assign T726 = T771 ? T749 : T727;
  assign T727 = T748 ? T738 : T728;
  assign T728 = T737 ? counts_113 : counts_112;
  assign T10457 = reset ? 4'h0 : T729;
  assign T729 = T731 ? T52 : T730;
  assign T730 = io_resetCounts ? 4'h0 : counts_112;
  assign T731 = T10320 & T732;
  assign T732 = T76[7'h70:7'h70];
  assign T10458 = reset ? 4'h0 : T733;
  assign T733 = T735 ? T52 : T734;
  assign T734 = io_resetCounts ? 4'h0 : counts_113;
  assign T735 = T10320 & T736;
  assign T736 = T76[7'h71:7'h71];
  assign T737 = T68[1'h0:1'h0];
  assign T738 = T747 ? counts_115 : counts_114;
  assign T10459 = reset ? 4'h0 : T739;
  assign T739 = T741 ? T52 : T740;
  assign T740 = io_resetCounts ? 4'h0 : counts_114;
  assign T741 = T10320 & T742;
  assign T742 = T76[7'h72:7'h72];
  assign T10460 = reset ? 4'h0 : T743;
  assign T743 = T745 ? T52 : T744;
  assign T744 = io_resetCounts ? 4'h0 : counts_115;
  assign T745 = T10320 & T746;
  assign T746 = T76[7'h73:7'h73];
  assign T747 = T68[1'h0:1'h0];
  assign T748 = T68[1'h1:1'h1];
  assign T749 = T770 ? T760 : T750;
  assign T750 = T759 ? counts_117 : counts_116;
  assign T10461 = reset ? 4'h0 : T751;
  assign T751 = T753 ? T52 : T752;
  assign T752 = io_resetCounts ? 4'h0 : counts_116;
  assign T753 = T10320 & T754;
  assign T754 = T76[7'h74:7'h74];
  assign T10462 = reset ? 4'h0 : T755;
  assign T755 = T757 ? T52 : T756;
  assign T756 = io_resetCounts ? 4'h0 : counts_117;
  assign T757 = T10320 & T758;
  assign T758 = T76[7'h75:7'h75];
  assign T759 = T68[1'h0:1'h0];
  assign T760 = T769 ? counts_119 : counts_118;
  assign T10463 = reset ? 4'h0 : T761;
  assign T761 = T763 ? T52 : T762;
  assign T762 = io_resetCounts ? 4'h0 : counts_118;
  assign T763 = T10320 & T764;
  assign T764 = T76[7'h76:7'h76];
  assign T10464 = reset ? 4'h0 : T765;
  assign T765 = T767 ? T52 : T766;
  assign T766 = io_resetCounts ? 4'h0 : counts_119;
  assign T767 = T10320 & T768;
  assign T768 = T76[7'h77:7'h77];
  assign T769 = T68[1'h0:1'h0];
  assign T770 = T68[1'h1:1'h1];
  assign T771 = T68[2'h2:2'h2];
  assign T772 = T817 ? T795 : T773;
  assign T773 = T794 ? T784 : T774;
  assign T774 = T783 ? counts_121 : counts_120;
  assign T10465 = reset ? 4'h0 : T775;
  assign T775 = T777 ? T52 : T776;
  assign T776 = io_resetCounts ? 4'h0 : counts_120;
  assign T777 = T10320 & T778;
  assign T778 = T76[7'h78:7'h78];
  assign T10466 = reset ? 4'h0 : T779;
  assign T779 = T781 ? T52 : T780;
  assign T780 = io_resetCounts ? 4'h0 : counts_121;
  assign T781 = T10320 & T782;
  assign T782 = T76[7'h79:7'h79];
  assign T783 = T68[1'h0:1'h0];
  assign T784 = T793 ? counts_123 : counts_122;
  assign T10467 = reset ? 4'h0 : T785;
  assign T785 = T787 ? T52 : T786;
  assign T786 = io_resetCounts ? 4'h0 : counts_122;
  assign T787 = T10320 & T788;
  assign T788 = T76[7'h7a:7'h7a];
  assign T10468 = reset ? 4'h0 : T789;
  assign T789 = T791 ? T52 : T790;
  assign T790 = io_resetCounts ? 4'h0 : counts_123;
  assign T791 = T10320 & T792;
  assign T792 = T76[7'h7b:7'h7b];
  assign T793 = T68[1'h0:1'h0];
  assign T794 = T68[1'h1:1'h1];
  assign T795 = T816 ? T806 : T796;
  assign T796 = T805 ? counts_125 : counts_124;
  assign T10469 = reset ? 4'h0 : T797;
  assign T797 = T799 ? T52 : T798;
  assign T798 = io_resetCounts ? 4'h0 : counts_124;
  assign T799 = T10320 & T800;
  assign T800 = T76[7'h7c:7'h7c];
  assign T10470 = reset ? 4'h0 : T801;
  assign T801 = T803 ? T52 : T802;
  assign T802 = io_resetCounts ? 4'h0 : counts_125;
  assign T803 = T10320 & T804;
  assign T804 = T76[7'h7d:7'h7d];
  assign T805 = T68[1'h0:1'h0];
  assign T806 = T815 ? counts_127 : counts_126;
  assign T10471 = reset ? 4'h0 : T807;
  assign T807 = T809 ? T52 : T808;
  assign T808 = io_resetCounts ? 4'h0 : counts_126;
  assign T809 = T10320 & T810;
  assign T810 = T76[7'h7e:7'h7e];
  assign T10472 = reset ? 4'h0 : T811;
  assign T811 = T813 ? T52 : T812;
  assign T812 = io_resetCounts ? 4'h0 : counts_127;
  assign T813 = T10320 & T814;
  assign T814 = T76[7'h7f:7'h7f];
  assign T815 = T68[1'h0:1'h0];
  assign T816 = T68[1'h1:1'h1];
  assign T817 = T68[2'h2:2'h2];
  assign T818 = T68[2'h3:2'h3];
  assign T819 = T68[3'h4:3'h4];
  assign T820 = T68[3'h5:3'h5];
  assign T821 = T68[3'h6:3'h6];
  assign T822 = T1587 ? T1205 : T823;
  assign T823 = T1204 ? T1014 : T824;
  assign T824 = T1013 ? T919 : T825;
  assign T825 = T918 ? T872 : T826;
  assign T826 = T871 ? T849 : T827;
  assign T827 = T848 ? T838 : T828;
  assign T828 = T837 ? counts_129 : counts_128;
  assign T10473 = reset ? 4'h0 : T829;
  assign T829 = T831 ? T52 : T830;
  assign T830 = io_resetCounts ? 4'h0 : counts_128;
  assign T831 = T10320 & T832;
  assign T832 = T76[8'h80:8'h80];
  assign T10474 = reset ? 4'h0 : T833;
  assign T833 = T835 ? T52 : T834;
  assign T834 = io_resetCounts ? 4'h0 : counts_129;
  assign T835 = T10320 & T836;
  assign T836 = T76[8'h81:8'h81];
  assign T837 = T68[1'h0:1'h0];
  assign T838 = T847 ? counts_131 : counts_130;
  assign T10475 = reset ? 4'h0 : T839;
  assign T839 = T841 ? T52 : T840;
  assign T840 = io_resetCounts ? 4'h0 : counts_130;
  assign T841 = T10320 & T842;
  assign T842 = T76[8'h82:8'h82];
  assign T10476 = reset ? 4'h0 : T843;
  assign T843 = T845 ? T52 : T844;
  assign T844 = io_resetCounts ? 4'h0 : counts_131;
  assign T845 = T10320 & T846;
  assign T846 = T76[8'h83:8'h83];
  assign T847 = T68[1'h0:1'h0];
  assign T848 = T68[1'h1:1'h1];
  assign T849 = T870 ? T860 : T850;
  assign T850 = T859 ? counts_133 : counts_132;
  assign T10477 = reset ? 4'h0 : T851;
  assign T851 = T853 ? T52 : T852;
  assign T852 = io_resetCounts ? 4'h0 : counts_132;
  assign T853 = T10320 & T854;
  assign T854 = T76[8'h84:8'h84];
  assign T10478 = reset ? 4'h0 : T855;
  assign T855 = T857 ? T52 : T856;
  assign T856 = io_resetCounts ? 4'h0 : counts_133;
  assign T857 = T10320 & T858;
  assign T858 = T76[8'h85:8'h85];
  assign T859 = T68[1'h0:1'h0];
  assign T860 = T869 ? counts_135 : counts_134;
  assign T10479 = reset ? 4'h0 : T861;
  assign T861 = T863 ? T52 : T862;
  assign T862 = io_resetCounts ? 4'h0 : counts_134;
  assign T863 = T10320 & T864;
  assign T864 = T76[8'h86:8'h86];
  assign T10480 = reset ? 4'h0 : T865;
  assign T865 = T867 ? T52 : T866;
  assign T866 = io_resetCounts ? 4'h0 : counts_135;
  assign T867 = T10320 & T868;
  assign T868 = T76[8'h87:8'h87];
  assign T869 = T68[1'h0:1'h0];
  assign T870 = T68[1'h1:1'h1];
  assign T871 = T68[2'h2:2'h2];
  assign T872 = T917 ? T895 : T873;
  assign T873 = T894 ? T884 : T874;
  assign T874 = T883 ? counts_137 : counts_136;
  assign T10481 = reset ? 4'h0 : T875;
  assign T875 = T877 ? T52 : T876;
  assign T876 = io_resetCounts ? 4'h0 : counts_136;
  assign T877 = T10320 & T878;
  assign T878 = T76[8'h88:8'h88];
  assign T10482 = reset ? 4'h0 : T879;
  assign T879 = T881 ? T52 : T880;
  assign T880 = io_resetCounts ? 4'h0 : counts_137;
  assign T881 = T10320 & T882;
  assign T882 = T76[8'h89:8'h89];
  assign T883 = T68[1'h0:1'h0];
  assign T884 = T893 ? counts_139 : counts_138;
  assign T10483 = reset ? 4'h0 : T885;
  assign T885 = T887 ? T52 : T886;
  assign T886 = io_resetCounts ? 4'h0 : counts_138;
  assign T887 = T10320 & T888;
  assign T888 = T76[8'h8a:8'h8a];
  assign T10484 = reset ? 4'h0 : T889;
  assign T889 = T891 ? T52 : T890;
  assign T890 = io_resetCounts ? 4'h0 : counts_139;
  assign T891 = T10320 & T892;
  assign T892 = T76[8'h8b:8'h8b];
  assign T893 = T68[1'h0:1'h0];
  assign T894 = T68[1'h1:1'h1];
  assign T895 = T916 ? T906 : T896;
  assign T896 = T905 ? counts_141 : counts_140;
  assign T10485 = reset ? 4'h0 : T897;
  assign T897 = T899 ? T52 : T898;
  assign T898 = io_resetCounts ? 4'h0 : counts_140;
  assign T899 = T10320 & T900;
  assign T900 = T76[8'h8c:8'h8c];
  assign T10486 = reset ? 4'h0 : T901;
  assign T901 = T903 ? T52 : T902;
  assign T902 = io_resetCounts ? 4'h0 : counts_141;
  assign T903 = T10320 & T904;
  assign T904 = T76[8'h8d:8'h8d];
  assign T905 = T68[1'h0:1'h0];
  assign T906 = T915 ? counts_143 : counts_142;
  assign T10487 = reset ? 4'h0 : T907;
  assign T907 = T909 ? T52 : T908;
  assign T908 = io_resetCounts ? 4'h0 : counts_142;
  assign T909 = T10320 & T910;
  assign T910 = T76[8'h8e:8'h8e];
  assign T10488 = reset ? 4'h0 : T911;
  assign T911 = T913 ? T52 : T912;
  assign T912 = io_resetCounts ? 4'h0 : counts_143;
  assign T913 = T10320 & T914;
  assign T914 = T76[8'h8f:8'h8f];
  assign T915 = T68[1'h0:1'h0];
  assign T916 = T68[1'h1:1'h1];
  assign T917 = T68[2'h2:2'h2];
  assign T918 = T68[2'h3:2'h3];
  assign T919 = T1012 ? T966 : T920;
  assign T920 = T965 ? T943 : T921;
  assign T921 = T942 ? T932 : T922;
  assign T922 = T931 ? counts_145 : counts_144;
  assign T10489 = reset ? 4'h0 : T923;
  assign T923 = T925 ? T52 : T924;
  assign T924 = io_resetCounts ? 4'h0 : counts_144;
  assign T925 = T10320 & T926;
  assign T926 = T76[8'h90:8'h90];
  assign T10490 = reset ? 4'h0 : T927;
  assign T927 = T929 ? T52 : T928;
  assign T928 = io_resetCounts ? 4'h0 : counts_145;
  assign T929 = T10320 & T930;
  assign T930 = T76[8'h91:8'h91];
  assign T931 = T68[1'h0:1'h0];
  assign T932 = T941 ? counts_147 : counts_146;
  assign T10491 = reset ? 4'h0 : T933;
  assign T933 = T935 ? T52 : T934;
  assign T934 = io_resetCounts ? 4'h0 : counts_146;
  assign T935 = T10320 & T936;
  assign T936 = T76[8'h92:8'h92];
  assign T10492 = reset ? 4'h0 : T937;
  assign T937 = T939 ? T52 : T938;
  assign T938 = io_resetCounts ? 4'h0 : counts_147;
  assign T939 = T10320 & T940;
  assign T940 = T76[8'h93:8'h93];
  assign T941 = T68[1'h0:1'h0];
  assign T942 = T68[1'h1:1'h1];
  assign T943 = T964 ? T954 : T944;
  assign T944 = T953 ? counts_149 : counts_148;
  assign T10493 = reset ? 4'h0 : T945;
  assign T945 = T947 ? T52 : T946;
  assign T946 = io_resetCounts ? 4'h0 : counts_148;
  assign T947 = T10320 & T948;
  assign T948 = T76[8'h94:8'h94];
  assign T10494 = reset ? 4'h0 : T949;
  assign T949 = T951 ? T52 : T950;
  assign T950 = io_resetCounts ? 4'h0 : counts_149;
  assign T951 = T10320 & T952;
  assign T952 = T76[8'h95:8'h95];
  assign T953 = T68[1'h0:1'h0];
  assign T954 = T963 ? counts_151 : counts_150;
  assign T10495 = reset ? 4'h0 : T955;
  assign T955 = T957 ? T52 : T956;
  assign T956 = io_resetCounts ? 4'h0 : counts_150;
  assign T957 = T10320 & T958;
  assign T958 = T76[8'h96:8'h96];
  assign T10496 = reset ? 4'h0 : T959;
  assign T959 = T961 ? T52 : T960;
  assign T960 = io_resetCounts ? 4'h0 : counts_151;
  assign T961 = T10320 & T962;
  assign T962 = T76[8'h97:8'h97];
  assign T963 = T68[1'h0:1'h0];
  assign T964 = T68[1'h1:1'h1];
  assign T965 = T68[2'h2:2'h2];
  assign T966 = T1011 ? T989 : T967;
  assign T967 = T988 ? T978 : T968;
  assign T968 = T977 ? counts_153 : counts_152;
  assign T10497 = reset ? 4'h0 : T969;
  assign T969 = T971 ? T52 : T970;
  assign T970 = io_resetCounts ? 4'h0 : counts_152;
  assign T971 = T10320 & T972;
  assign T972 = T76[8'h98:8'h98];
  assign T10498 = reset ? 4'h0 : T973;
  assign T973 = T975 ? T52 : T974;
  assign T974 = io_resetCounts ? 4'h0 : counts_153;
  assign T975 = T10320 & T976;
  assign T976 = T76[8'h99:8'h99];
  assign T977 = T68[1'h0:1'h0];
  assign T978 = T987 ? counts_155 : counts_154;
  assign T10499 = reset ? 4'h0 : T979;
  assign T979 = T981 ? T52 : T980;
  assign T980 = io_resetCounts ? 4'h0 : counts_154;
  assign T981 = T10320 & T982;
  assign T982 = T76[8'h9a:8'h9a];
  assign T10500 = reset ? 4'h0 : T983;
  assign T983 = T985 ? T52 : T984;
  assign T984 = io_resetCounts ? 4'h0 : counts_155;
  assign T985 = T10320 & T986;
  assign T986 = T76[8'h9b:8'h9b];
  assign T987 = T68[1'h0:1'h0];
  assign T988 = T68[1'h1:1'h1];
  assign T989 = T1010 ? T1000 : T990;
  assign T990 = T999 ? counts_157 : counts_156;
  assign T10501 = reset ? 4'h0 : T991;
  assign T991 = T993 ? T52 : T992;
  assign T992 = io_resetCounts ? 4'h0 : counts_156;
  assign T993 = T10320 & T994;
  assign T994 = T76[8'h9c:8'h9c];
  assign T10502 = reset ? 4'h0 : T995;
  assign T995 = T997 ? T52 : T996;
  assign T996 = io_resetCounts ? 4'h0 : counts_157;
  assign T997 = T10320 & T998;
  assign T998 = T76[8'h9d:8'h9d];
  assign T999 = T68[1'h0:1'h0];
  assign T1000 = T1009 ? counts_159 : counts_158;
  assign T10503 = reset ? 4'h0 : T1001;
  assign T1001 = T1003 ? T52 : T1002;
  assign T1002 = io_resetCounts ? 4'h0 : counts_158;
  assign T1003 = T10320 & T1004;
  assign T1004 = T76[8'h9e:8'h9e];
  assign T10504 = reset ? 4'h0 : T1005;
  assign T1005 = T1007 ? T52 : T1006;
  assign T1006 = io_resetCounts ? 4'h0 : counts_159;
  assign T1007 = T10320 & T1008;
  assign T1008 = T76[8'h9f:8'h9f];
  assign T1009 = T68[1'h0:1'h0];
  assign T1010 = T68[1'h1:1'h1];
  assign T1011 = T68[2'h2:2'h2];
  assign T1012 = T68[2'h3:2'h3];
  assign T1013 = T68[3'h4:3'h4];
  assign T1014 = T1203 ? T1109 : T1015;
  assign T1015 = T1108 ? T1062 : T1016;
  assign T1016 = T1061 ? T1039 : T1017;
  assign T1017 = T1038 ? T1028 : T1018;
  assign T1018 = T1027 ? counts_161 : counts_160;
  assign T10505 = reset ? 4'h0 : T1019;
  assign T1019 = T1021 ? T52 : T1020;
  assign T1020 = io_resetCounts ? 4'h0 : counts_160;
  assign T1021 = T10320 & T1022;
  assign T1022 = T76[8'ha0:8'ha0];
  assign T10506 = reset ? 4'h0 : T1023;
  assign T1023 = T1025 ? T52 : T1024;
  assign T1024 = io_resetCounts ? 4'h0 : counts_161;
  assign T1025 = T10320 & T1026;
  assign T1026 = T76[8'ha1:8'ha1];
  assign T1027 = T68[1'h0:1'h0];
  assign T1028 = T1037 ? counts_163 : counts_162;
  assign T10507 = reset ? 4'h0 : T1029;
  assign T1029 = T1031 ? T52 : T1030;
  assign T1030 = io_resetCounts ? 4'h0 : counts_162;
  assign T1031 = T10320 & T1032;
  assign T1032 = T76[8'ha2:8'ha2];
  assign T10508 = reset ? 4'h0 : T1033;
  assign T1033 = T1035 ? T52 : T1034;
  assign T1034 = io_resetCounts ? 4'h0 : counts_163;
  assign T1035 = T10320 & T1036;
  assign T1036 = T76[8'ha3:8'ha3];
  assign T1037 = T68[1'h0:1'h0];
  assign T1038 = T68[1'h1:1'h1];
  assign T1039 = T1060 ? T1050 : T1040;
  assign T1040 = T1049 ? counts_165 : counts_164;
  assign T10509 = reset ? 4'h0 : T1041;
  assign T1041 = T1043 ? T52 : T1042;
  assign T1042 = io_resetCounts ? 4'h0 : counts_164;
  assign T1043 = T10320 & T1044;
  assign T1044 = T76[8'ha4:8'ha4];
  assign T10510 = reset ? 4'h0 : T1045;
  assign T1045 = T1047 ? T52 : T1046;
  assign T1046 = io_resetCounts ? 4'h0 : counts_165;
  assign T1047 = T10320 & T1048;
  assign T1048 = T76[8'ha5:8'ha5];
  assign T1049 = T68[1'h0:1'h0];
  assign T1050 = T1059 ? counts_167 : counts_166;
  assign T10511 = reset ? 4'h0 : T1051;
  assign T1051 = T1053 ? T52 : T1052;
  assign T1052 = io_resetCounts ? 4'h0 : counts_166;
  assign T1053 = T10320 & T1054;
  assign T1054 = T76[8'ha6:8'ha6];
  assign T10512 = reset ? 4'h0 : T1055;
  assign T1055 = T1057 ? T52 : T1056;
  assign T1056 = io_resetCounts ? 4'h0 : counts_167;
  assign T1057 = T10320 & T1058;
  assign T1058 = T76[8'ha7:8'ha7];
  assign T1059 = T68[1'h0:1'h0];
  assign T1060 = T68[1'h1:1'h1];
  assign T1061 = T68[2'h2:2'h2];
  assign T1062 = T1107 ? T1085 : T1063;
  assign T1063 = T1084 ? T1074 : T1064;
  assign T1064 = T1073 ? counts_169 : counts_168;
  assign T10513 = reset ? 4'h0 : T1065;
  assign T1065 = T1067 ? T52 : T1066;
  assign T1066 = io_resetCounts ? 4'h0 : counts_168;
  assign T1067 = T10320 & T1068;
  assign T1068 = T76[8'ha8:8'ha8];
  assign T10514 = reset ? 4'h0 : T1069;
  assign T1069 = T1071 ? T52 : T1070;
  assign T1070 = io_resetCounts ? 4'h0 : counts_169;
  assign T1071 = T10320 & T1072;
  assign T1072 = T76[8'ha9:8'ha9];
  assign T1073 = T68[1'h0:1'h0];
  assign T1074 = T1083 ? counts_171 : counts_170;
  assign T10515 = reset ? 4'h0 : T1075;
  assign T1075 = T1077 ? T52 : T1076;
  assign T1076 = io_resetCounts ? 4'h0 : counts_170;
  assign T1077 = T10320 & T1078;
  assign T1078 = T76[8'haa:8'haa];
  assign T10516 = reset ? 4'h0 : T1079;
  assign T1079 = T1081 ? T52 : T1080;
  assign T1080 = io_resetCounts ? 4'h0 : counts_171;
  assign T1081 = T10320 & T1082;
  assign T1082 = T76[8'hab:8'hab];
  assign T1083 = T68[1'h0:1'h0];
  assign T1084 = T68[1'h1:1'h1];
  assign T1085 = T1106 ? T1096 : T1086;
  assign T1086 = T1095 ? counts_173 : counts_172;
  assign T10517 = reset ? 4'h0 : T1087;
  assign T1087 = T1089 ? T52 : T1088;
  assign T1088 = io_resetCounts ? 4'h0 : counts_172;
  assign T1089 = T10320 & T1090;
  assign T1090 = T76[8'hac:8'hac];
  assign T10518 = reset ? 4'h0 : T1091;
  assign T1091 = T1093 ? T52 : T1092;
  assign T1092 = io_resetCounts ? 4'h0 : counts_173;
  assign T1093 = T10320 & T1094;
  assign T1094 = T76[8'had:8'had];
  assign T1095 = T68[1'h0:1'h0];
  assign T1096 = T1105 ? counts_175 : counts_174;
  assign T10519 = reset ? 4'h0 : T1097;
  assign T1097 = T1099 ? T52 : T1098;
  assign T1098 = io_resetCounts ? 4'h0 : counts_174;
  assign T1099 = T10320 & T1100;
  assign T1100 = T76[8'hae:8'hae];
  assign T10520 = reset ? 4'h0 : T1101;
  assign T1101 = T1103 ? T52 : T1102;
  assign T1102 = io_resetCounts ? 4'h0 : counts_175;
  assign T1103 = T10320 & T1104;
  assign T1104 = T76[8'haf:8'haf];
  assign T1105 = T68[1'h0:1'h0];
  assign T1106 = T68[1'h1:1'h1];
  assign T1107 = T68[2'h2:2'h2];
  assign T1108 = T68[2'h3:2'h3];
  assign T1109 = T1202 ? T1156 : T1110;
  assign T1110 = T1155 ? T1133 : T1111;
  assign T1111 = T1132 ? T1122 : T1112;
  assign T1112 = T1121 ? counts_177 : counts_176;
  assign T10521 = reset ? 4'h0 : T1113;
  assign T1113 = T1115 ? T52 : T1114;
  assign T1114 = io_resetCounts ? 4'h0 : counts_176;
  assign T1115 = T10320 & T1116;
  assign T1116 = T76[8'hb0:8'hb0];
  assign T10522 = reset ? 4'h0 : T1117;
  assign T1117 = T1119 ? T52 : T1118;
  assign T1118 = io_resetCounts ? 4'h0 : counts_177;
  assign T1119 = T10320 & T1120;
  assign T1120 = T76[8'hb1:8'hb1];
  assign T1121 = T68[1'h0:1'h0];
  assign T1122 = T1131 ? counts_179 : counts_178;
  assign T10523 = reset ? 4'h0 : T1123;
  assign T1123 = T1125 ? T52 : T1124;
  assign T1124 = io_resetCounts ? 4'h0 : counts_178;
  assign T1125 = T10320 & T1126;
  assign T1126 = T76[8'hb2:8'hb2];
  assign T10524 = reset ? 4'h0 : T1127;
  assign T1127 = T1129 ? T52 : T1128;
  assign T1128 = io_resetCounts ? 4'h0 : counts_179;
  assign T1129 = T10320 & T1130;
  assign T1130 = T76[8'hb3:8'hb3];
  assign T1131 = T68[1'h0:1'h0];
  assign T1132 = T68[1'h1:1'h1];
  assign T1133 = T1154 ? T1144 : T1134;
  assign T1134 = T1143 ? counts_181 : counts_180;
  assign T10525 = reset ? 4'h0 : T1135;
  assign T1135 = T1137 ? T52 : T1136;
  assign T1136 = io_resetCounts ? 4'h0 : counts_180;
  assign T1137 = T10320 & T1138;
  assign T1138 = T76[8'hb4:8'hb4];
  assign T10526 = reset ? 4'h0 : T1139;
  assign T1139 = T1141 ? T52 : T1140;
  assign T1140 = io_resetCounts ? 4'h0 : counts_181;
  assign T1141 = T10320 & T1142;
  assign T1142 = T76[8'hb5:8'hb5];
  assign T1143 = T68[1'h0:1'h0];
  assign T1144 = T1153 ? counts_183 : counts_182;
  assign T10527 = reset ? 4'h0 : T1145;
  assign T1145 = T1147 ? T52 : T1146;
  assign T1146 = io_resetCounts ? 4'h0 : counts_182;
  assign T1147 = T10320 & T1148;
  assign T1148 = T76[8'hb6:8'hb6];
  assign T10528 = reset ? 4'h0 : T1149;
  assign T1149 = T1151 ? T52 : T1150;
  assign T1150 = io_resetCounts ? 4'h0 : counts_183;
  assign T1151 = T10320 & T1152;
  assign T1152 = T76[8'hb7:8'hb7];
  assign T1153 = T68[1'h0:1'h0];
  assign T1154 = T68[1'h1:1'h1];
  assign T1155 = T68[2'h2:2'h2];
  assign T1156 = T1201 ? T1179 : T1157;
  assign T1157 = T1178 ? T1168 : T1158;
  assign T1158 = T1167 ? counts_185 : counts_184;
  assign T10529 = reset ? 4'h0 : T1159;
  assign T1159 = T1161 ? T52 : T1160;
  assign T1160 = io_resetCounts ? 4'h0 : counts_184;
  assign T1161 = T10320 & T1162;
  assign T1162 = T76[8'hb8:8'hb8];
  assign T10530 = reset ? 4'h0 : T1163;
  assign T1163 = T1165 ? T52 : T1164;
  assign T1164 = io_resetCounts ? 4'h0 : counts_185;
  assign T1165 = T10320 & T1166;
  assign T1166 = T76[8'hb9:8'hb9];
  assign T1167 = T68[1'h0:1'h0];
  assign T1168 = T1177 ? counts_187 : counts_186;
  assign T10531 = reset ? 4'h0 : T1169;
  assign T1169 = T1171 ? T52 : T1170;
  assign T1170 = io_resetCounts ? 4'h0 : counts_186;
  assign T1171 = T10320 & T1172;
  assign T1172 = T76[8'hba:8'hba];
  assign T10532 = reset ? 4'h0 : T1173;
  assign T1173 = T1175 ? T52 : T1174;
  assign T1174 = io_resetCounts ? 4'h0 : counts_187;
  assign T1175 = T10320 & T1176;
  assign T1176 = T76[8'hbb:8'hbb];
  assign T1177 = T68[1'h0:1'h0];
  assign T1178 = T68[1'h1:1'h1];
  assign T1179 = T1200 ? T1190 : T1180;
  assign T1180 = T1189 ? counts_189 : counts_188;
  assign T10533 = reset ? 4'h0 : T1181;
  assign T1181 = T1183 ? T52 : T1182;
  assign T1182 = io_resetCounts ? 4'h0 : counts_188;
  assign T1183 = T10320 & T1184;
  assign T1184 = T76[8'hbc:8'hbc];
  assign T10534 = reset ? 4'h0 : T1185;
  assign T1185 = T1187 ? T52 : T1186;
  assign T1186 = io_resetCounts ? 4'h0 : counts_189;
  assign T1187 = T10320 & T1188;
  assign T1188 = T76[8'hbd:8'hbd];
  assign T1189 = T68[1'h0:1'h0];
  assign T1190 = T1199 ? counts_191 : counts_190;
  assign T10535 = reset ? 4'h0 : T1191;
  assign T1191 = T1193 ? T52 : T1192;
  assign T1192 = io_resetCounts ? 4'h0 : counts_190;
  assign T1193 = T10320 & T1194;
  assign T1194 = T76[8'hbe:8'hbe];
  assign T10536 = reset ? 4'h0 : T1195;
  assign T1195 = T1197 ? T52 : T1196;
  assign T1196 = io_resetCounts ? 4'h0 : counts_191;
  assign T1197 = T10320 & T1198;
  assign T1198 = T76[8'hbf:8'hbf];
  assign T1199 = T68[1'h0:1'h0];
  assign T1200 = T68[1'h1:1'h1];
  assign T1201 = T68[2'h2:2'h2];
  assign T1202 = T68[2'h3:2'h3];
  assign T1203 = T68[3'h4:3'h4];
  assign T1204 = T68[3'h5:3'h5];
  assign T1205 = T1586 ? T1396 : T1206;
  assign T1206 = T1395 ? T1301 : T1207;
  assign T1207 = T1300 ? T1254 : T1208;
  assign T1208 = T1253 ? T1231 : T1209;
  assign T1209 = T1230 ? T1220 : T1210;
  assign T1210 = T1219 ? counts_193 : counts_192;
  assign T10537 = reset ? 4'h0 : T1211;
  assign T1211 = T1213 ? T52 : T1212;
  assign T1212 = io_resetCounts ? 4'h0 : counts_192;
  assign T1213 = T10320 & T1214;
  assign T1214 = T76[8'hc0:8'hc0];
  assign T10538 = reset ? 4'h0 : T1215;
  assign T1215 = T1217 ? T52 : T1216;
  assign T1216 = io_resetCounts ? 4'h0 : counts_193;
  assign T1217 = T10320 & T1218;
  assign T1218 = T76[8'hc1:8'hc1];
  assign T1219 = T68[1'h0:1'h0];
  assign T1220 = T1229 ? counts_195 : counts_194;
  assign T10539 = reset ? 4'h0 : T1221;
  assign T1221 = T1223 ? T52 : T1222;
  assign T1222 = io_resetCounts ? 4'h0 : counts_194;
  assign T1223 = T10320 & T1224;
  assign T1224 = T76[8'hc2:8'hc2];
  assign T10540 = reset ? 4'h0 : T1225;
  assign T1225 = T1227 ? T52 : T1226;
  assign T1226 = io_resetCounts ? 4'h0 : counts_195;
  assign T1227 = T10320 & T1228;
  assign T1228 = T76[8'hc3:8'hc3];
  assign T1229 = T68[1'h0:1'h0];
  assign T1230 = T68[1'h1:1'h1];
  assign T1231 = T1252 ? T1242 : T1232;
  assign T1232 = T1241 ? counts_197 : counts_196;
  assign T10541 = reset ? 4'h0 : T1233;
  assign T1233 = T1235 ? T52 : T1234;
  assign T1234 = io_resetCounts ? 4'h0 : counts_196;
  assign T1235 = T10320 & T1236;
  assign T1236 = T76[8'hc4:8'hc4];
  assign T10542 = reset ? 4'h0 : T1237;
  assign T1237 = T1239 ? T52 : T1238;
  assign T1238 = io_resetCounts ? 4'h0 : counts_197;
  assign T1239 = T10320 & T1240;
  assign T1240 = T76[8'hc5:8'hc5];
  assign T1241 = T68[1'h0:1'h0];
  assign T1242 = T1251 ? counts_199 : counts_198;
  assign T10543 = reset ? 4'h0 : T1243;
  assign T1243 = T1245 ? T52 : T1244;
  assign T1244 = io_resetCounts ? 4'h0 : counts_198;
  assign T1245 = T10320 & T1246;
  assign T1246 = T76[8'hc6:8'hc6];
  assign T10544 = reset ? 4'h0 : T1247;
  assign T1247 = T1249 ? T52 : T1248;
  assign T1248 = io_resetCounts ? 4'h0 : counts_199;
  assign T1249 = T10320 & T1250;
  assign T1250 = T76[8'hc7:8'hc7];
  assign T1251 = T68[1'h0:1'h0];
  assign T1252 = T68[1'h1:1'h1];
  assign T1253 = T68[2'h2:2'h2];
  assign T1254 = T1299 ? T1277 : T1255;
  assign T1255 = T1276 ? T1266 : T1256;
  assign T1256 = T1265 ? counts_201 : counts_200;
  assign T10545 = reset ? 4'h0 : T1257;
  assign T1257 = T1259 ? T52 : T1258;
  assign T1258 = io_resetCounts ? 4'h0 : counts_200;
  assign T1259 = T10320 & T1260;
  assign T1260 = T76[8'hc8:8'hc8];
  assign T10546 = reset ? 4'h0 : T1261;
  assign T1261 = T1263 ? T52 : T1262;
  assign T1262 = io_resetCounts ? 4'h0 : counts_201;
  assign T1263 = T10320 & T1264;
  assign T1264 = T76[8'hc9:8'hc9];
  assign T1265 = T68[1'h0:1'h0];
  assign T1266 = T1275 ? counts_203 : counts_202;
  assign T10547 = reset ? 4'h0 : T1267;
  assign T1267 = T1269 ? T52 : T1268;
  assign T1268 = io_resetCounts ? 4'h0 : counts_202;
  assign T1269 = T10320 & T1270;
  assign T1270 = T76[8'hca:8'hca];
  assign T10548 = reset ? 4'h0 : T1271;
  assign T1271 = T1273 ? T52 : T1272;
  assign T1272 = io_resetCounts ? 4'h0 : counts_203;
  assign T1273 = T10320 & T1274;
  assign T1274 = T76[8'hcb:8'hcb];
  assign T1275 = T68[1'h0:1'h0];
  assign T1276 = T68[1'h1:1'h1];
  assign T1277 = T1298 ? T1288 : T1278;
  assign T1278 = T1287 ? counts_205 : counts_204;
  assign T10549 = reset ? 4'h0 : T1279;
  assign T1279 = T1281 ? T52 : T1280;
  assign T1280 = io_resetCounts ? 4'h0 : counts_204;
  assign T1281 = T10320 & T1282;
  assign T1282 = T76[8'hcc:8'hcc];
  assign T10550 = reset ? 4'h0 : T1283;
  assign T1283 = T1285 ? T52 : T1284;
  assign T1284 = io_resetCounts ? 4'h0 : counts_205;
  assign T1285 = T10320 & T1286;
  assign T1286 = T76[8'hcd:8'hcd];
  assign T1287 = T68[1'h0:1'h0];
  assign T1288 = T1297 ? counts_207 : counts_206;
  assign T10551 = reset ? 4'h0 : T1289;
  assign T1289 = T1291 ? T52 : T1290;
  assign T1290 = io_resetCounts ? 4'h0 : counts_206;
  assign T1291 = T10320 & T1292;
  assign T1292 = T76[8'hce:8'hce];
  assign T10552 = reset ? 4'h0 : T1293;
  assign T1293 = T1295 ? T52 : T1294;
  assign T1294 = io_resetCounts ? 4'h0 : counts_207;
  assign T1295 = T10320 & T1296;
  assign T1296 = T76[8'hcf:8'hcf];
  assign T1297 = T68[1'h0:1'h0];
  assign T1298 = T68[1'h1:1'h1];
  assign T1299 = T68[2'h2:2'h2];
  assign T1300 = T68[2'h3:2'h3];
  assign T1301 = T1394 ? T1348 : T1302;
  assign T1302 = T1347 ? T1325 : T1303;
  assign T1303 = T1324 ? T1314 : T1304;
  assign T1304 = T1313 ? counts_209 : counts_208;
  assign T10553 = reset ? 4'h0 : T1305;
  assign T1305 = T1307 ? T52 : T1306;
  assign T1306 = io_resetCounts ? 4'h0 : counts_208;
  assign T1307 = T10320 & T1308;
  assign T1308 = T76[8'hd0:8'hd0];
  assign T10554 = reset ? 4'h0 : T1309;
  assign T1309 = T1311 ? T52 : T1310;
  assign T1310 = io_resetCounts ? 4'h0 : counts_209;
  assign T1311 = T10320 & T1312;
  assign T1312 = T76[8'hd1:8'hd1];
  assign T1313 = T68[1'h0:1'h0];
  assign T1314 = T1323 ? counts_211 : counts_210;
  assign T10555 = reset ? 4'h0 : T1315;
  assign T1315 = T1317 ? T52 : T1316;
  assign T1316 = io_resetCounts ? 4'h0 : counts_210;
  assign T1317 = T10320 & T1318;
  assign T1318 = T76[8'hd2:8'hd2];
  assign T10556 = reset ? 4'h0 : T1319;
  assign T1319 = T1321 ? T52 : T1320;
  assign T1320 = io_resetCounts ? 4'h0 : counts_211;
  assign T1321 = T10320 & T1322;
  assign T1322 = T76[8'hd3:8'hd3];
  assign T1323 = T68[1'h0:1'h0];
  assign T1324 = T68[1'h1:1'h1];
  assign T1325 = T1346 ? T1336 : T1326;
  assign T1326 = T1335 ? counts_213 : counts_212;
  assign T10557 = reset ? 4'h0 : T1327;
  assign T1327 = T1329 ? T52 : T1328;
  assign T1328 = io_resetCounts ? 4'h0 : counts_212;
  assign T1329 = T10320 & T1330;
  assign T1330 = T76[8'hd4:8'hd4];
  assign T10558 = reset ? 4'h0 : T1331;
  assign T1331 = T1333 ? T52 : T1332;
  assign T1332 = io_resetCounts ? 4'h0 : counts_213;
  assign T1333 = T10320 & T1334;
  assign T1334 = T76[8'hd5:8'hd5];
  assign T1335 = T68[1'h0:1'h0];
  assign T1336 = T1345 ? counts_215 : counts_214;
  assign T10559 = reset ? 4'h0 : T1337;
  assign T1337 = T1339 ? T52 : T1338;
  assign T1338 = io_resetCounts ? 4'h0 : counts_214;
  assign T1339 = T10320 & T1340;
  assign T1340 = T76[8'hd6:8'hd6];
  assign T10560 = reset ? 4'h0 : T1341;
  assign T1341 = T1343 ? T52 : T1342;
  assign T1342 = io_resetCounts ? 4'h0 : counts_215;
  assign T1343 = T10320 & T1344;
  assign T1344 = T76[8'hd7:8'hd7];
  assign T1345 = T68[1'h0:1'h0];
  assign T1346 = T68[1'h1:1'h1];
  assign T1347 = T68[2'h2:2'h2];
  assign T1348 = T1393 ? T1371 : T1349;
  assign T1349 = T1370 ? T1360 : T1350;
  assign T1350 = T1359 ? counts_217 : counts_216;
  assign T10561 = reset ? 4'h0 : T1351;
  assign T1351 = T1353 ? T52 : T1352;
  assign T1352 = io_resetCounts ? 4'h0 : counts_216;
  assign T1353 = T10320 & T1354;
  assign T1354 = T76[8'hd8:8'hd8];
  assign T10562 = reset ? 4'h0 : T1355;
  assign T1355 = T1357 ? T52 : T1356;
  assign T1356 = io_resetCounts ? 4'h0 : counts_217;
  assign T1357 = T10320 & T1358;
  assign T1358 = T76[8'hd9:8'hd9];
  assign T1359 = T68[1'h0:1'h0];
  assign T1360 = T1369 ? counts_219 : counts_218;
  assign T10563 = reset ? 4'h0 : T1361;
  assign T1361 = T1363 ? T52 : T1362;
  assign T1362 = io_resetCounts ? 4'h0 : counts_218;
  assign T1363 = T10320 & T1364;
  assign T1364 = T76[8'hda:8'hda];
  assign T10564 = reset ? 4'h0 : T1365;
  assign T1365 = T1367 ? T52 : T1366;
  assign T1366 = io_resetCounts ? 4'h0 : counts_219;
  assign T1367 = T10320 & T1368;
  assign T1368 = T76[8'hdb:8'hdb];
  assign T1369 = T68[1'h0:1'h0];
  assign T1370 = T68[1'h1:1'h1];
  assign T1371 = T1392 ? T1382 : T1372;
  assign T1372 = T1381 ? counts_221 : counts_220;
  assign T10565 = reset ? 4'h0 : T1373;
  assign T1373 = T1375 ? T52 : T1374;
  assign T1374 = io_resetCounts ? 4'h0 : counts_220;
  assign T1375 = T10320 & T1376;
  assign T1376 = T76[8'hdc:8'hdc];
  assign T10566 = reset ? 4'h0 : T1377;
  assign T1377 = T1379 ? T52 : T1378;
  assign T1378 = io_resetCounts ? 4'h0 : counts_221;
  assign T1379 = T10320 & T1380;
  assign T1380 = T76[8'hdd:8'hdd];
  assign T1381 = T68[1'h0:1'h0];
  assign T1382 = T1391 ? counts_223 : counts_222;
  assign T10567 = reset ? 4'h0 : T1383;
  assign T1383 = T1385 ? T52 : T1384;
  assign T1384 = io_resetCounts ? 4'h0 : counts_222;
  assign T1385 = T10320 & T1386;
  assign T1386 = T76[8'hde:8'hde];
  assign T10568 = reset ? 4'h0 : T1387;
  assign T1387 = T1389 ? T52 : T1388;
  assign T1388 = io_resetCounts ? 4'h0 : counts_223;
  assign T1389 = T10320 & T1390;
  assign T1390 = T76[8'hdf:8'hdf];
  assign T1391 = T68[1'h0:1'h0];
  assign T1392 = T68[1'h1:1'h1];
  assign T1393 = T68[2'h2:2'h2];
  assign T1394 = T68[2'h3:2'h3];
  assign T1395 = T68[3'h4:3'h4];
  assign T1396 = T1585 ? T1491 : T1397;
  assign T1397 = T1490 ? T1444 : T1398;
  assign T1398 = T1443 ? T1421 : T1399;
  assign T1399 = T1420 ? T1410 : T1400;
  assign T1400 = T1409 ? counts_225 : counts_224;
  assign T10569 = reset ? 4'h0 : T1401;
  assign T1401 = T1403 ? T52 : T1402;
  assign T1402 = io_resetCounts ? 4'h0 : counts_224;
  assign T1403 = T10320 & T1404;
  assign T1404 = T76[8'he0:8'he0];
  assign T10570 = reset ? 4'h0 : T1405;
  assign T1405 = T1407 ? T52 : T1406;
  assign T1406 = io_resetCounts ? 4'h0 : counts_225;
  assign T1407 = T10320 & T1408;
  assign T1408 = T76[8'he1:8'he1];
  assign T1409 = T68[1'h0:1'h0];
  assign T1410 = T1419 ? counts_227 : counts_226;
  assign T10571 = reset ? 4'h0 : T1411;
  assign T1411 = T1413 ? T52 : T1412;
  assign T1412 = io_resetCounts ? 4'h0 : counts_226;
  assign T1413 = T10320 & T1414;
  assign T1414 = T76[8'he2:8'he2];
  assign T10572 = reset ? 4'h0 : T1415;
  assign T1415 = T1417 ? T52 : T1416;
  assign T1416 = io_resetCounts ? 4'h0 : counts_227;
  assign T1417 = T10320 & T1418;
  assign T1418 = T76[8'he3:8'he3];
  assign T1419 = T68[1'h0:1'h0];
  assign T1420 = T68[1'h1:1'h1];
  assign T1421 = T1442 ? T1432 : T1422;
  assign T1422 = T1431 ? counts_229 : counts_228;
  assign T10573 = reset ? 4'h0 : T1423;
  assign T1423 = T1425 ? T52 : T1424;
  assign T1424 = io_resetCounts ? 4'h0 : counts_228;
  assign T1425 = T10320 & T1426;
  assign T1426 = T76[8'he4:8'he4];
  assign T10574 = reset ? 4'h0 : T1427;
  assign T1427 = T1429 ? T52 : T1428;
  assign T1428 = io_resetCounts ? 4'h0 : counts_229;
  assign T1429 = T10320 & T1430;
  assign T1430 = T76[8'he5:8'he5];
  assign T1431 = T68[1'h0:1'h0];
  assign T1432 = T1441 ? counts_231 : counts_230;
  assign T10575 = reset ? 4'h0 : T1433;
  assign T1433 = T1435 ? T52 : T1434;
  assign T1434 = io_resetCounts ? 4'h0 : counts_230;
  assign T1435 = T10320 & T1436;
  assign T1436 = T76[8'he6:8'he6];
  assign T10576 = reset ? 4'h0 : T1437;
  assign T1437 = T1439 ? T52 : T1438;
  assign T1438 = io_resetCounts ? 4'h0 : counts_231;
  assign T1439 = T10320 & T1440;
  assign T1440 = T76[8'he7:8'he7];
  assign T1441 = T68[1'h0:1'h0];
  assign T1442 = T68[1'h1:1'h1];
  assign T1443 = T68[2'h2:2'h2];
  assign T1444 = T1489 ? T1467 : T1445;
  assign T1445 = T1466 ? T1456 : T1446;
  assign T1446 = T1455 ? counts_233 : counts_232;
  assign T10577 = reset ? 4'h0 : T1447;
  assign T1447 = T1449 ? T52 : T1448;
  assign T1448 = io_resetCounts ? 4'h0 : counts_232;
  assign T1449 = T10320 & T1450;
  assign T1450 = T76[8'he8:8'he8];
  assign T10578 = reset ? 4'h0 : T1451;
  assign T1451 = T1453 ? T52 : T1452;
  assign T1452 = io_resetCounts ? 4'h0 : counts_233;
  assign T1453 = T10320 & T1454;
  assign T1454 = T76[8'he9:8'he9];
  assign T1455 = T68[1'h0:1'h0];
  assign T1456 = T1465 ? counts_235 : counts_234;
  assign T10579 = reset ? 4'h0 : T1457;
  assign T1457 = T1459 ? T52 : T1458;
  assign T1458 = io_resetCounts ? 4'h0 : counts_234;
  assign T1459 = T10320 & T1460;
  assign T1460 = T76[8'hea:8'hea];
  assign T10580 = reset ? 4'h0 : T1461;
  assign T1461 = T1463 ? T52 : T1462;
  assign T1462 = io_resetCounts ? 4'h0 : counts_235;
  assign T1463 = T10320 & T1464;
  assign T1464 = T76[8'heb:8'heb];
  assign T1465 = T68[1'h0:1'h0];
  assign T1466 = T68[1'h1:1'h1];
  assign T1467 = T1488 ? T1478 : T1468;
  assign T1468 = T1477 ? counts_237 : counts_236;
  assign T10581 = reset ? 4'h0 : T1469;
  assign T1469 = T1471 ? T52 : T1470;
  assign T1470 = io_resetCounts ? 4'h0 : counts_236;
  assign T1471 = T10320 & T1472;
  assign T1472 = T76[8'hec:8'hec];
  assign T10582 = reset ? 4'h0 : T1473;
  assign T1473 = T1475 ? T52 : T1474;
  assign T1474 = io_resetCounts ? 4'h0 : counts_237;
  assign T1475 = T10320 & T1476;
  assign T1476 = T76[8'hed:8'hed];
  assign T1477 = T68[1'h0:1'h0];
  assign T1478 = T1487 ? counts_239 : counts_238;
  assign T10583 = reset ? 4'h0 : T1479;
  assign T1479 = T1481 ? T52 : T1480;
  assign T1480 = io_resetCounts ? 4'h0 : counts_238;
  assign T1481 = T10320 & T1482;
  assign T1482 = T76[8'hee:8'hee];
  assign T10584 = reset ? 4'h0 : T1483;
  assign T1483 = T1485 ? T52 : T1484;
  assign T1484 = io_resetCounts ? 4'h0 : counts_239;
  assign T1485 = T10320 & T1486;
  assign T1486 = T76[8'hef:8'hef];
  assign T1487 = T68[1'h0:1'h0];
  assign T1488 = T68[1'h1:1'h1];
  assign T1489 = T68[2'h2:2'h2];
  assign T1490 = T68[2'h3:2'h3];
  assign T1491 = T1584 ? T1538 : T1492;
  assign T1492 = T1537 ? T1515 : T1493;
  assign T1493 = T1514 ? T1504 : T1494;
  assign T1494 = T1503 ? counts_241 : counts_240;
  assign T10585 = reset ? 4'h0 : T1495;
  assign T1495 = T1497 ? T52 : T1496;
  assign T1496 = io_resetCounts ? 4'h0 : counts_240;
  assign T1497 = T10320 & T1498;
  assign T1498 = T76[8'hf0:8'hf0];
  assign T10586 = reset ? 4'h0 : T1499;
  assign T1499 = T1501 ? T52 : T1500;
  assign T1500 = io_resetCounts ? 4'h0 : counts_241;
  assign T1501 = T10320 & T1502;
  assign T1502 = T76[8'hf1:8'hf1];
  assign T1503 = T68[1'h0:1'h0];
  assign T1504 = T1513 ? counts_243 : counts_242;
  assign T10587 = reset ? 4'h0 : T1505;
  assign T1505 = T1507 ? T52 : T1506;
  assign T1506 = io_resetCounts ? 4'h0 : counts_242;
  assign T1507 = T10320 & T1508;
  assign T1508 = T76[8'hf2:8'hf2];
  assign T10588 = reset ? 4'h0 : T1509;
  assign T1509 = T1511 ? T52 : T1510;
  assign T1510 = io_resetCounts ? 4'h0 : counts_243;
  assign T1511 = T10320 & T1512;
  assign T1512 = T76[8'hf3:8'hf3];
  assign T1513 = T68[1'h0:1'h0];
  assign T1514 = T68[1'h1:1'h1];
  assign T1515 = T1536 ? T1526 : T1516;
  assign T1516 = T1525 ? counts_245 : counts_244;
  assign T10589 = reset ? 4'h0 : T1517;
  assign T1517 = T1519 ? T52 : T1518;
  assign T1518 = io_resetCounts ? 4'h0 : counts_244;
  assign T1519 = T10320 & T1520;
  assign T1520 = T76[8'hf4:8'hf4];
  assign T10590 = reset ? 4'h0 : T1521;
  assign T1521 = T1523 ? T52 : T1522;
  assign T1522 = io_resetCounts ? 4'h0 : counts_245;
  assign T1523 = T10320 & T1524;
  assign T1524 = T76[8'hf5:8'hf5];
  assign T1525 = T68[1'h0:1'h0];
  assign T1526 = T1535 ? counts_247 : counts_246;
  assign T10591 = reset ? 4'h0 : T1527;
  assign T1527 = T1529 ? T52 : T1528;
  assign T1528 = io_resetCounts ? 4'h0 : counts_246;
  assign T1529 = T10320 & T1530;
  assign T1530 = T76[8'hf6:8'hf6];
  assign T10592 = reset ? 4'h0 : T1531;
  assign T1531 = T1533 ? T52 : T1532;
  assign T1532 = io_resetCounts ? 4'h0 : counts_247;
  assign T1533 = T10320 & T1534;
  assign T1534 = T76[8'hf7:8'hf7];
  assign T1535 = T68[1'h0:1'h0];
  assign T1536 = T68[1'h1:1'h1];
  assign T1537 = T68[2'h2:2'h2];
  assign T1538 = T1583 ? T1561 : T1539;
  assign T1539 = T1560 ? T1550 : T1540;
  assign T1540 = T1549 ? counts_249 : counts_248;
  assign T10593 = reset ? 4'h0 : T1541;
  assign T1541 = T1543 ? T52 : T1542;
  assign T1542 = io_resetCounts ? 4'h0 : counts_248;
  assign T1543 = T10320 & T1544;
  assign T1544 = T76[8'hf8:8'hf8];
  assign T10594 = reset ? 4'h0 : T1545;
  assign T1545 = T1547 ? T52 : T1546;
  assign T1546 = io_resetCounts ? 4'h0 : counts_249;
  assign T1547 = T10320 & T1548;
  assign T1548 = T76[8'hf9:8'hf9];
  assign T1549 = T68[1'h0:1'h0];
  assign T1550 = T1559 ? counts_251 : counts_250;
  assign T10595 = reset ? 4'h0 : T1551;
  assign T1551 = T1553 ? T52 : T1552;
  assign T1552 = io_resetCounts ? 4'h0 : counts_250;
  assign T1553 = T10320 & T1554;
  assign T1554 = T76[8'hfa:8'hfa];
  assign T10596 = reset ? 4'h0 : T1555;
  assign T1555 = T1557 ? T52 : T1556;
  assign T1556 = io_resetCounts ? 4'h0 : counts_251;
  assign T1557 = T10320 & T1558;
  assign T1558 = T76[8'hfb:8'hfb];
  assign T1559 = T68[1'h0:1'h0];
  assign T1560 = T68[1'h1:1'h1];
  assign T1561 = T1582 ? T1572 : T1562;
  assign T1562 = T1571 ? counts_253 : counts_252;
  assign T10597 = reset ? 4'h0 : T1563;
  assign T1563 = T1565 ? T52 : T1564;
  assign T1564 = io_resetCounts ? 4'h0 : counts_252;
  assign T1565 = T10320 & T1566;
  assign T1566 = T76[8'hfc:8'hfc];
  assign T10598 = reset ? 4'h0 : T1567;
  assign T1567 = T1569 ? T52 : T1568;
  assign T1568 = io_resetCounts ? 4'h0 : counts_253;
  assign T1569 = T10320 & T1570;
  assign T1570 = T76[8'hfd:8'hfd];
  assign T1571 = T68[1'h0:1'h0];
  assign T1572 = T1581 ? counts_255 : counts_254;
  assign T10599 = reset ? 4'h0 : T1573;
  assign T1573 = T1575 ? T52 : T1574;
  assign T1574 = io_resetCounts ? 4'h0 : counts_254;
  assign T1575 = T10320 & T1576;
  assign T1576 = T76[8'hfe:8'hfe];
  assign T10600 = reset ? 4'h0 : T1577;
  assign T1577 = T1579 ? T52 : T1578;
  assign T1578 = io_resetCounts ? 4'h0 : counts_255;
  assign T1579 = T10320 & T1580;
  assign T1580 = T76[8'hff:8'hff];
  assign T1581 = T68[1'h0:1'h0];
  assign T1582 = T68[1'h1:1'h1];
  assign T1583 = T68[2'h2:2'h2];
  assign T1584 = T68[2'h3:2'h3];
  assign T1585 = T68[3'h4:3'h4];
  assign T1586 = T68[3'h5:3'h5];
  assign T1587 = T68[3'h6:3'h6];
  assign T1588 = T68[3'h7:3'h7];
  assign T1589 = T3122 ? T2356 : T1590;
  assign T1590 = T2355 ? T1973 : T1591;
  assign T1591 = T1972 ? T1782 : T1592;
  assign T1592 = T1781 ? T1687 : T1593;
  assign T1593 = T1686 ? T1640 : T1594;
  assign T1594 = T1639 ? T1617 : T1595;
  assign T1595 = T1616 ? T1606 : T1596;
  assign T1596 = T1605 ? counts_257 : counts_256;
  assign T10601 = reset ? 4'h0 : T1597;
  assign T1597 = T1599 ? T52 : T1598;
  assign T1598 = io_resetCounts ? 4'h0 : counts_256;
  assign T1599 = T10320 & T1600;
  assign T1600 = T76[9'h100:9'h100];
  assign T10602 = reset ? 4'h0 : T1601;
  assign T1601 = T1603 ? T52 : T1602;
  assign T1602 = io_resetCounts ? 4'h0 : counts_257;
  assign T1603 = T10320 & T1604;
  assign T1604 = T76[9'h101:9'h101];
  assign T1605 = T68[1'h0:1'h0];
  assign T1606 = T1615 ? counts_259 : counts_258;
  assign T10603 = reset ? 4'h0 : T1607;
  assign T1607 = T1609 ? T52 : T1608;
  assign T1608 = io_resetCounts ? 4'h0 : counts_258;
  assign T1609 = T10320 & T1610;
  assign T1610 = T76[9'h102:9'h102];
  assign T10604 = reset ? 4'h0 : T1611;
  assign T1611 = T1613 ? T52 : T1612;
  assign T1612 = io_resetCounts ? 4'h0 : counts_259;
  assign T1613 = T10320 & T1614;
  assign T1614 = T76[9'h103:9'h103];
  assign T1615 = T68[1'h0:1'h0];
  assign T1616 = T68[1'h1:1'h1];
  assign T1617 = T1638 ? T1628 : T1618;
  assign T1618 = T1627 ? counts_261 : counts_260;
  assign T10605 = reset ? 4'h0 : T1619;
  assign T1619 = T1621 ? T52 : T1620;
  assign T1620 = io_resetCounts ? 4'h0 : counts_260;
  assign T1621 = T10320 & T1622;
  assign T1622 = T76[9'h104:9'h104];
  assign T10606 = reset ? 4'h0 : T1623;
  assign T1623 = T1625 ? T52 : T1624;
  assign T1624 = io_resetCounts ? 4'h0 : counts_261;
  assign T1625 = T10320 & T1626;
  assign T1626 = T76[9'h105:9'h105];
  assign T1627 = T68[1'h0:1'h0];
  assign T1628 = T1637 ? counts_263 : counts_262;
  assign T10607 = reset ? 4'h0 : T1629;
  assign T1629 = T1631 ? T52 : T1630;
  assign T1630 = io_resetCounts ? 4'h0 : counts_262;
  assign T1631 = T10320 & T1632;
  assign T1632 = T76[9'h106:9'h106];
  assign T10608 = reset ? 4'h0 : T1633;
  assign T1633 = T1635 ? T52 : T1634;
  assign T1634 = io_resetCounts ? 4'h0 : counts_263;
  assign T1635 = T10320 & T1636;
  assign T1636 = T76[9'h107:9'h107];
  assign T1637 = T68[1'h0:1'h0];
  assign T1638 = T68[1'h1:1'h1];
  assign T1639 = T68[2'h2:2'h2];
  assign T1640 = T1685 ? T1663 : T1641;
  assign T1641 = T1662 ? T1652 : T1642;
  assign T1642 = T1651 ? counts_265 : counts_264;
  assign T10609 = reset ? 4'h0 : T1643;
  assign T1643 = T1645 ? T52 : T1644;
  assign T1644 = io_resetCounts ? 4'h0 : counts_264;
  assign T1645 = T10320 & T1646;
  assign T1646 = T76[9'h108:9'h108];
  assign T10610 = reset ? 4'h0 : T1647;
  assign T1647 = T1649 ? T52 : T1648;
  assign T1648 = io_resetCounts ? 4'h0 : counts_265;
  assign T1649 = T10320 & T1650;
  assign T1650 = T76[9'h109:9'h109];
  assign T1651 = T68[1'h0:1'h0];
  assign T1652 = T1661 ? counts_267 : counts_266;
  assign T10611 = reset ? 4'h0 : T1653;
  assign T1653 = T1655 ? T52 : T1654;
  assign T1654 = io_resetCounts ? 4'h0 : counts_266;
  assign T1655 = T10320 & T1656;
  assign T1656 = T76[9'h10a:9'h10a];
  assign T10612 = reset ? 4'h0 : T1657;
  assign T1657 = T1659 ? T52 : T1658;
  assign T1658 = io_resetCounts ? 4'h0 : counts_267;
  assign T1659 = T10320 & T1660;
  assign T1660 = T76[9'h10b:9'h10b];
  assign T1661 = T68[1'h0:1'h0];
  assign T1662 = T68[1'h1:1'h1];
  assign T1663 = T1684 ? T1674 : T1664;
  assign T1664 = T1673 ? counts_269 : counts_268;
  assign T10613 = reset ? 4'h0 : T1665;
  assign T1665 = T1667 ? T52 : T1666;
  assign T1666 = io_resetCounts ? 4'h0 : counts_268;
  assign T1667 = T10320 & T1668;
  assign T1668 = T76[9'h10c:9'h10c];
  assign T10614 = reset ? 4'h0 : T1669;
  assign T1669 = T1671 ? T52 : T1670;
  assign T1670 = io_resetCounts ? 4'h0 : counts_269;
  assign T1671 = T10320 & T1672;
  assign T1672 = T76[9'h10d:9'h10d];
  assign T1673 = T68[1'h0:1'h0];
  assign T1674 = T1683 ? counts_271 : counts_270;
  assign T10615 = reset ? 4'h0 : T1675;
  assign T1675 = T1677 ? T52 : T1676;
  assign T1676 = io_resetCounts ? 4'h0 : counts_270;
  assign T1677 = T10320 & T1678;
  assign T1678 = T76[9'h10e:9'h10e];
  assign T10616 = reset ? 4'h0 : T1679;
  assign T1679 = T1681 ? T52 : T1680;
  assign T1680 = io_resetCounts ? 4'h0 : counts_271;
  assign T1681 = T10320 & T1682;
  assign T1682 = T76[9'h10f:9'h10f];
  assign T1683 = T68[1'h0:1'h0];
  assign T1684 = T68[1'h1:1'h1];
  assign T1685 = T68[2'h2:2'h2];
  assign T1686 = T68[2'h3:2'h3];
  assign T1687 = T1780 ? T1734 : T1688;
  assign T1688 = T1733 ? T1711 : T1689;
  assign T1689 = T1710 ? T1700 : T1690;
  assign T1690 = T1699 ? counts_273 : counts_272;
  assign T10617 = reset ? 4'h0 : T1691;
  assign T1691 = T1693 ? T52 : T1692;
  assign T1692 = io_resetCounts ? 4'h0 : counts_272;
  assign T1693 = T10320 & T1694;
  assign T1694 = T76[9'h110:9'h110];
  assign T10618 = reset ? 4'h0 : T1695;
  assign T1695 = T1697 ? T52 : T1696;
  assign T1696 = io_resetCounts ? 4'h0 : counts_273;
  assign T1697 = T10320 & T1698;
  assign T1698 = T76[9'h111:9'h111];
  assign T1699 = T68[1'h0:1'h0];
  assign T1700 = T1709 ? counts_275 : counts_274;
  assign T10619 = reset ? 4'h0 : T1701;
  assign T1701 = T1703 ? T52 : T1702;
  assign T1702 = io_resetCounts ? 4'h0 : counts_274;
  assign T1703 = T10320 & T1704;
  assign T1704 = T76[9'h112:9'h112];
  assign T10620 = reset ? 4'h0 : T1705;
  assign T1705 = T1707 ? T52 : T1706;
  assign T1706 = io_resetCounts ? 4'h0 : counts_275;
  assign T1707 = T10320 & T1708;
  assign T1708 = T76[9'h113:9'h113];
  assign T1709 = T68[1'h0:1'h0];
  assign T1710 = T68[1'h1:1'h1];
  assign T1711 = T1732 ? T1722 : T1712;
  assign T1712 = T1721 ? counts_277 : counts_276;
  assign T10621 = reset ? 4'h0 : T1713;
  assign T1713 = T1715 ? T52 : T1714;
  assign T1714 = io_resetCounts ? 4'h0 : counts_276;
  assign T1715 = T10320 & T1716;
  assign T1716 = T76[9'h114:9'h114];
  assign T10622 = reset ? 4'h0 : T1717;
  assign T1717 = T1719 ? T52 : T1718;
  assign T1718 = io_resetCounts ? 4'h0 : counts_277;
  assign T1719 = T10320 & T1720;
  assign T1720 = T76[9'h115:9'h115];
  assign T1721 = T68[1'h0:1'h0];
  assign T1722 = T1731 ? counts_279 : counts_278;
  assign T10623 = reset ? 4'h0 : T1723;
  assign T1723 = T1725 ? T52 : T1724;
  assign T1724 = io_resetCounts ? 4'h0 : counts_278;
  assign T1725 = T10320 & T1726;
  assign T1726 = T76[9'h116:9'h116];
  assign T10624 = reset ? 4'h0 : T1727;
  assign T1727 = T1729 ? T52 : T1728;
  assign T1728 = io_resetCounts ? 4'h0 : counts_279;
  assign T1729 = T10320 & T1730;
  assign T1730 = T76[9'h117:9'h117];
  assign T1731 = T68[1'h0:1'h0];
  assign T1732 = T68[1'h1:1'h1];
  assign T1733 = T68[2'h2:2'h2];
  assign T1734 = T1779 ? T1757 : T1735;
  assign T1735 = T1756 ? T1746 : T1736;
  assign T1736 = T1745 ? counts_281 : counts_280;
  assign T10625 = reset ? 4'h0 : T1737;
  assign T1737 = T1739 ? T52 : T1738;
  assign T1738 = io_resetCounts ? 4'h0 : counts_280;
  assign T1739 = T10320 & T1740;
  assign T1740 = T76[9'h118:9'h118];
  assign T10626 = reset ? 4'h0 : T1741;
  assign T1741 = T1743 ? T52 : T1742;
  assign T1742 = io_resetCounts ? 4'h0 : counts_281;
  assign T1743 = T10320 & T1744;
  assign T1744 = T76[9'h119:9'h119];
  assign T1745 = T68[1'h0:1'h0];
  assign T1746 = T1755 ? counts_283 : counts_282;
  assign T10627 = reset ? 4'h0 : T1747;
  assign T1747 = T1749 ? T52 : T1748;
  assign T1748 = io_resetCounts ? 4'h0 : counts_282;
  assign T1749 = T10320 & T1750;
  assign T1750 = T76[9'h11a:9'h11a];
  assign T10628 = reset ? 4'h0 : T1751;
  assign T1751 = T1753 ? T52 : T1752;
  assign T1752 = io_resetCounts ? 4'h0 : counts_283;
  assign T1753 = T10320 & T1754;
  assign T1754 = T76[9'h11b:9'h11b];
  assign T1755 = T68[1'h0:1'h0];
  assign T1756 = T68[1'h1:1'h1];
  assign T1757 = T1778 ? T1768 : T1758;
  assign T1758 = T1767 ? counts_285 : counts_284;
  assign T10629 = reset ? 4'h0 : T1759;
  assign T1759 = T1761 ? T52 : T1760;
  assign T1760 = io_resetCounts ? 4'h0 : counts_284;
  assign T1761 = T10320 & T1762;
  assign T1762 = T76[9'h11c:9'h11c];
  assign T10630 = reset ? 4'h0 : T1763;
  assign T1763 = T1765 ? T52 : T1764;
  assign T1764 = io_resetCounts ? 4'h0 : counts_285;
  assign T1765 = T10320 & T1766;
  assign T1766 = T76[9'h11d:9'h11d];
  assign T1767 = T68[1'h0:1'h0];
  assign T1768 = T1777 ? counts_287 : counts_286;
  assign T10631 = reset ? 4'h0 : T1769;
  assign T1769 = T1771 ? T52 : T1770;
  assign T1770 = io_resetCounts ? 4'h0 : counts_286;
  assign T1771 = T10320 & T1772;
  assign T1772 = T76[9'h11e:9'h11e];
  assign T10632 = reset ? 4'h0 : T1773;
  assign T1773 = T1775 ? T52 : T1774;
  assign T1774 = io_resetCounts ? 4'h0 : counts_287;
  assign T1775 = T10320 & T1776;
  assign T1776 = T76[9'h11f:9'h11f];
  assign T1777 = T68[1'h0:1'h0];
  assign T1778 = T68[1'h1:1'h1];
  assign T1779 = T68[2'h2:2'h2];
  assign T1780 = T68[2'h3:2'h3];
  assign T1781 = T68[3'h4:3'h4];
  assign T1782 = T1971 ? T1877 : T1783;
  assign T1783 = T1876 ? T1830 : T1784;
  assign T1784 = T1829 ? T1807 : T1785;
  assign T1785 = T1806 ? T1796 : T1786;
  assign T1786 = T1795 ? counts_289 : counts_288;
  assign T10633 = reset ? 4'h0 : T1787;
  assign T1787 = T1789 ? T52 : T1788;
  assign T1788 = io_resetCounts ? 4'h0 : counts_288;
  assign T1789 = T10320 & T1790;
  assign T1790 = T76[9'h120:9'h120];
  assign T10634 = reset ? 4'h0 : T1791;
  assign T1791 = T1793 ? T52 : T1792;
  assign T1792 = io_resetCounts ? 4'h0 : counts_289;
  assign T1793 = T10320 & T1794;
  assign T1794 = T76[9'h121:9'h121];
  assign T1795 = T68[1'h0:1'h0];
  assign T1796 = T1805 ? counts_291 : counts_290;
  assign T10635 = reset ? 4'h0 : T1797;
  assign T1797 = T1799 ? T52 : T1798;
  assign T1798 = io_resetCounts ? 4'h0 : counts_290;
  assign T1799 = T10320 & T1800;
  assign T1800 = T76[9'h122:9'h122];
  assign T10636 = reset ? 4'h0 : T1801;
  assign T1801 = T1803 ? T52 : T1802;
  assign T1802 = io_resetCounts ? 4'h0 : counts_291;
  assign T1803 = T10320 & T1804;
  assign T1804 = T76[9'h123:9'h123];
  assign T1805 = T68[1'h0:1'h0];
  assign T1806 = T68[1'h1:1'h1];
  assign T1807 = T1828 ? T1818 : T1808;
  assign T1808 = T1817 ? counts_293 : counts_292;
  assign T10637 = reset ? 4'h0 : T1809;
  assign T1809 = T1811 ? T52 : T1810;
  assign T1810 = io_resetCounts ? 4'h0 : counts_292;
  assign T1811 = T10320 & T1812;
  assign T1812 = T76[9'h124:9'h124];
  assign T10638 = reset ? 4'h0 : T1813;
  assign T1813 = T1815 ? T52 : T1814;
  assign T1814 = io_resetCounts ? 4'h0 : counts_293;
  assign T1815 = T10320 & T1816;
  assign T1816 = T76[9'h125:9'h125];
  assign T1817 = T68[1'h0:1'h0];
  assign T1818 = T1827 ? counts_295 : counts_294;
  assign T10639 = reset ? 4'h0 : T1819;
  assign T1819 = T1821 ? T52 : T1820;
  assign T1820 = io_resetCounts ? 4'h0 : counts_294;
  assign T1821 = T10320 & T1822;
  assign T1822 = T76[9'h126:9'h126];
  assign T10640 = reset ? 4'h0 : T1823;
  assign T1823 = T1825 ? T52 : T1824;
  assign T1824 = io_resetCounts ? 4'h0 : counts_295;
  assign T1825 = T10320 & T1826;
  assign T1826 = T76[9'h127:9'h127];
  assign T1827 = T68[1'h0:1'h0];
  assign T1828 = T68[1'h1:1'h1];
  assign T1829 = T68[2'h2:2'h2];
  assign T1830 = T1875 ? T1853 : T1831;
  assign T1831 = T1852 ? T1842 : T1832;
  assign T1832 = T1841 ? counts_297 : counts_296;
  assign T10641 = reset ? 4'h0 : T1833;
  assign T1833 = T1835 ? T52 : T1834;
  assign T1834 = io_resetCounts ? 4'h0 : counts_296;
  assign T1835 = T10320 & T1836;
  assign T1836 = T76[9'h128:9'h128];
  assign T10642 = reset ? 4'h0 : T1837;
  assign T1837 = T1839 ? T52 : T1838;
  assign T1838 = io_resetCounts ? 4'h0 : counts_297;
  assign T1839 = T10320 & T1840;
  assign T1840 = T76[9'h129:9'h129];
  assign T1841 = T68[1'h0:1'h0];
  assign T1842 = T1851 ? counts_299 : counts_298;
  assign T10643 = reset ? 4'h0 : T1843;
  assign T1843 = T1845 ? T52 : T1844;
  assign T1844 = io_resetCounts ? 4'h0 : counts_298;
  assign T1845 = T10320 & T1846;
  assign T1846 = T76[9'h12a:9'h12a];
  assign T10644 = reset ? 4'h0 : T1847;
  assign T1847 = T1849 ? T52 : T1848;
  assign T1848 = io_resetCounts ? 4'h0 : counts_299;
  assign T1849 = T10320 & T1850;
  assign T1850 = T76[9'h12b:9'h12b];
  assign T1851 = T68[1'h0:1'h0];
  assign T1852 = T68[1'h1:1'h1];
  assign T1853 = T1874 ? T1864 : T1854;
  assign T1854 = T1863 ? counts_301 : counts_300;
  assign T10645 = reset ? 4'h0 : T1855;
  assign T1855 = T1857 ? T52 : T1856;
  assign T1856 = io_resetCounts ? 4'h0 : counts_300;
  assign T1857 = T10320 & T1858;
  assign T1858 = T76[9'h12c:9'h12c];
  assign T10646 = reset ? 4'h0 : T1859;
  assign T1859 = T1861 ? T52 : T1860;
  assign T1860 = io_resetCounts ? 4'h0 : counts_301;
  assign T1861 = T10320 & T1862;
  assign T1862 = T76[9'h12d:9'h12d];
  assign T1863 = T68[1'h0:1'h0];
  assign T1864 = T1873 ? counts_303 : counts_302;
  assign T10647 = reset ? 4'h0 : T1865;
  assign T1865 = T1867 ? T52 : T1866;
  assign T1866 = io_resetCounts ? 4'h0 : counts_302;
  assign T1867 = T10320 & T1868;
  assign T1868 = T76[9'h12e:9'h12e];
  assign T10648 = reset ? 4'h0 : T1869;
  assign T1869 = T1871 ? T52 : T1870;
  assign T1870 = io_resetCounts ? 4'h0 : counts_303;
  assign T1871 = T10320 & T1872;
  assign T1872 = T76[9'h12f:9'h12f];
  assign T1873 = T68[1'h0:1'h0];
  assign T1874 = T68[1'h1:1'h1];
  assign T1875 = T68[2'h2:2'h2];
  assign T1876 = T68[2'h3:2'h3];
  assign T1877 = T1970 ? T1924 : T1878;
  assign T1878 = T1923 ? T1901 : T1879;
  assign T1879 = T1900 ? T1890 : T1880;
  assign T1880 = T1889 ? counts_305 : counts_304;
  assign T10649 = reset ? 4'h0 : T1881;
  assign T1881 = T1883 ? T52 : T1882;
  assign T1882 = io_resetCounts ? 4'h0 : counts_304;
  assign T1883 = T10320 & T1884;
  assign T1884 = T76[9'h130:9'h130];
  assign T10650 = reset ? 4'h0 : T1885;
  assign T1885 = T1887 ? T52 : T1886;
  assign T1886 = io_resetCounts ? 4'h0 : counts_305;
  assign T1887 = T10320 & T1888;
  assign T1888 = T76[9'h131:9'h131];
  assign T1889 = T68[1'h0:1'h0];
  assign T1890 = T1899 ? counts_307 : counts_306;
  assign T10651 = reset ? 4'h0 : T1891;
  assign T1891 = T1893 ? T52 : T1892;
  assign T1892 = io_resetCounts ? 4'h0 : counts_306;
  assign T1893 = T10320 & T1894;
  assign T1894 = T76[9'h132:9'h132];
  assign T10652 = reset ? 4'h0 : T1895;
  assign T1895 = T1897 ? T52 : T1896;
  assign T1896 = io_resetCounts ? 4'h0 : counts_307;
  assign T1897 = T10320 & T1898;
  assign T1898 = T76[9'h133:9'h133];
  assign T1899 = T68[1'h0:1'h0];
  assign T1900 = T68[1'h1:1'h1];
  assign T1901 = T1922 ? T1912 : T1902;
  assign T1902 = T1911 ? counts_309 : counts_308;
  assign T10653 = reset ? 4'h0 : T1903;
  assign T1903 = T1905 ? T52 : T1904;
  assign T1904 = io_resetCounts ? 4'h0 : counts_308;
  assign T1905 = T10320 & T1906;
  assign T1906 = T76[9'h134:9'h134];
  assign T10654 = reset ? 4'h0 : T1907;
  assign T1907 = T1909 ? T52 : T1908;
  assign T1908 = io_resetCounts ? 4'h0 : counts_309;
  assign T1909 = T10320 & T1910;
  assign T1910 = T76[9'h135:9'h135];
  assign T1911 = T68[1'h0:1'h0];
  assign T1912 = T1921 ? counts_311 : counts_310;
  assign T10655 = reset ? 4'h0 : T1913;
  assign T1913 = T1915 ? T52 : T1914;
  assign T1914 = io_resetCounts ? 4'h0 : counts_310;
  assign T1915 = T10320 & T1916;
  assign T1916 = T76[9'h136:9'h136];
  assign T10656 = reset ? 4'h0 : T1917;
  assign T1917 = T1919 ? T52 : T1918;
  assign T1918 = io_resetCounts ? 4'h0 : counts_311;
  assign T1919 = T10320 & T1920;
  assign T1920 = T76[9'h137:9'h137];
  assign T1921 = T68[1'h0:1'h0];
  assign T1922 = T68[1'h1:1'h1];
  assign T1923 = T68[2'h2:2'h2];
  assign T1924 = T1969 ? T1947 : T1925;
  assign T1925 = T1946 ? T1936 : T1926;
  assign T1926 = T1935 ? counts_313 : counts_312;
  assign T10657 = reset ? 4'h0 : T1927;
  assign T1927 = T1929 ? T52 : T1928;
  assign T1928 = io_resetCounts ? 4'h0 : counts_312;
  assign T1929 = T10320 & T1930;
  assign T1930 = T76[9'h138:9'h138];
  assign T10658 = reset ? 4'h0 : T1931;
  assign T1931 = T1933 ? T52 : T1932;
  assign T1932 = io_resetCounts ? 4'h0 : counts_313;
  assign T1933 = T10320 & T1934;
  assign T1934 = T76[9'h139:9'h139];
  assign T1935 = T68[1'h0:1'h0];
  assign T1936 = T1945 ? counts_315 : counts_314;
  assign T10659 = reset ? 4'h0 : T1937;
  assign T1937 = T1939 ? T52 : T1938;
  assign T1938 = io_resetCounts ? 4'h0 : counts_314;
  assign T1939 = T10320 & T1940;
  assign T1940 = T76[9'h13a:9'h13a];
  assign T10660 = reset ? 4'h0 : T1941;
  assign T1941 = T1943 ? T52 : T1942;
  assign T1942 = io_resetCounts ? 4'h0 : counts_315;
  assign T1943 = T10320 & T1944;
  assign T1944 = T76[9'h13b:9'h13b];
  assign T1945 = T68[1'h0:1'h0];
  assign T1946 = T68[1'h1:1'h1];
  assign T1947 = T1968 ? T1958 : T1948;
  assign T1948 = T1957 ? counts_317 : counts_316;
  assign T10661 = reset ? 4'h0 : T1949;
  assign T1949 = T1951 ? T52 : T1950;
  assign T1950 = io_resetCounts ? 4'h0 : counts_316;
  assign T1951 = T10320 & T1952;
  assign T1952 = T76[9'h13c:9'h13c];
  assign T10662 = reset ? 4'h0 : T1953;
  assign T1953 = T1955 ? T52 : T1954;
  assign T1954 = io_resetCounts ? 4'h0 : counts_317;
  assign T1955 = T10320 & T1956;
  assign T1956 = T76[9'h13d:9'h13d];
  assign T1957 = T68[1'h0:1'h0];
  assign T1958 = T1967 ? counts_319 : counts_318;
  assign T10663 = reset ? 4'h0 : T1959;
  assign T1959 = T1961 ? T52 : T1960;
  assign T1960 = io_resetCounts ? 4'h0 : counts_318;
  assign T1961 = T10320 & T1962;
  assign T1962 = T76[9'h13e:9'h13e];
  assign T10664 = reset ? 4'h0 : T1963;
  assign T1963 = T1965 ? T52 : T1964;
  assign T1964 = io_resetCounts ? 4'h0 : counts_319;
  assign T1965 = T10320 & T1966;
  assign T1966 = T76[9'h13f:9'h13f];
  assign T1967 = T68[1'h0:1'h0];
  assign T1968 = T68[1'h1:1'h1];
  assign T1969 = T68[2'h2:2'h2];
  assign T1970 = T68[2'h3:2'h3];
  assign T1971 = T68[3'h4:3'h4];
  assign T1972 = T68[3'h5:3'h5];
  assign T1973 = T2354 ? T2164 : T1974;
  assign T1974 = T2163 ? T2069 : T1975;
  assign T1975 = T2068 ? T2022 : T1976;
  assign T1976 = T2021 ? T1999 : T1977;
  assign T1977 = T1998 ? T1988 : T1978;
  assign T1978 = T1987 ? counts_321 : counts_320;
  assign T10665 = reset ? 4'h0 : T1979;
  assign T1979 = T1981 ? T52 : T1980;
  assign T1980 = io_resetCounts ? 4'h0 : counts_320;
  assign T1981 = T10320 & T1982;
  assign T1982 = T76[9'h140:9'h140];
  assign T10666 = reset ? 4'h0 : T1983;
  assign T1983 = T1985 ? T52 : T1984;
  assign T1984 = io_resetCounts ? 4'h0 : counts_321;
  assign T1985 = T10320 & T1986;
  assign T1986 = T76[9'h141:9'h141];
  assign T1987 = T68[1'h0:1'h0];
  assign T1988 = T1997 ? counts_323 : counts_322;
  assign T10667 = reset ? 4'h0 : T1989;
  assign T1989 = T1991 ? T52 : T1990;
  assign T1990 = io_resetCounts ? 4'h0 : counts_322;
  assign T1991 = T10320 & T1992;
  assign T1992 = T76[9'h142:9'h142];
  assign T10668 = reset ? 4'h0 : T1993;
  assign T1993 = T1995 ? T52 : T1994;
  assign T1994 = io_resetCounts ? 4'h0 : counts_323;
  assign T1995 = T10320 & T1996;
  assign T1996 = T76[9'h143:9'h143];
  assign T1997 = T68[1'h0:1'h0];
  assign T1998 = T68[1'h1:1'h1];
  assign T1999 = T2020 ? T2010 : T2000;
  assign T2000 = T2009 ? counts_325 : counts_324;
  assign T10669 = reset ? 4'h0 : T2001;
  assign T2001 = T2003 ? T52 : T2002;
  assign T2002 = io_resetCounts ? 4'h0 : counts_324;
  assign T2003 = T10320 & T2004;
  assign T2004 = T76[9'h144:9'h144];
  assign T10670 = reset ? 4'h0 : T2005;
  assign T2005 = T2007 ? T52 : T2006;
  assign T2006 = io_resetCounts ? 4'h0 : counts_325;
  assign T2007 = T10320 & T2008;
  assign T2008 = T76[9'h145:9'h145];
  assign T2009 = T68[1'h0:1'h0];
  assign T2010 = T2019 ? counts_327 : counts_326;
  assign T10671 = reset ? 4'h0 : T2011;
  assign T2011 = T2013 ? T52 : T2012;
  assign T2012 = io_resetCounts ? 4'h0 : counts_326;
  assign T2013 = T10320 & T2014;
  assign T2014 = T76[9'h146:9'h146];
  assign T10672 = reset ? 4'h0 : T2015;
  assign T2015 = T2017 ? T52 : T2016;
  assign T2016 = io_resetCounts ? 4'h0 : counts_327;
  assign T2017 = T10320 & T2018;
  assign T2018 = T76[9'h147:9'h147];
  assign T2019 = T68[1'h0:1'h0];
  assign T2020 = T68[1'h1:1'h1];
  assign T2021 = T68[2'h2:2'h2];
  assign T2022 = T2067 ? T2045 : T2023;
  assign T2023 = T2044 ? T2034 : T2024;
  assign T2024 = T2033 ? counts_329 : counts_328;
  assign T10673 = reset ? 4'h0 : T2025;
  assign T2025 = T2027 ? T52 : T2026;
  assign T2026 = io_resetCounts ? 4'h0 : counts_328;
  assign T2027 = T10320 & T2028;
  assign T2028 = T76[9'h148:9'h148];
  assign T10674 = reset ? 4'h0 : T2029;
  assign T2029 = T2031 ? T52 : T2030;
  assign T2030 = io_resetCounts ? 4'h0 : counts_329;
  assign T2031 = T10320 & T2032;
  assign T2032 = T76[9'h149:9'h149];
  assign T2033 = T68[1'h0:1'h0];
  assign T2034 = T2043 ? counts_331 : counts_330;
  assign T10675 = reset ? 4'h0 : T2035;
  assign T2035 = T2037 ? T52 : T2036;
  assign T2036 = io_resetCounts ? 4'h0 : counts_330;
  assign T2037 = T10320 & T2038;
  assign T2038 = T76[9'h14a:9'h14a];
  assign T10676 = reset ? 4'h0 : T2039;
  assign T2039 = T2041 ? T52 : T2040;
  assign T2040 = io_resetCounts ? 4'h0 : counts_331;
  assign T2041 = T10320 & T2042;
  assign T2042 = T76[9'h14b:9'h14b];
  assign T2043 = T68[1'h0:1'h0];
  assign T2044 = T68[1'h1:1'h1];
  assign T2045 = T2066 ? T2056 : T2046;
  assign T2046 = T2055 ? counts_333 : counts_332;
  assign T10677 = reset ? 4'h0 : T2047;
  assign T2047 = T2049 ? T52 : T2048;
  assign T2048 = io_resetCounts ? 4'h0 : counts_332;
  assign T2049 = T10320 & T2050;
  assign T2050 = T76[9'h14c:9'h14c];
  assign T10678 = reset ? 4'h0 : T2051;
  assign T2051 = T2053 ? T52 : T2052;
  assign T2052 = io_resetCounts ? 4'h0 : counts_333;
  assign T2053 = T10320 & T2054;
  assign T2054 = T76[9'h14d:9'h14d];
  assign T2055 = T68[1'h0:1'h0];
  assign T2056 = T2065 ? counts_335 : counts_334;
  assign T10679 = reset ? 4'h0 : T2057;
  assign T2057 = T2059 ? T52 : T2058;
  assign T2058 = io_resetCounts ? 4'h0 : counts_334;
  assign T2059 = T10320 & T2060;
  assign T2060 = T76[9'h14e:9'h14e];
  assign T10680 = reset ? 4'h0 : T2061;
  assign T2061 = T2063 ? T52 : T2062;
  assign T2062 = io_resetCounts ? 4'h0 : counts_335;
  assign T2063 = T10320 & T2064;
  assign T2064 = T76[9'h14f:9'h14f];
  assign T2065 = T68[1'h0:1'h0];
  assign T2066 = T68[1'h1:1'h1];
  assign T2067 = T68[2'h2:2'h2];
  assign T2068 = T68[2'h3:2'h3];
  assign T2069 = T2162 ? T2116 : T2070;
  assign T2070 = T2115 ? T2093 : T2071;
  assign T2071 = T2092 ? T2082 : T2072;
  assign T2072 = T2081 ? counts_337 : counts_336;
  assign T10681 = reset ? 4'h0 : T2073;
  assign T2073 = T2075 ? T52 : T2074;
  assign T2074 = io_resetCounts ? 4'h0 : counts_336;
  assign T2075 = T10320 & T2076;
  assign T2076 = T76[9'h150:9'h150];
  assign T10682 = reset ? 4'h0 : T2077;
  assign T2077 = T2079 ? T52 : T2078;
  assign T2078 = io_resetCounts ? 4'h0 : counts_337;
  assign T2079 = T10320 & T2080;
  assign T2080 = T76[9'h151:9'h151];
  assign T2081 = T68[1'h0:1'h0];
  assign T2082 = T2091 ? counts_339 : counts_338;
  assign T10683 = reset ? 4'h0 : T2083;
  assign T2083 = T2085 ? T52 : T2084;
  assign T2084 = io_resetCounts ? 4'h0 : counts_338;
  assign T2085 = T10320 & T2086;
  assign T2086 = T76[9'h152:9'h152];
  assign T10684 = reset ? 4'h0 : T2087;
  assign T2087 = T2089 ? T52 : T2088;
  assign T2088 = io_resetCounts ? 4'h0 : counts_339;
  assign T2089 = T10320 & T2090;
  assign T2090 = T76[9'h153:9'h153];
  assign T2091 = T68[1'h0:1'h0];
  assign T2092 = T68[1'h1:1'h1];
  assign T2093 = T2114 ? T2104 : T2094;
  assign T2094 = T2103 ? counts_341 : counts_340;
  assign T10685 = reset ? 4'h0 : T2095;
  assign T2095 = T2097 ? T52 : T2096;
  assign T2096 = io_resetCounts ? 4'h0 : counts_340;
  assign T2097 = T10320 & T2098;
  assign T2098 = T76[9'h154:9'h154];
  assign T10686 = reset ? 4'h0 : T2099;
  assign T2099 = T2101 ? T52 : T2100;
  assign T2100 = io_resetCounts ? 4'h0 : counts_341;
  assign T2101 = T10320 & T2102;
  assign T2102 = T76[9'h155:9'h155];
  assign T2103 = T68[1'h0:1'h0];
  assign T2104 = T2113 ? counts_343 : counts_342;
  assign T10687 = reset ? 4'h0 : T2105;
  assign T2105 = T2107 ? T52 : T2106;
  assign T2106 = io_resetCounts ? 4'h0 : counts_342;
  assign T2107 = T10320 & T2108;
  assign T2108 = T76[9'h156:9'h156];
  assign T10688 = reset ? 4'h0 : T2109;
  assign T2109 = T2111 ? T52 : T2110;
  assign T2110 = io_resetCounts ? 4'h0 : counts_343;
  assign T2111 = T10320 & T2112;
  assign T2112 = T76[9'h157:9'h157];
  assign T2113 = T68[1'h0:1'h0];
  assign T2114 = T68[1'h1:1'h1];
  assign T2115 = T68[2'h2:2'h2];
  assign T2116 = T2161 ? T2139 : T2117;
  assign T2117 = T2138 ? T2128 : T2118;
  assign T2118 = T2127 ? counts_345 : counts_344;
  assign T10689 = reset ? 4'h0 : T2119;
  assign T2119 = T2121 ? T52 : T2120;
  assign T2120 = io_resetCounts ? 4'h0 : counts_344;
  assign T2121 = T10320 & T2122;
  assign T2122 = T76[9'h158:9'h158];
  assign T10690 = reset ? 4'h0 : T2123;
  assign T2123 = T2125 ? T52 : T2124;
  assign T2124 = io_resetCounts ? 4'h0 : counts_345;
  assign T2125 = T10320 & T2126;
  assign T2126 = T76[9'h159:9'h159];
  assign T2127 = T68[1'h0:1'h0];
  assign T2128 = T2137 ? counts_347 : counts_346;
  assign T10691 = reset ? 4'h0 : T2129;
  assign T2129 = T2131 ? T52 : T2130;
  assign T2130 = io_resetCounts ? 4'h0 : counts_346;
  assign T2131 = T10320 & T2132;
  assign T2132 = T76[9'h15a:9'h15a];
  assign T10692 = reset ? 4'h0 : T2133;
  assign T2133 = T2135 ? T52 : T2134;
  assign T2134 = io_resetCounts ? 4'h0 : counts_347;
  assign T2135 = T10320 & T2136;
  assign T2136 = T76[9'h15b:9'h15b];
  assign T2137 = T68[1'h0:1'h0];
  assign T2138 = T68[1'h1:1'h1];
  assign T2139 = T2160 ? T2150 : T2140;
  assign T2140 = T2149 ? counts_349 : counts_348;
  assign T10693 = reset ? 4'h0 : T2141;
  assign T2141 = T2143 ? T52 : T2142;
  assign T2142 = io_resetCounts ? 4'h0 : counts_348;
  assign T2143 = T10320 & T2144;
  assign T2144 = T76[9'h15c:9'h15c];
  assign T10694 = reset ? 4'h0 : T2145;
  assign T2145 = T2147 ? T52 : T2146;
  assign T2146 = io_resetCounts ? 4'h0 : counts_349;
  assign T2147 = T10320 & T2148;
  assign T2148 = T76[9'h15d:9'h15d];
  assign T2149 = T68[1'h0:1'h0];
  assign T2150 = T2159 ? counts_351 : counts_350;
  assign T10695 = reset ? 4'h0 : T2151;
  assign T2151 = T2153 ? T52 : T2152;
  assign T2152 = io_resetCounts ? 4'h0 : counts_350;
  assign T2153 = T10320 & T2154;
  assign T2154 = T76[9'h15e:9'h15e];
  assign T10696 = reset ? 4'h0 : T2155;
  assign T2155 = T2157 ? T52 : T2156;
  assign T2156 = io_resetCounts ? 4'h0 : counts_351;
  assign T2157 = T10320 & T2158;
  assign T2158 = T76[9'h15f:9'h15f];
  assign T2159 = T68[1'h0:1'h0];
  assign T2160 = T68[1'h1:1'h1];
  assign T2161 = T68[2'h2:2'h2];
  assign T2162 = T68[2'h3:2'h3];
  assign T2163 = T68[3'h4:3'h4];
  assign T2164 = T2353 ? T2259 : T2165;
  assign T2165 = T2258 ? T2212 : T2166;
  assign T2166 = T2211 ? T2189 : T2167;
  assign T2167 = T2188 ? T2178 : T2168;
  assign T2168 = T2177 ? counts_353 : counts_352;
  assign T10697 = reset ? 4'h0 : T2169;
  assign T2169 = T2171 ? T52 : T2170;
  assign T2170 = io_resetCounts ? 4'h0 : counts_352;
  assign T2171 = T10320 & T2172;
  assign T2172 = T76[9'h160:9'h160];
  assign T10698 = reset ? 4'h0 : T2173;
  assign T2173 = T2175 ? T52 : T2174;
  assign T2174 = io_resetCounts ? 4'h0 : counts_353;
  assign T2175 = T10320 & T2176;
  assign T2176 = T76[9'h161:9'h161];
  assign T2177 = T68[1'h0:1'h0];
  assign T2178 = T2187 ? counts_355 : counts_354;
  assign T10699 = reset ? 4'h0 : T2179;
  assign T2179 = T2181 ? T52 : T2180;
  assign T2180 = io_resetCounts ? 4'h0 : counts_354;
  assign T2181 = T10320 & T2182;
  assign T2182 = T76[9'h162:9'h162];
  assign T10700 = reset ? 4'h0 : T2183;
  assign T2183 = T2185 ? T52 : T2184;
  assign T2184 = io_resetCounts ? 4'h0 : counts_355;
  assign T2185 = T10320 & T2186;
  assign T2186 = T76[9'h163:9'h163];
  assign T2187 = T68[1'h0:1'h0];
  assign T2188 = T68[1'h1:1'h1];
  assign T2189 = T2210 ? T2200 : T2190;
  assign T2190 = T2199 ? counts_357 : counts_356;
  assign T10701 = reset ? 4'h0 : T2191;
  assign T2191 = T2193 ? T52 : T2192;
  assign T2192 = io_resetCounts ? 4'h0 : counts_356;
  assign T2193 = T10320 & T2194;
  assign T2194 = T76[9'h164:9'h164];
  assign T10702 = reset ? 4'h0 : T2195;
  assign T2195 = T2197 ? T52 : T2196;
  assign T2196 = io_resetCounts ? 4'h0 : counts_357;
  assign T2197 = T10320 & T2198;
  assign T2198 = T76[9'h165:9'h165];
  assign T2199 = T68[1'h0:1'h0];
  assign T2200 = T2209 ? counts_359 : counts_358;
  assign T10703 = reset ? 4'h0 : T2201;
  assign T2201 = T2203 ? T52 : T2202;
  assign T2202 = io_resetCounts ? 4'h0 : counts_358;
  assign T2203 = T10320 & T2204;
  assign T2204 = T76[9'h166:9'h166];
  assign T10704 = reset ? 4'h0 : T2205;
  assign T2205 = T2207 ? T52 : T2206;
  assign T2206 = io_resetCounts ? 4'h0 : counts_359;
  assign T2207 = T10320 & T2208;
  assign T2208 = T76[9'h167:9'h167];
  assign T2209 = T68[1'h0:1'h0];
  assign T2210 = T68[1'h1:1'h1];
  assign T2211 = T68[2'h2:2'h2];
  assign T2212 = T2257 ? T2235 : T2213;
  assign T2213 = T2234 ? T2224 : T2214;
  assign T2214 = T2223 ? counts_361 : counts_360;
  assign T10705 = reset ? 4'h0 : T2215;
  assign T2215 = T2217 ? T52 : T2216;
  assign T2216 = io_resetCounts ? 4'h0 : counts_360;
  assign T2217 = T10320 & T2218;
  assign T2218 = T76[9'h168:9'h168];
  assign T10706 = reset ? 4'h0 : T2219;
  assign T2219 = T2221 ? T52 : T2220;
  assign T2220 = io_resetCounts ? 4'h0 : counts_361;
  assign T2221 = T10320 & T2222;
  assign T2222 = T76[9'h169:9'h169];
  assign T2223 = T68[1'h0:1'h0];
  assign T2224 = T2233 ? counts_363 : counts_362;
  assign T10707 = reset ? 4'h0 : T2225;
  assign T2225 = T2227 ? T52 : T2226;
  assign T2226 = io_resetCounts ? 4'h0 : counts_362;
  assign T2227 = T10320 & T2228;
  assign T2228 = T76[9'h16a:9'h16a];
  assign T10708 = reset ? 4'h0 : T2229;
  assign T2229 = T2231 ? T52 : T2230;
  assign T2230 = io_resetCounts ? 4'h0 : counts_363;
  assign T2231 = T10320 & T2232;
  assign T2232 = T76[9'h16b:9'h16b];
  assign T2233 = T68[1'h0:1'h0];
  assign T2234 = T68[1'h1:1'h1];
  assign T2235 = T2256 ? T2246 : T2236;
  assign T2236 = T2245 ? counts_365 : counts_364;
  assign T10709 = reset ? 4'h0 : T2237;
  assign T2237 = T2239 ? T52 : T2238;
  assign T2238 = io_resetCounts ? 4'h0 : counts_364;
  assign T2239 = T10320 & T2240;
  assign T2240 = T76[9'h16c:9'h16c];
  assign T10710 = reset ? 4'h0 : T2241;
  assign T2241 = T2243 ? T52 : T2242;
  assign T2242 = io_resetCounts ? 4'h0 : counts_365;
  assign T2243 = T10320 & T2244;
  assign T2244 = T76[9'h16d:9'h16d];
  assign T2245 = T68[1'h0:1'h0];
  assign T2246 = T2255 ? counts_367 : counts_366;
  assign T10711 = reset ? 4'h0 : T2247;
  assign T2247 = T2249 ? T52 : T2248;
  assign T2248 = io_resetCounts ? 4'h0 : counts_366;
  assign T2249 = T10320 & T2250;
  assign T2250 = T76[9'h16e:9'h16e];
  assign T10712 = reset ? 4'h0 : T2251;
  assign T2251 = T2253 ? T52 : T2252;
  assign T2252 = io_resetCounts ? 4'h0 : counts_367;
  assign T2253 = T10320 & T2254;
  assign T2254 = T76[9'h16f:9'h16f];
  assign T2255 = T68[1'h0:1'h0];
  assign T2256 = T68[1'h1:1'h1];
  assign T2257 = T68[2'h2:2'h2];
  assign T2258 = T68[2'h3:2'h3];
  assign T2259 = T2352 ? T2306 : T2260;
  assign T2260 = T2305 ? T2283 : T2261;
  assign T2261 = T2282 ? T2272 : T2262;
  assign T2262 = T2271 ? counts_369 : counts_368;
  assign T10713 = reset ? 4'h0 : T2263;
  assign T2263 = T2265 ? T52 : T2264;
  assign T2264 = io_resetCounts ? 4'h0 : counts_368;
  assign T2265 = T10320 & T2266;
  assign T2266 = T76[9'h170:9'h170];
  assign T10714 = reset ? 4'h0 : T2267;
  assign T2267 = T2269 ? T52 : T2268;
  assign T2268 = io_resetCounts ? 4'h0 : counts_369;
  assign T2269 = T10320 & T2270;
  assign T2270 = T76[9'h171:9'h171];
  assign T2271 = T68[1'h0:1'h0];
  assign T2272 = T2281 ? counts_371 : counts_370;
  assign T10715 = reset ? 4'h0 : T2273;
  assign T2273 = T2275 ? T52 : T2274;
  assign T2274 = io_resetCounts ? 4'h0 : counts_370;
  assign T2275 = T10320 & T2276;
  assign T2276 = T76[9'h172:9'h172];
  assign T10716 = reset ? 4'h0 : T2277;
  assign T2277 = T2279 ? T52 : T2278;
  assign T2278 = io_resetCounts ? 4'h0 : counts_371;
  assign T2279 = T10320 & T2280;
  assign T2280 = T76[9'h173:9'h173];
  assign T2281 = T68[1'h0:1'h0];
  assign T2282 = T68[1'h1:1'h1];
  assign T2283 = T2304 ? T2294 : T2284;
  assign T2284 = T2293 ? counts_373 : counts_372;
  assign T10717 = reset ? 4'h0 : T2285;
  assign T2285 = T2287 ? T52 : T2286;
  assign T2286 = io_resetCounts ? 4'h0 : counts_372;
  assign T2287 = T10320 & T2288;
  assign T2288 = T76[9'h174:9'h174];
  assign T10718 = reset ? 4'h0 : T2289;
  assign T2289 = T2291 ? T52 : T2290;
  assign T2290 = io_resetCounts ? 4'h0 : counts_373;
  assign T2291 = T10320 & T2292;
  assign T2292 = T76[9'h175:9'h175];
  assign T2293 = T68[1'h0:1'h0];
  assign T2294 = T2303 ? counts_375 : counts_374;
  assign T10719 = reset ? 4'h0 : T2295;
  assign T2295 = T2297 ? T52 : T2296;
  assign T2296 = io_resetCounts ? 4'h0 : counts_374;
  assign T2297 = T10320 & T2298;
  assign T2298 = T76[9'h176:9'h176];
  assign T10720 = reset ? 4'h0 : T2299;
  assign T2299 = T2301 ? T52 : T2300;
  assign T2300 = io_resetCounts ? 4'h0 : counts_375;
  assign T2301 = T10320 & T2302;
  assign T2302 = T76[9'h177:9'h177];
  assign T2303 = T68[1'h0:1'h0];
  assign T2304 = T68[1'h1:1'h1];
  assign T2305 = T68[2'h2:2'h2];
  assign T2306 = T2351 ? T2329 : T2307;
  assign T2307 = T2328 ? T2318 : T2308;
  assign T2308 = T2317 ? counts_377 : counts_376;
  assign T10721 = reset ? 4'h0 : T2309;
  assign T2309 = T2311 ? T52 : T2310;
  assign T2310 = io_resetCounts ? 4'h0 : counts_376;
  assign T2311 = T10320 & T2312;
  assign T2312 = T76[9'h178:9'h178];
  assign T10722 = reset ? 4'h0 : T2313;
  assign T2313 = T2315 ? T52 : T2314;
  assign T2314 = io_resetCounts ? 4'h0 : counts_377;
  assign T2315 = T10320 & T2316;
  assign T2316 = T76[9'h179:9'h179];
  assign T2317 = T68[1'h0:1'h0];
  assign T2318 = T2327 ? counts_379 : counts_378;
  assign T10723 = reset ? 4'h0 : T2319;
  assign T2319 = T2321 ? T52 : T2320;
  assign T2320 = io_resetCounts ? 4'h0 : counts_378;
  assign T2321 = T10320 & T2322;
  assign T2322 = T76[9'h17a:9'h17a];
  assign T10724 = reset ? 4'h0 : T2323;
  assign T2323 = T2325 ? T52 : T2324;
  assign T2324 = io_resetCounts ? 4'h0 : counts_379;
  assign T2325 = T10320 & T2326;
  assign T2326 = T76[9'h17b:9'h17b];
  assign T2327 = T68[1'h0:1'h0];
  assign T2328 = T68[1'h1:1'h1];
  assign T2329 = T2350 ? T2340 : T2330;
  assign T2330 = T2339 ? counts_381 : counts_380;
  assign T10725 = reset ? 4'h0 : T2331;
  assign T2331 = T2333 ? T52 : T2332;
  assign T2332 = io_resetCounts ? 4'h0 : counts_380;
  assign T2333 = T10320 & T2334;
  assign T2334 = T76[9'h17c:9'h17c];
  assign T10726 = reset ? 4'h0 : T2335;
  assign T2335 = T2337 ? T52 : T2336;
  assign T2336 = io_resetCounts ? 4'h0 : counts_381;
  assign T2337 = T10320 & T2338;
  assign T2338 = T76[9'h17d:9'h17d];
  assign T2339 = T68[1'h0:1'h0];
  assign T2340 = T2349 ? counts_383 : counts_382;
  assign T10727 = reset ? 4'h0 : T2341;
  assign T2341 = T2343 ? T52 : T2342;
  assign T2342 = io_resetCounts ? 4'h0 : counts_382;
  assign T2343 = T10320 & T2344;
  assign T2344 = T76[9'h17e:9'h17e];
  assign T10728 = reset ? 4'h0 : T2345;
  assign T2345 = T2347 ? T52 : T2346;
  assign T2346 = io_resetCounts ? 4'h0 : counts_383;
  assign T2347 = T10320 & T2348;
  assign T2348 = T76[9'h17f:9'h17f];
  assign T2349 = T68[1'h0:1'h0];
  assign T2350 = T68[1'h1:1'h1];
  assign T2351 = T68[2'h2:2'h2];
  assign T2352 = T68[2'h3:2'h3];
  assign T2353 = T68[3'h4:3'h4];
  assign T2354 = T68[3'h5:3'h5];
  assign T2355 = T68[3'h6:3'h6];
  assign T2356 = T3121 ? T2739 : T2357;
  assign T2357 = T2738 ? T2548 : T2358;
  assign T2358 = T2547 ? T2453 : T2359;
  assign T2359 = T2452 ? T2406 : T2360;
  assign T2360 = T2405 ? T2383 : T2361;
  assign T2361 = T2382 ? T2372 : T2362;
  assign T2362 = T2371 ? counts_385 : counts_384;
  assign T10729 = reset ? 4'h0 : T2363;
  assign T2363 = T2365 ? T52 : T2364;
  assign T2364 = io_resetCounts ? 4'h0 : counts_384;
  assign T2365 = T10320 & T2366;
  assign T2366 = T76[9'h180:9'h180];
  assign T10730 = reset ? 4'h0 : T2367;
  assign T2367 = T2369 ? T52 : T2368;
  assign T2368 = io_resetCounts ? 4'h0 : counts_385;
  assign T2369 = T10320 & T2370;
  assign T2370 = T76[9'h181:9'h181];
  assign T2371 = T68[1'h0:1'h0];
  assign T2372 = T2381 ? counts_387 : counts_386;
  assign T10731 = reset ? 4'h0 : T2373;
  assign T2373 = T2375 ? T52 : T2374;
  assign T2374 = io_resetCounts ? 4'h0 : counts_386;
  assign T2375 = T10320 & T2376;
  assign T2376 = T76[9'h182:9'h182];
  assign T10732 = reset ? 4'h0 : T2377;
  assign T2377 = T2379 ? T52 : T2378;
  assign T2378 = io_resetCounts ? 4'h0 : counts_387;
  assign T2379 = T10320 & T2380;
  assign T2380 = T76[9'h183:9'h183];
  assign T2381 = T68[1'h0:1'h0];
  assign T2382 = T68[1'h1:1'h1];
  assign T2383 = T2404 ? T2394 : T2384;
  assign T2384 = T2393 ? counts_389 : counts_388;
  assign T10733 = reset ? 4'h0 : T2385;
  assign T2385 = T2387 ? T52 : T2386;
  assign T2386 = io_resetCounts ? 4'h0 : counts_388;
  assign T2387 = T10320 & T2388;
  assign T2388 = T76[9'h184:9'h184];
  assign T10734 = reset ? 4'h0 : T2389;
  assign T2389 = T2391 ? T52 : T2390;
  assign T2390 = io_resetCounts ? 4'h0 : counts_389;
  assign T2391 = T10320 & T2392;
  assign T2392 = T76[9'h185:9'h185];
  assign T2393 = T68[1'h0:1'h0];
  assign T2394 = T2403 ? counts_391 : counts_390;
  assign T10735 = reset ? 4'h0 : T2395;
  assign T2395 = T2397 ? T52 : T2396;
  assign T2396 = io_resetCounts ? 4'h0 : counts_390;
  assign T2397 = T10320 & T2398;
  assign T2398 = T76[9'h186:9'h186];
  assign T10736 = reset ? 4'h0 : T2399;
  assign T2399 = T2401 ? T52 : T2400;
  assign T2400 = io_resetCounts ? 4'h0 : counts_391;
  assign T2401 = T10320 & T2402;
  assign T2402 = T76[9'h187:9'h187];
  assign T2403 = T68[1'h0:1'h0];
  assign T2404 = T68[1'h1:1'h1];
  assign T2405 = T68[2'h2:2'h2];
  assign T2406 = T2451 ? T2429 : T2407;
  assign T2407 = T2428 ? T2418 : T2408;
  assign T2408 = T2417 ? counts_393 : counts_392;
  assign T10737 = reset ? 4'h0 : T2409;
  assign T2409 = T2411 ? T52 : T2410;
  assign T2410 = io_resetCounts ? 4'h0 : counts_392;
  assign T2411 = T10320 & T2412;
  assign T2412 = T76[9'h188:9'h188];
  assign T10738 = reset ? 4'h0 : T2413;
  assign T2413 = T2415 ? T52 : T2414;
  assign T2414 = io_resetCounts ? 4'h0 : counts_393;
  assign T2415 = T10320 & T2416;
  assign T2416 = T76[9'h189:9'h189];
  assign T2417 = T68[1'h0:1'h0];
  assign T2418 = T2427 ? counts_395 : counts_394;
  assign T10739 = reset ? 4'h0 : T2419;
  assign T2419 = T2421 ? T52 : T2420;
  assign T2420 = io_resetCounts ? 4'h0 : counts_394;
  assign T2421 = T10320 & T2422;
  assign T2422 = T76[9'h18a:9'h18a];
  assign T10740 = reset ? 4'h0 : T2423;
  assign T2423 = T2425 ? T52 : T2424;
  assign T2424 = io_resetCounts ? 4'h0 : counts_395;
  assign T2425 = T10320 & T2426;
  assign T2426 = T76[9'h18b:9'h18b];
  assign T2427 = T68[1'h0:1'h0];
  assign T2428 = T68[1'h1:1'h1];
  assign T2429 = T2450 ? T2440 : T2430;
  assign T2430 = T2439 ? counts_397 : counts_396;
  assign T10741 = reset ? 4'h0 : T2431;
  assign T2431 = T2433 ? T52 : T2432;
  assign T2432 = io_resetCounts ? 4'h0 : counts_396;
  assign T2433 = T10320 & T2434;
  assign T2434 = T76[9'h18c:9'h18c];
  assign T10742 = reset ? 4'h0 : T2435;
  assign T2435 = T2437 ? T52 : T2436;
  assign T2436 = io_resetCounts ? 4'h0 : counts_397;
  assign T2437 = T10320 & T2438;
  assign T2438 = T76[9'h18d:9'h18d];
  assign T2439 = T68[1'h0:1'h0];
  assign T2440 = T2449 ? counts_399 : counts_398;
  assign T10743 = reset ? 4'h0 : T2441;
  assign T2441 = T2443 ? T52 : T2442;
  assign T2442 = io_resetCounts ? 4'h0 : counts_398;
  assign T2443 = T10320 & T2444;
  assign T2444 = T76[9'h18e:9'h18e];
  assign T10744 = reset ? 4'h0 : T2445;
  assign T2445 = T2447 ? T52 : T2446;
  assign T2446 = io_resetCounts ? 4'h0 : counts_399;
  assign T2447 = T10320 & T2448;
  assign T2448 = T76[9'h18f:9'h18f];
  assign T2449 = T68[1'h0:1'h0];
  assign T2450 = T68[1'h1:1'h1];
  assign T2451 = T68[2'h2:2'h2];
  assign T2452 = T68[2'h3:2'h3];
  assign T2453 = T2546 ? T2500 : T2454;
  assign T2454 = T2499 ? T2477 : T2455;
  assign T2455 = T2476 ? T2466 : T2456;
  assign T2456 = T2465 ? counts_401 : counts_400;
  assign T10745 = reset ? 4'h0 : T2457;
  assign T2457 = T2459 ? T52 : T2458;
  assign T2458 = io_resetCounts ? 4'h0 : counts_400;
  assign T2459 = T10320 & T2460;
  assign T2460 = T76[9'h190:9'h190];
  assign T10746 = reset ? 4'h0 : T2461;
  assign T2461 = T2463 ? T52 : T2462;
  assign T2462 = io_resetCounts ? 4'h0 : counts_401;
  assign T2463 = T10320 & T2464;
  assign T2464 = T76[9'h191:9'h191];
  assign T2465 = T68[1'h0:1'h0];
  assign T2466 = T2475 ? counts_403 : counts_402;
  assign T10747 = reset ? 4'h0 : T2467;
  assign T2467 = T2469 ? T52 : T2468;
  assign T2468 = io_resetCounts ? 4'h0 : counts_402;
  assign T2469 = T10320 & T2470;
  assign T2470 = T76[9'h192:9'h192];
  assign T10748 = reset ? 4'h0 : T2471;
  assign T2471 = T2473 ? T52 : T2472;
  assign T2472 = io_resetCounts ? 4'h0 : counts_403;
  assign T2473 = T10320 & T2474;
  assign T2474 = T76[9'h193:9'h193];
  assign T2475 = T68[1'h0:1'h0];
  assign T2476 = T68[1'h1:1'h1];
  assign T2477 = T2498 ? T2488 : T2478;
  assign T2478 = T2487 ? counts_405 : counts_404;
  assign T10749 = reset ? 4'h0 : T2479;
  assign T2479 = T2481 ? T52 : T2480;
  assign T2480 = io_resetCounts ? 4'h0 : counts_404;
  assign T2481 = T10320 & T2482;
  assign T2482 = T76[9'h194:9'h194];
  assign T10750 = reset ? 4'h0 : T2483;
  assign T2483 = T2485 ? T52 : T2484;
  assign T2484 = io_resetCounts ? 4'h0 : counts_405;
  assign T2485 = T10320 & T2486;
  assign T2486 = T76[9'h195:9'h195];
  assign T2487 = T68[1'h0:1'h0];
  assign T2488 = T2497 ? counts_407 : counts_406;
  assign T10751 = reset ? 4'h0 : T2489;
  assign T2489 = T2491 ? T52 : T2490;
  assign T2490 = io_resetCounts ? 4'h0 : counts_406;
  assign T2491 = T10320 & T2492;
  assign T2492 = T76[9'h196:9'h196];
  assign T10752 = reset ? 4'h0 : T2493;
  assign T2493 = T2495 ? T52 : T2494;
  assign T2494 = io_resetCounts ? 4'h0 : counts_407;
  assign T2495 = T10320 & T2496;
  assign T2496 = T76[9'h197:9'h197];
  assign T2497 = T68[1'h0:1'h0];
  assign T2498 = T68[1'h1:1'h1];
  assign T2499 = T68[2'h2:2'h2];
  assign T2500 = T2545 ? T2523 : T2501;
  assign T2501 = T2522 ? T2512 : T2502;
  assign T2502 = T2511 ? counts_409 : counts_408;
  assign T10753 = reset ? 4'h0 : T2503;
  assign T2503 = T2505 ? T52 : T2504;
  assign T2504 = io_resetCounts ? 4'h0 : counts_408;
  assign T2505 = T10320 & T2506;
  assign T2506 = T76[9'h198:9'h198];
  assign T10754 = reset ? 4'h0 : T2507;
  assign T2507 = T2509 ? T52 : T2508;
  assign T2508 = io_resetCounts ? 4'h0 : counts_409;
  assign T2509 = T10320 & T2510;
  assign T2510 = T76[9'h199:9'h199];
  assign T2511 = T68[1'h0:1'h0];
  assign T2512 = T2521 ? counts_411 : counts_410;
  assign T10755 = reset ? 4'h0 : T2513;
  assign T2513 = T2515 ? T52 : T2514;
  assign T2514 = io_resetCounts ? 4'h0 : counts_410;
  assign T2515 = T10320 & T2516;
  assign T2516 = T76[9'h19a:9'h19a];
  assign T10756 = reset ? 4'h0 : T2517;
  assign T2517 = T2519 ? T52 : T2518;
  assign T2518 = io_resetCounts ? 4'h0 : counts_411;
  assign T2519 = T10320 & T2520;
  assign T2520 = T76[9'h19b:9'h19b];
  assign T2521 = T68[1'h0:1'h0];
  assign T2522 = T68[1'h1:1'h1];
  assign T2523 = T2544 ? T2534 : T2524;
  assign T2524 = T2533 ? counts_413 : counts_412;
  assign T10757 = reset ? 4'h0 : T2525;
  assign T2525 = T2527 ? T52 : T2526;
  assign T2526 = io_resetCounts ? 4'h0 : counts_412;
  assign T2527 = T10320 & T2528;
  assign T2528 = T76[9'h19c:9'h19c];
  assign T10758 = reset ? 4'h0 : T2529;
  assign T2529 = T2531 ? T52 : T2530;
  assign T2530 = io_resetCounts ? 4'h0 : counts_413;
  assign T2531 = T10320 & T2532;
  assign T2532 = T76[9'h19d:9'h19d];
  assign T2533 = T68[1'h0:1'h0];
  assign T2534 = T2543 ? counts_415 : counts_414;
  assign T10759 = reset ? 4'h0 : T2535;
  assign T2535 = T2537 ? T52 : T2536;
  assign T2536 = io_resetCounts ? 4'h0 : counts_414;
  assign T2537 = T10320 & T2538;
  assign T2538 = T76[9'h19e:9'h19e];
  assign T10760 = reset ? 4'h0 : T2539;
  assign T2539 = T2541 ? T52 : T2540;
  assign T2540 = io_resetCounts ? 4'h0 : counts_415;
  assign T2541 = T10320 & T2542;
  assign T2542 = T76[9'h19f:9'h19f];
  assign T2543 = T68[1'h0:1'h0];
  assign T2544 = T68[1'h1:1'h1];
  assign T2545 = T68[2'h2:2'h2];
  assign T2546 = T68[2'h3:2'h3];
  assign T2547 = T68[3'h4:3'h4];
  assign T2548 = T2737 ? T2643 : T2549;
  assign T2549 = T2642 ? T2596 : T2550;
  assign T2550 = T2595 ? T2573 : T2551;
  assign T2551 = T2572 ? T2562 : T2552;
  assign T2552 = T2561 ? counts_417 : counts_416;
  assign T10761 = reset ? 4'h0 : T2553;
  assign T2553 = T2555 ? T52 : T2554;
  assign T2554 = io_resetCounts ? 4'h0 : counts_416;
  assign T2555 = T10320 & T2556;
  assign T2556 = T76[9'h1a0:9'h1a0];
  assign T10762 = reset ? 4'h0 : T2557;
  assign T2557 = T2559 ? T52 : T2558;
  assign T2558 = io_resetCounts ? 4'h0 : counts_417;
  assign T2559 = T10320 & T2560;
  assign T2560 = T76[9'h1a1:9'h1a1];
  assign T2561 = T68[1'h0:1'h0];
  assign T2562 = T2571 ? counts_419 : counts_418;
  assign T10763 = reset ? 4'h0 : T2563;
  assign T2563 = T2565 ? T52 : T2564;
  assign T2564 = io_resetCounts ? 4'h0 : counts_418;
  assign T2565 = T10320 & T2566;
  assign T2566 = T76[9'h1a2:9'h1a2];
  assign T10764 = reset ? 4'h0 : T2567;
  assign T2567 = T2569 ? T52 : T2568;
  assign T2568 = io_resetCounts ? 4'h0 : counts_419;
  assign T2569 = T10320 & T2570;
  assign T2570 = T76[9'h1a3:9'h1a3];
  assign T2571 = T68[1'h0:1'h0];
  assign T2572 = T68[1'h1:1'h1];
  assign T2573 = T2594 ? T2584 : T2574;
  assign T2574 = T2583 ? counts_421 : counts_420;
  assign T10765 = reset ? 4'h0 : T2575;
  assign T2575 = T2577 ? T52 : T2576;
  assign T2576 = io_resetCounts ? 4'h0 : counts_420;
  assign T2577 = T10320 & T2578;
  assign T2578 = T76[9'h1a4:9'h1a4];
  assign T10766 = reset ? 4'h0 : T2579;
  assign T2579 = T2581 ? T52 : T2580;
  assign T2580 = io_resetCounts ? 4'h0 : counts_421;
  assign T2581 = T10320 & T2582;
  assign T2582 = T76[9'h1a5:9'h1a5];
  assign T2583 = T68[1'h0:1'h0];
  assign T2584 = T2593 ? counts_423 : counts_422;
  assign T10767 = reset ? 4'h0 : T2585;
  assign T2585 = T2587 ? T52 : T2586;
  assign T2586 = io_resetCounts ? 4'h0 : counts_422;
  assign T2587 = T10320 & T2588;
  assign T2588 = T76[9'h1a6:9'h1a6];
  assign T10768 = reset ? 4'h0 : T2589;
  assign T2589 = T2591 ? T52 : T2590;
  assign T2590 = io_resetCounts ? 4'h0 : counts_423;
  assign T2591 = T10320 & T2592;
  assign T2592 = T76[9'h1a7:9'h1a7];
  assign T2593 = T68[1'h0:1'h0];
  assign T2594 = T68[1'h1:1'h1];
  assign T2595 = T68[2'h2:2'h2];
  assign T2596 = T2641 ? T2619 : T2597;
  assign T2597 = T2618 ? T2608 : T2598;
  assign T2598 = T2607 ? counts_425 : counts_424;
  assign T10769 = reset ? 4'h0 : T2599;
  assign T2599 = T2601 ? T52 : T2600;
  assign T2600 = io_resetCounts ? 4'h0 : counts_424;
  assign T2601 = T10320 & T2602;
  assign T2602 = T76[9'h1a8:9'h1a8];
  assign T10770 = reset ? 4'h0 : T2603;
  assign T2603 = T2605 ? T52 : T2604;
  assign T2604 = io_resetCounts ? 4'h0 : counts_425;
  assign T2605 = T10320 & T2606;
  assign T2606 = T76[9'h1a9:9'h1a9];
  assign T2607 = T68[1'h0:1'h0];
  assign T2608 = T2617 ? counts_427 : counts_426;
  assign T10771 = reset ? 4'h0 : T2609;
  assign T2609 = T2611 ? T52 : T2610;
  assign T2610 = io_resetCounts ? 4'h0 : counts_426;
  assign T2611 = T10320 & T2612;
  assign T2612 = T76[9'h1aa:9'h1aa];
  assign T10772 = reset ? 4'h0 : T2613;
  assign T2613 = T2615 ? T52 : T2614;
  assign T2614 = io_resetCounts ? 4'h0 : counts_427;
  assign T2615 = T10320 & T2616;
  assign T2616 = T76[9'h1ab:9'h1ab];
  assign T2617 = T68[1'h0:1'h0];
  assign T2618 = T68[1'h1:1'h1];
  assign T2619 = T2640 ? T2630 : T2620;
  assign T2620 = T2629 ? counts_429 : counts_428;
  assign T10773 = reset ? 4'h0 : T2621;
  assign T2621 = T2623 ? T52 : T2622;
  assign T2622 = io_resetCounts ? 4'h0 : counts_428;
  assign T2623 = T10320 & T2624;
  assign T2624 = T76[9'h1ac:9'h1ac];
  assign T10774 = reset ? 4'h0 : T2625;
  assign T2625 = T2627 ? T52 : T2626;
  assign T2626 = io_resetCounts ? 4'h0 : counts_429;
  assign T2627 = T10320 & T2628;
  assign T2628 = T76[9'h1ad:9'h1ad];
  assign T2629 = T68[1'h0:1'h0];
  assign T2630 = T2639 ? counts_431 : counts_430;
  assign T10775 = reset ? 4'h0 : T2631;
  assign T2631 = T2633 ? T52 : T2632;
  assign T2632 = io_resetCounts ? 4'h0 : counts_430;
  assign T2633 = T10320 & T2634;
  assign T2634 = T76[9'h1ae:9'h1ae];
  assign T10776 = reset ? 4'h0 : T2635;
  assign T2635 = T2637 ? T52 : T2636;
  assign T2636 = io_resetCounts ? 4'h0 : counts_431;
  assign T2637 = T10320 & T2638;
  assign T2638 = T76[9'h1af:9'h1af];
  assign T2639 = T68[1'h0:1'h0];
  assign T2640 = T68[1'h1:1'h1];
  assign T2641 = T68[2'h2:2'h2];
  assign T2642 = T68[2'h3:2'h3];
  assign T2643 = T2736 ? T2690 : T2644;
  assign T2644 = T2689 ? T2667 : T2645;
  assign T2645 = T2666 ? T2656 : T2646;
  assign T2646 = T2655 ? counts_433 : counts_432;
  assign T10777 = reset ? 4'h0 : T2647;
  assign T2647 = T2649 ? T52 : T2648;
  assign T2648 = io_resetCounts ? 4'h0 : counts_432;
  assign T2649 = T10320 & T2650;
  assign T2650 = T76[9'h1b0:9'h1b0];
  assign T10778 = reset ? 4'h0 : T2651;
  assign T2651 = T2653 ? T52 : T2652;
  assign T2652 = io_resetCounts ? 4'h0 : counts_433;
  assign T2653 = T10320 & T2654;
  assign T2654 = T76[9'h1b1:9'h1b1];
  assign T2655 = T68[1'h0:1'h0];
  assign T2656 = T2665 ? counts_435 : counts_434;
  assign T10779 = reset ? 4'h0 : T2657;
  assign T2657 = T2659 ? T52 : T2658;
  assign T2658 = io_resetCounts ? 4'h0 : counts_434;
  assign T2659 = T10320 & T2660;
  assign T2660 = T76[9'h1b2:9'h1b2];
  assign T10780 = reset ? 4'h0 : T2661;
  assign T2661 = T2663 ? T52 : T2662;
  assign T2662 = io_resetCounts ? 4'h0 : counts_435;
  assign T2663 = T10320 & T2664;
  assign T2664 = T76[9'h1b3:9'h1b3];
  assign T2665 = T68[1'h0:1'h0];
  assign T2666 = T68[1'h1:1'h1];
  assign T2667 = T2688 ? T2678 : T2668;
  assign T2668 = T2677 ? counts_437 : counts_436;
  assign T10781 = reset ? 4'h0 : T2669;
  assign T2669 = T2671 ? T52 : T2670;
  assign T2670 = io_resetCounts ? 4'h0 : counts_436;
  assign T2671 = T10320 & T2672;
  assign T2672 = T76[9'h1b4:9'h1b4];
  assign T10782 = reset ? 4'h0 : T2673;
  assign T2673 = T2675 ? T52 : T2674;
  assign T2674 = io_resetCounts ? 4'h0 : counts_437;
  assign T2675 = T10320 & T2676;
  assign T2676 = T76[9'h1b5:9'h1b5];
  assign T2677 = T68[1'h0:1'h0];
  assign T2678 = T2687 ? counts_439 : counts_438;
  assign T10783 = reset ? 4'h0 : T2679;
  assign T2679 = T2681 ? T52 : T2680;
  assign T2680 = io_resetCounts ? 4'h0 : counts_438;
  assign T2681 = T10320 & T2682;
  assign T2682 = T76[9'h1b6:9'h1b6];
  assign T10784 = reset ? 4'h0 : T2683;
  assign T2683 = T2685 ? T52 : T2684;
  assign T2684 = io_resetCounts ? 4'h0 : counts_439;
  assign T2685 = T10320 & T2686;
  assign T2686 = T76[9'h1b7:9'h1b7];
  assign T2687 = T68[1'h0:1'h0];
  assign T2688 = T68[1'h1:1'h1];
  assign T2689 = T68[2'h2:2'h2];
  assign T2690 = T2735 ? T2713 : T2691;
  assign T2691 = T2712 ? T2702 : T2692;
  assign T2692 = T2701 ? counts_441 : counts_440;
  assign T10785 = reset ? 4'h0 : T2693;
  assign T2693 = T2695 ? T52 : T2694;
  assign T2694 = io_resetCounts ? 4'h0 : counts_440;
  assign T2695 = T10320 & T2696;
  assign T2696 = T76[9'h1b8:9'h1b8];
  assign T10786 = reset ? 4'h0 : T2697;
  assign T2697 = T2699 ? T52 : T2698;
  assign T2698 = io_resetCounts ? 4'h0 : counts_441;
  assign T2699 = T10320 & T2700;
  assign T2700 = T76[9'h1b9:9'h1b9];
  assign T2701 = T68[1'h0:1'h0];
  assign T2702 = T2711 ? counts_443 : counts_442;
  assign T10787 = reset ? 4'h0 : T2703;
  assign T2703 = T2705 ? T52 : T2704;
  assign T2704 = io_resetCounts ? 4'h0 : counts_442;
  assign T2705 = T10320 & T2706;
  assign T2706 = T76[9'h1ba:9'h1ba];
  assign T10788 = reset ? 4'h0 : T2707;
  assign T2707 = T2709 ? T52 : T2708;
  assign T2708 = io_resetCounts ? 4'h0 : counts_443;
  assign T2709 = T10320 & T2710;
  assign T2710 = T76[9'h1bb:9'h1bb];
  assign T2711 = T68[1'h0:1'h0];
  assign T2712 = T68[1'h1:1'h1];
  assign T2713 = T2734 ? T2724 : T2714;
  assign T2714 = T2723 ? counts_445 : counts_444;
  assign T10789 = reset ? 4'h0 : T2715;
  assign T2715 = T2717 ? T52 : T2716;
  assign T2716 = io_resetCounts ? 4'h0 : counts_444;
  assign T2717 = T10320 & T2718;
  assign T2718 = T76[9'h1bc:9'h1bc];
  assign T10790 = reset ? 4'h0 : T2719;
  assign T2719 = T2721 ? T52 : T2720;
  assign T2720 = io_resetCounts ? 4'h0 : counts_445;
  assign T2721 = T10320 & T2722;
  assign T2722 = T76[9'h1bd:9'h1bd];
  assign T2723 = T68[1'h0:1'h0];
  assign T2724 = T2733 ? counts_447 : counts_446;
  assign T10791 = reset ? 4'h0 : T2725;
  assign T2725 = T2727 ? T52 : T2726;
  assign T2726 = io_resetCounts ? 4'h0 : counts_446;
  assign T2727 = T10320 & T2728;
  assign T2728 = T76[9'h1be:9'h1be];
  assign T10792 = reset ? 4'h0 : T2729;
  assign T2729 = T2731 ? T52 : T2730;
  assign T2730 = io_resetCounts ? 4'h0 : counts_447;
  assign T2731 = T10320 & T2732;
  assign T2732 = T76[9'h1bf:9'h1bf];
  assign T2733 = T68[1'h0:1'h0];
  assign T2734 = T68[1'h1:1'h1];
  assign T2735 = T68[2'h2:2'h2];
  assign T2736 = T68[2'h3:2'h3];
  assign T2737 = T68[3'h4:3'h4];
  assign T2738 = T68[3'h5:3'h5];
  assign T2739 = T3120 ? T2930 : T2740;
  assign T2740 = T2929 ? T2835 : T2741;
  assign T2741 = T2834 ? T2788 : T2742;
  assign T2742 = T2787 ? T2765 : T2743;
  assign T2743 = T2764 ? T2754 : T2744;
  assign T2744 = T2753 ? counts_449 : counts_448;
  assign T10793 = reset ? 4'h0 : T2745;
  assign T2745 = T2747 ? T52 : T2746;
  assign T2746 = io_resetCounts ? 4'h0 : counts_448;
  assign T2747 = T10320 & T2748;
  assign T2748 = T76[9'h1c0:9'h1c0];
  assign T10794 = reset ? 4'h0 : T2749;
  assign T2749 = T2751 ? T52 : T2750;
  assign T2750 = io_resetCounts ? 4'h0 : counts_449;
  assign T2751 = T10320 & T2752;
  assign T2752 = T76[9'h1c1:9'h1c1];
  assign T2753 = T68[1'h0:1'h0];
  assign T2754 = T2763 ? counts_451 : counts_450;
  assign T10795 = reset ? 4'h0 : T2755;
  assign T2755 = T2757 ? T52 : T2756;
  assign T2756 = io_resetCounts ? 4'h0 : counts_450;
  assign T2757 = T10320 & T2758;
  assign T2758 = T76[9'h1c2:9'h1c2];
  assign T10796 = reset ? 4'h0 : T2759;
  assign T2759 = T2761 ? T52 : T2760;
  assign T2760 = io_resetCounts ? 4'h0 : counts_451;
  assign T2761 = T10320 & T2762;
  assign T2762 = T76[9'h1c3:9'h1c3];
  assign T2763 = T68[1'h0:1'h0];
  assign T2764 = T68[1'h1:1'h1];
  assign T2765 = T2786 ? T2776 : T2766;
  assign T2766 = T2775 ? counts_453 : counts_452;
  assign T10797 = reset ? 4'h0 : T2767;
  assign T2767 = T2769 ? T52 : T2768;
  assign T2768 = io_resetCounts ? 4'h0 : counts_452;
  assign T2769 = T10320 & T2770;
  assign T2770 = T76[9'h1c4:9'h1c4];
  assign T10798 = reset ? 4'h0 : T2771;
  assign T2771 = T2773 ? T52 : T2772;
  assign T2772 = io_resetCounts ? 4'h0 : counts_453;
  assign T2773 = T10320 & T2774;
  assign T2774 = T76[9'h1c5:9'h1c5];
  assign T2775 = T68[1'h0:1'h0];
  assign T2776 = T2785 ? counts_455 : counts_454;
  assign T10799 = reset ? 4'h0 : T2777;
  assign T2777 = T2779 ? T52 : T2778;
  assign T2778 = io_resetCounts ? 4'h0 : counts_454;
  assign T2779 = T10320 & T2780;
  assign T2780 = T76[9'h1c6:9'h1c6];
  assign T10800 = reset ? 4'h0 : T2781;
  assign T2781 = T2783 ? T52 : T2782;
  assign T2782 = io_resetCounts ? 4'h0 : counts_455;
  assign T2783 = T10320 & T2784;
  assign T2784 = T76[9'h1c7:9'h1c7];
  assign T2785 = T68[1'h0:1'h0];
  assign T2786 = T68[1'h1:1'h1];
  assign T2787 = T68[2'h2:2'h2];
  assign T2788 = T2833 ? T2811 : T2789;
  assign T2789 = T2810 ? T2800 : T2790;
  assign T2790 = T2799 ? counts_457 : counts_456;
  assign T10801 = reset ? 4'h0 : T2791;
  assign T2791 = T2793 ? T52 : T2792;
  assign T2792 = io_resetCounts ? 4'h0 : counts_456;
  assign T2793 = T10320 & T2794;
  assign T2794 = T76[9'h1c8:9'h1c8];
  assign T10802 = reset ? 4'h0 : T2795;
  assign T2795 = T2797 ? T52 : T2796;
  assign T2796 = io_resetCounts ? 4'h0 : counts_457;
  assign T2797 = T10320 & T2798;
  assign T2798 = T76[9'h1c9:9'h1c9];
  assign T2799 = T68[1'h0:1'h0];
  assign T2800 = T2809 ? counts_459 : counts_458;
  assign T10803 = reset ? 4'h0 : T2801;
  assign T2801 = T2803 ? T52 : T2802;
  assign T2802 = io_resetCounts ? 4'h0 : counts_458;
  assign T2803 = T10320 & T2804;
  assign T2804 = T76[9'h1ca:9'h1ca];
  assign T10804 = reset ? 4'h0 : T2805;
  assign T2805 = T2807 ? T52 : T2806;
  assign T2806 = io_resetCounts ? 4'h0 : counts_459;
  assign T2807 = T10320 & T2808;
  assign T2808 = T76[9'h1cb:9'h1cb];
  assign T2809 = T68[1'h0:1'h0];
  assign T2810 = T68[1'h1:1'h1];
  assign T2811 = T2832 ? T2822 : T2812;
  assign T2812 = T2821 ? counts_461 : counts_460;
  assign T10805 = reset ? 4'h0 : T2813;
  assign T2813 = T2815 ? T52 : T2814;
  assign T2814 = io_resetCounts ? 4'h0 : counts_460;
  assign T2815 = T10320 & T2816;
  assign T2816 = T76[9'h1cc:9'h1cc];
  assign T10806 = reset ? 4'h0 : T2817;
  assign T2817 = T2819 ? T52 : T2818;
  assign T2818 = io_resetCounts ? 4'h0 : counts_461;
  assign T2819 = T10320 & T2820;
  assign T2820 = T76[9'h1cd:9'h1cd];
  assign T2821 = T68[1'h0:1'h0];
  assign T2822 = T2831 ? counts_463 : counts_462;
  assign T10807 = reset ? 4'h0 : T2823;
  assign T2823 = T2825 ? T52 : T2824;
  assign T2824 = io_resetCounts ? 4'h0 : counts_462;
  assign T2825 = T10320 & T2826;
  assign T2826 = T76[9'h1ce:9'h1ce];
  assign T10808 = reset ? 4'h0 : T2827;
  assign T2827 = T2829 ? T52 : T2828;
  assign T2828 = io_resetCounts ? 4'h0 : counts_463;
  assign T2829 = T10320 & T2830;
  assign T2830 = T76[9'h1cf:9'h1cf];
  assign T2831 = T68[1'h0:1'h0];
  assign T2832 = T68[1'h1:1'h1];
  assign T2833 = T68[2'h2:2'h2];
  assign T2834 = T68[2'h3:2'h3];
  assign T2835 = T2928 ? T2882 : T2836;
  assign T2836 = T2881 ? T2859 : T2837;
  assign T2837 = T2858 ? T2848 : T2838;
  assign T2838 = T2847 ? counts_465 : counts_464;
  assign T10809 = reset ? 4'h0 : T2839;
  assign T2839 = T2841 ? T52 : T2840;
  assign T2840 = io_resetCounts ? 4'h0 : counts_464;
  assign T2841 = T10320 & T2842;
  assign T2842 = T76[9'h1d0:9'h1d0];
  assign T10810 = reset ? 4'h0 : T2843;
  assign T2843 = T2845 ? T52 : T2844;
  assign T2844 = io_resetCounts ? 4'h0 : counts_465;
  assign T2845 = T10320 & T2846;
  assign T2846 = T76[9'h1d1:9'h1d1];
  assign T2847 = T68[1'h0:1'h0];
  assign T2848 = T2857 ? counts_467 : counts_466;
  assign T10811 = reset ? 4'h0 : T2849;
  assign T2849 = T2851 ? T52 : T2850;
  assign T2850 = io_resetCounts ? 4'h0 : counts_466;
  assign T2851 = T10320 & T2852;
  assign T2852 = T76[9'h1d2:9'h1d2];
  assign T10812 = reset ? 4'h0 : T2853;
  assign T2853 = T2855 ? T52 : T2854;
  assign T2854 = io_resetCounts ? 4'h0 : counts_467;
  assign T2855 = T10320 & T2856;
  assign T2856 = T76[9'h1d3:9'h1d3];
  assign T2857 = T68[1'h0:1'h0];
  assign T2858 = T68[1'h1:1'h1];
  assign T2859 = T2880 ? T2870 : T2860;
  assign T2860 = T2869 ? counts_469 : counts_468;
  assign T10813 = reset ? 4'h0 : T2861;
  assign T2861 = T2863 ? T52 : T2862;
  assign T2862 = io_resetCounts ? 4'h0 : counts_468;
  assign T2863 = T10320 & T2864;
  assign T2864 = T76[9'h1d4:9'h1d4];
  assign T10814 = reset ? 4'h0 : T2865;
  assign T2865 = T2867 ? T52 : T2866;
  assign T2866 = io_resetCounts ? 4'h0 : counts_469;
  assign T2867 = T10320 & T2868;
  assign T2868 = T76[9'h1d5:9'h1d5];
  assign T2869 = T68[1'h0:1'h0];
  assign T2870 = T2879 ? counts_471 : counts_470;
  assign T10815 = reset ? 4'h0 : T2871;
  assign T2871 = T2873 ? T52 : T2872;
  assign T2872 = io_resetCounts ? 4'h0 : counts_470;
  assign T2873 = T10320 & T2874;
  assign T2874 = T76[9'h1d6:9'h1d6];
  assign T10816 = reset ? 4'h0 : T2875;
  assign T2875 = T2877 ? T52 : T2876;
  assign T2876 = io_resetCounts ? 4'h0 : counts_471;
  assign T2877 = T10320 & T2878;
  assign T2878 = T76[9'h1d7:9'h1d7];
  assign T2879 = T68[1'h0:1'h0];
  assign T2880 = T68[1'h1:1'h1];
  assign T2881 = T68[2'h2:2'h2];
  assign T2882 = T2927 ? T2905 : T2883;
  assign T2883 = T2904 ? T2894 : T2884;
  assign T2884 = T2893 ? counts_473 : counts_472;
  assign T10817 = reset ? 4'h0 : T2885;
  assign T2885 = T2887 ? T52 : T2886;
  assign T2886 = io_resetCounts ? 4'h0 : counts_472;
  assign T2887 = T10320 & T2888;
  assign T2888 = T76[9'h1d8:9'h1d8];
  assign T10818 = reset ? 4'h0 : T2889;
  assign T2889 = T2891 ? T52 : T2890;
  assign T2890 = io_resetCounts ? 4'h0 : counts_473;
  assign T2891 = T10320 & T2892;
  assign T2892 = T76[9'h1d9:9'h1d9];
  assign T2893 = T68[1'h0:1'h0];
  assign T2894 = T2903 ? counts_475 : counts_474;
  assign T10819 = reset ? 4'h0 : T2895;
  assign T2895 = T2897 ? T52 : T2896;
  assign T2896 = io_resetCounts ? 4'h0 : counts_474;
  assign T2897 = T10320 & T2898;
  assign T2898 = T76[9'h1da:9'h1da];
  assign T10820 = reset ? 4'h0 : T2899;
  assign T2899 = T2901 ? T52 : T2900;
  assign T2900 = io_resetCounts ? 4'h0 : counts_475;
  assign T2901 = T10320 & T2902;
  assign T2902 = T76[9'h1db:9'h1db];
  assign T2903 = T68[1'h0:1'h0];
  assign T2904 = T68[1'h1:1'h1];
  assign T2905 = T2926 ? T2916 : T2906;
  assign T2906 = T2915 ? counts_477 : counts_476;
  assign T10821 = reset ? 4'h0 : T2907;
  assign T2907 = T2909 ? T52 : T2908;
  assign T2908 = io_resetCounts ? 4'h0 : counts_476;
  assign T2909 = T10320 & T2910;
  assign T2910 = T76[9'h1dc:9'h1dc];
  assign T10822 = reset ? 4'h0 : T2911;
  assign T2911 = T2913 ? T52 : T2912;
  assign T2912 = io_resetCounts ? 4'h0 : counts_477;
  assign T2913 = T10320 & T2914;
  assign T2914 = T76[9'h1dd:9'h1dd];
  assign T2915 = T68[1'h0:1'h0];
  assign T2916 = T2925 ? counts_479 : counts_478;
  assign T10823 = reset ? 4'h0 : T2917;
  assign T2917 = T2919 ? T52 : T2918;
  assign T2918 = io_resetCounts ? 4'h0 : counts_478;
  assign T2919 = T10320 & T2920;
  assign T2920 = T76[9'h1de:9'h1de];
  assign T10824 = reset ? 4'h0 : T2921;
  assign T2921 = T2923 ? T52 : T2922;
  assign T2922 = io_resetCounts ? 4'h0 : counts_479;
  assign T2923 = T10320 & T2924;
  assign T2924 = T76[9'h1df:9'h1df];
  assign T2925 = T68[1'h0:1'h0];
  assign T2926 = T68[1'h1:1'h1];
  assign T2927 = T68[2'h2:2'h2];
  assign T2928 = T68[2'h3:2'h3];
  assign T2929 = T68[3'h4:3'h4];
  assign T2930 = T3119 ? T3025 : T2931;
  assign T2931 = T3024 ? T2978 : T2932;
  assign T2932 = T2977 ? T2955 : T2933;
  assign T2933 = T2954 ? T2944 : T2934;
  assign T2934 = T2943 ? counts_481 : counts_480;
  assign T10825 = reset ? 4'h0 : T2935;
  assign T2935 = T2937 ? T52 : T2936;
  assign T2936 = io_resetCounts ? 4'h0 : counts_480;
  assign T2937 = T10320 & T2938;
  assign T2938 = T76[9'h1e0:9'h1e0];
  assign T10826 = reset ? 4'h0 : T2939;
  assign T2939 = T2941 ? T52 : T2940;
  assign T2940 = io_resetCounts ? 4'h0 : counts_481;
  assign T2941 = T10320 & T2942;
  assign T2942 = T76[9'h1e1:9'h1e1];
  assign T2943 = T68[1'h0:1'h0];
  assign T2944 = T2953 ? counts_483 : counts_482;
  assign T10827 = reset ? 4'h0 : T2945;
  assign T2945 = T2947 ? T52 : T2946;
  assign T2946 = io_resetCounts ? 4'h0 : counts_482;
  assign T2947 = T10320 & T2948;
  assign T2948 = T76[9'h1e2:9'h1e2];
  assign T10828 = reset ? 4'h0 : T2949;
  assign T2949 = T2951 ? T52 : T2950;
  assign T2950 = io_resetCounts ? 4'h0 : counts_483;
  assign T2951 = T10320 & T2952;
  assign T2952 = T76[9'h1e3:9'h1e3];
  assign T2953 = T68[1'h0:1'h0];
  assign T2954 = T68[1'h1:1'h1];
  assign T2955 = T2976 ? T2966 : T2956;
  assign T2956 = T2965 ? counts_485 : counts_484;
  assign T10829 = reset ? 4'h0 : T2957;
  assign T2957 = T2959 ? T52 : T2958;
  assign T2958 = io_resetCounts ? 4'h0 : counts_484;
  assign T2959 = T10320 & T2960;
  assign T2960 = T76[9'h1e4:9'h1e4];
  assign T10830 = reset ? 4'h0 : T2961;
  assign T2961 = T2963 ? T52 : T2962;
  assign T2962 = io_resetCounts ? 4'h0 : counts_485;
  assign T2963 = T10320 & T2964;
  assign T2964 = T76[9'h1e5:9'h1e5];
  assign T2965 = T68[1'h0:1'h0];
  assign T2966 = T2975 ? counts_487 : counts_486;
  assign T10831 = reset ? 4'h0 : T2967;
  assign T2967 = T2969 ? T52 : T2968;
  assign T2968 = io_resetCounts ? 4'h0 : counts_486;
  assign T2969 = T10320 & T2970;
  assign T2970 = T76[9'h1e6:9'h1e6];
  assign T10832 = reset ? 4'h0 : T2971;
  assign T2971 = T2973 ? T52 : T2972;
  assign T2972 = io_resetCounts ? 4'h0 : counts_487;
  assign T2973 = T10320 & T2974;
  assign T2974 = T76[9'h1e7:9'h1e7];
  assign T2975 = T68[1'h0:1'h0];
  assign T2976 = T68[1'h1:1'h1];
  assign T2977 = T68[2'h2:2'h2];
  assign T2978 = T3023 ? T3001 : T2979;
  assign T2979 = T3000 ? T2990 : T2980;
  assign T2980 = T2989 ? counts_489 : counts_488;
  assign T10833 = reset ? 4'h0 : T2981;
  assign T2981 = T2983 ? T52 : T2982;
  assign T2982 = io_resetCounts ? 4'h0 : counts_488;
  assign T2983 = T10320 & T2984;
  assign T2984 = T76[9'h1e8:9'h1e8];
  assign T10834 = reset ? 4'h0 : T2985;
  assign T2985 = T2987 ? T52 : T2986;
  assign T2986 = io_resetCounts ? 4'h0 : counts_489;
  assign T2987 = T10320 & T2988;
  assign T2988 = T76[9'h1e9:9'h1e9];
  assign T2989 = T68[1'h0:1'h0];
  assign T2990 = T2999 ? counts_491 : counts_490;
  assign T10835 = reset ? 4'h0 : T2991;
  assign T2991 = T2993 ? T52 : T2992;
  assign T2992 = io_resetCounts ? 4'h0 : counts_490;
  assign T2993 = T10320 & T2994;
  assign T2994 = T76[9'h1ea:9'h1ea];
  assign T10836 = reset ? 4'h0 : T2995;
  assign T2995 = T2997 ? T52 : T2996;
  assign T2996 = io_resetCounts ? 4'h0 : counts_491;
  assign T2997 = T10320 & T2998;
  assign T2998 = T76[9'h1eb:9'h1eb];
  assign T2999 = T68[1'h0:1'h0];
  assign T3000 = T68[1'h1:1'h1];
  assign T3001 = T3022 ? T3012 : T3002;
  assign T3002 = T3011 ? counts_493 : counts_492;
  assign T10837 = reset ? 4'h0 : T3003;
  assign T3003 = T3005 ? T52 : T3004;
  assign T3004 = io_resetCounts ? 4'h0 : counts_492;
  assign T3005 = T10320 & T3006;
  assign T3006 = T76[9'h1ec:9'h1ec];
  assign T10838 = reset ? 4'h0 : T3007;
  assign T3007 = T3009 ? T52 : T3008;
  assign T3008 = io_resetCounts ? 4'h0 : counts_493;
  assign T3009 = T10320 & T3010;
  assign T3010 = T76[9'h1ed:9'h1ed];
  assign T3011 = T68[1'h0:1'h0];
  assign T3012 = T3021 ? counts_495 : counts_494;
  assign T10839 = reset ? 4'h0 : T3013;
  assign T3013 = T3015 ? T52 : T3014;
  assign T3014 = io_resetCounts ? 4'h0 : counts_494;
  assign T3015 = T10320 & T3016;
  assign T3016 = T76[9'h1ee:9'h1ee];
  assign T10840 = reset ? 4'h0 : T3017;
  assign T3017 = T3019 ? T52 : T3018;
  assign T3018 = io_resetCounts ? 4'h0 : counts_495;
  assign T3019 = T10320 & T3020;
  assign T3020 = T76[9'h1ef:9'h1ef];
  assign T3021 = T68[1'h0:1'h0];
  assign T3022 = T68[1'h1:1'h1];
  assign T3023 = T68[2'h2:2'h2];
  assign T3024 = T68[2'h3:2'h3];
  assign T3025 = T3118 ? T3072 : T3026;
  assign T3026 = T3071 ? T3049 : T3027;
  assign T3027 = T3048 ? T3038 : T3028;
  assign T3028 = T3037 ? counts_497 : counts_496;
  assign T10841 = reset ? 4'h0 : T3029;
  assign T3029 = T3031 ? T52 : T3030;
  assign T3030 = io_resetCounts ? 4'h0 : counts_496;
  assign T3031 = T10320 & T3032;
  assign T3032 = T76[9'h1f0:9'h1f0];
  assign T10842 = reset ? 4'h0 : T3033;
  assign T3033 = T3035 ? T52 : T3034;
  assign T3034 = io_resetCounts ? 4'h0 : counts_497;
  assign T3035 = T10320 & T3036;
  assign T3036 = T76[9'h1f1:9'h1f1];
  assign T3037 = T68[1'h0:1'h0];
  assign T3038 = T3047 ? counts_499 : counts_498;
  assign T10843 = reset ? 4'h0 : T3039;
  assign T3039 = T3041 ? T52 : T3040;
  assign T3040 = io_resetCounts ? 4'h0 : counts_498;
  assign T3041 = T10320 & T3042;
  assign T3042 = T76[9'h1f2:9'h1f2];
  assign T10844 = reset ? 4'h0 : T3043;
  assign T3043 = T3045 ? T52 : T3044;
  assign T3044 = io_resetCounts ? 4'h0 : counts_499;
  assign T3045 = T10320 & T3046;
  assign T3046 = T76[9'h1f3:9'h1f3];
  assign T3047 = T68[1'h0:1'h0];
  assign T3048 = T68[1'h1:1'h1];
  assign T3049 = T3070 ? T3060 : T3050;
  assign T3050 = T3059 ? counts_501 : counts_500;
  assign T10845 = reset ? 4'h0 : T3051;
  assign T3051 = T3053 ? T52 : T3052;
  assign T3052 = io_resetCounts ? 4'h0 : counts_500;
  assign T3053 = T10320 & T3054;
  assign T3054 = T76[9'h1f4:9'h1f4];
  assign T10846 = reset ? 4'h0 : T3055;
  assign T3055 = T3057 ? T52 : T3056;
  assign T3056 = io_resetCounts ? 4'h0 : counts_501;
  assign T3057 = T10320 & T3058;
  assign T3058 = T76[9'h1f5:9'h1f5];
  assign T3059 = T68[1'h0:1'h0];
  assign T3060 = T3069 ? counts_503 : counts_502;
  assign T10847 = reset ? 4'h0 : T3061;
  assign T3061 = T3063 ? T52 : T3062;
  assign T3062 = io_resetCounts ? 4'h0 : counts_502;
  assign T3063 = T10320 & T3064;
  assign T3064 = T76[9'h1f6:9'h1f6];
  assign T10848 = reset ? 4'h0 : T3065;
  assign T3065 = T3067 ? T52 : T3066;
  assign T3066 = io_resetCounts ? 4'h0 : counts_503;
  assign T3067 = T10320 & T3068;
  assign T3068 = T76[9'h1f7:9'h1f7];
  assign T3069 = T68[1'h0:1'h0];
  assign T3070 = T68[1'h1:1'h1];
  assign T3071 = T68[2'h2:2'h2];
  assign T3072 = T3117 ? T3095 : T3073;
  assign T3073 = T3094 ? T3084 : T3074;
  assign T3074 = T3083 ? counts_505 : counts_504;
  assign T10849 = reset ? 4'h0 : T3075;
  assign T3075 = T3077 ? T52 : T3076;
  assign T3076 = io_resetCounts ? 4'h0 : counts_504;
  assign T3077 = T10320 & T3078;
  assign T3078 = T76[9'h1f8:9'h1f8];
  assign T10850 = reset ? 4'h0 : T3079;
  assign T3079 = T3081 ? T52 : T3080;
  assign T3080 = io_resetCounts ? 4'h0 : counts_505;
  assign T3081 = T10320 & T3082;
  assign T3082 = T76[9'h1f9:9'h1f9];
  assign T3083 = T68[1'h0:1'h0];
  assign T3084 = T3093 ? counts_507 : counts_506;
  assign T10851 = reset ? 4'h0 : T3085;
  assign T3085 = T3087 ? T52 : T3086;
  assign T3086 = io_resetCounts ? 4'h0 : counts_506;
  assign T3087 = T10320 & T3088;
  assign T3088 = T76[9'h1fa:9'h1fa];
  assign T10852 = reset ? 4'h0 : T3089;
  assign T3089 = T3091 ? T52 : T3090;
  assign T3090 = io_resetCounts ? 4'h0 : counts_507;
  assign T3091 = T10320 & T3092;
  assign T3092 = T76[9'h1fb:9'h1fb];
  assign T3093 = T68[1'h0:1'h0];
  assign T3094 = T68[1'h1:1'h1];
  assign T3095 = T3116 ? T3106 : T3096;
  assign T3096 = T3105 ? counts_509 : counts_508;
  assign T10853 = reset ? 4'h0 : T3097;
  assign T3097 = T3099 ? T52 : T3098;
  assign T3098 = io_resetCounts ? 4'h0 : counts_508;
  assign T3099 = T10320 & T3100;
  assign T3100 = T76[9'h1fc:9'h1fc];
  assign T10854 = reset ? 4'h0 : T3101;
  assign T3101 = T3103 ? T52 : T3102;
  assign T3102 = io_resetCounts ? 4'h0 : counts_509;
  assign T3103 = T10320 & T3104;
  assign T3104 = T76[9'h1fd:9'h1fd];
  assign T3105 = T68[1'h0:1'h0];
  assign T3106 = T3115 ? counts_511 : counts_510;
  assign T10855 = reset ? 4'h0 : T3107;
  assign T3107 = T3109 ? T52 : T3108;
  assign T3108 = io_resetCounts ? 4'h0 : counts_510;
  assign T3109 = T10320 & T3110;
  assign T3110 = T76[9'h1fe:9'h1fe];
  assign T10856 = reset ? 4'h0 : T3111;
  assign T3111 = T3113 ? T52 : T3112;
  assign T3112 = io_resetCounts ? 4'h0 : counts_511;
  assign T3113 = T10320 & T3114;
  assign T3114 = T76[9'h1ff:9'h1ff];
  assign T3115 = T68[1'h0:1'h0];
  assign T3116 = T68[1'h1:1'h1];
  assign T3117 = T68[2'h2:2'h2];
  assign T3118 = T68[2'h3:2'h3];
  assign T3119 = T68[3'h4:3'h4];
  assign T3120 = T68[3'h5:3'h5];
  assign T3121 = T68[3'h6:3'h6];
  assign T3122 = T68[3'h7:3'h7];
  assign T3123 = T68[4'h8:4'h8];
  assign T3124 = T6193 ? T4659 : T3125;
  assign T3125 = T4658 ? T3892 : T3126;
  assign T3126 = T3891 ? T3509 : T3127;
  assign T3127 = T3508 ? T3318 : T3128;
  assign T3128 = T3317 ? T3223 : T3129;
  assign T3129 = T3222 ? T3176 : T3130;
  assign T3130 = T3175 ? T3153 : T3131;
  assign T3131 = T3152 ? T3142 : T3132;
  assign T3132 = T3141 ? counts_513 : counts_512;
  assign T10857 = reset ? 4'h0 : T3133;
  assign T3133 = T3135 ? T52 : T3134;
  assign T3134 = io_resetCounts ? 4'h0 : counts_512;
  assign T3135 = T10320 & T3136;
  assign T3136 = T76[10'h200:10'h200];
  assign T10858 = reset ? 4'h0 : T3137;
  assign T3137 = T3139 ? T52 : T3138;
  assign T3138 = io_resetCounts ? 4'h0 : counts_513;
  assign T3139 = T10320 & T3140;
  assign T3140 = T76[10'h201:10'h201];
  assign T3141 = T68[1'h0:1'h0];
  assign T3142 = T3151 ? counts_515 : counts_514;
  assign T10859 = reset ? 4'h0 : T3143;
  assign T3143 = T3145 ? T52 : T3144;
  assign T3144 = io_resetCounts ? 4'h0 : counts_514;
  assign T3145 = T10320 & T3146;
  assign T3146 = T76[10'h202:10'h202];
  assign T10860 = reset ? 4'h0 : T3147;
  assign T3147 = T3149 ? T52 : T3148;
  assign T3148 = io_resetCounts ? 4'h0 : counts_515;
  assign T3149 = T10320 & T3150;
  assign T3150 = T76[10'h203:10'h203];
  assign T3151 = T68[1'h0:1'h0];
  assign T3152 = T68[1'h1:1'h1];
  assign T3153 = T3174 ? T3164 : T3154;
  assign T3154 = T3163 ? counts_517 : counts_516;
  assign T10861 = reset ? 4'h0 : T3155;
  assign T3155 = T3157 ? T52 : T3156;
  assign T3156 = io_resetCounts ? 4'h0 : counts_516;
  assign T3157 = T10320 & T3158;
  assign T3158 = T76[10'h204:10'h204];
  assign T10862 = reset ? 4'h0 : T3159;
  assign T3159 = T3161 ? T52 : T3160;
  assign T3160 = io_resetCounts ? 4'h0 : counts_517;
  assign T3161 = T10320 & T3162;
  assign T3162 = T76[10'h205:10'h205];
  assign T3163 = T68[1'h0:1'h0];
  assign T3164 = T3173 ? counts_519 : counts_518;
  assign T10863 = reset ? 4'h0 : T3165;
  assign T3165 = T3167 ? T52 : T3166;
  assign T3166 = io_resetCounts ? 4'h0 : counts_518;
  assign T3167 = T10320 & T3168;
  assign T3168 = T76[10'h206:10'h206];
  assign T10864 = reset ? 4'h0 : T3169;
  assign T3169 = T3171 ? T52 : T3170;
  assign T3170 = io_resetCounts ? 4'h0 : counts_519;
  assign T3171 = T10320 & T3172;
  assign T3172 = T76[10'h207:10'h207];
  assign T3173 = T68[1'h0:1'h0];
  assign T3174 = T68[1'h1:1'h1];
  assign T3175 = T68[2'h2:2'h2];
  assign T3176 = T3221 ? T3199 : T3177;
  assign T3177 = T3198 ? T3188 : T3178;
  assign T3178 = T3187 ? counts_521 : counts_520;
  assign T10865 = reset ? 4'h0 : T3179;
  assign T3179 = T3181 ? T52 : T3180;
  assign T3180 = io_resetCounts ? 4'h0 : counts_520;
  assign T3181 = T10320 & T3182;
  assign T3182 = T76[10'h208:10'h208];
  assign T10866 = reset ? 4'h0 : T3183;
  assign T3183 = T3185 ? T52 : T3184;
  assign T3184 = io_resetCounts ? 4'h0 : counts_521;
  assign T3185 = T10320 & T3186;
  assign T3186 = T76[10'h209:10'h209];
  assign T3187 = T68[1'h0:1'h0];
  assign T3188 = T3197 ? counts_523 : counts_522;
  assign T10867 = reset ? 4'h0 : T3189;
  assign T3189 = T3191 ? T52 : T3190;
  assign T3190 = io_resetCounts ? 4'h0 : counts_522;
  assign T3191 = T10320 & T3192;
  assign T3192 = T76[10'h20a:10'h20a];
  assign T10868 = reset ? 4'h0 : T3193;
  assign T3193 = T3195 ? T52 : T3194;
  assign T3194 = io_resetCounts ? 4'h0 : counts_523;
  assign T3195 = T10320 & T3196;
  assign T3196 = T76[10'h20b:10'h20b];
  assign T3197 = T68[1'h0:1'h0];
  assign T3198 = T68[1'h1:1'h1];
  assign T3199 = T3220 ? T3210 : T3200;
  assign T3200 = T3209 ? counts_525 : counts_524;
  assign T10869 = reset ? 4'h0 : T3201;
  assign T3201 = T3203 ? T52 : T3202;
  assign T3202 = io_resetCounts ? 4'h0 : counts_524;
  assign T3203 = T10320 & T3204;
  assign T3204 = T76[10'h20c:10'h20c];
  assign T10870 = reset ? 4'h0 : T3205;
  assign T3205 = T3207 ? T52 : T3206;
  assign T3206 = io_resetCounts ? 4'h0 : counts_525;
  assign T3207 = T10320 & T3208;
  assign T3208 = T76[10'h20d:10'h20d];
  assign T3209 = T68[1'h0:1'h0];
  assign T3210 = T3219 ? counts_527 : counts_526;
  assign T10871 = reset ? 4'h0 : T3211;
  assign T3211 = T3213 ? T52 : T3212;
  assign T3212 = io_resetCounts ? 4'h0 : counts_526;
  assign T3213 = T10320 & T3214;
  assign T3214 = T76[10'h20e:10'h20e];
  assign T10872 = reset ? 4'h0 : T3215;
  assign T3215 = T3217 ? T52 : T3216;
  assign T3216 = io_resetCounts ? 4'h0 : counts_527;
  assign T3217 = T10320 & T3218;
  assign T3218 = T76[10'h20f:10'h20f];
  assign T3219 = T68[1'h0:1'h0];
  assign T3220 = T68[1'h1:1'h1];
  assign T3221 = T68[2'h2:2'h2];
  assign T3222 = T68[2'h3:2'h3];
  assign T3223 = T3316 ? T3270 : T3224;
  assign T3224 = T3269 ? T3247 : T3225;
  assign T3225 = T3246 ? T3236 : T3226;
  assign T3226 = T3235 ? counts_529 : counts_528;
  assign T10873 = reset ? 4'h0 : T3227;
  assign T3227 = T3229 ? T52 : T3228;
  assign T3228 = io_resetCounts ? 4'h0 : counts_528;
  assign T3229 = T10320 & T3230;
  assign T3230 = T76[10'h210:10'h210];
  assign T10874 = reset ? 4'h0 : T3231;
  assign T3231 = T3233 ? T52 : T3232;
  assign T3232 = io_resetCounts ? 4'h0 : counts_529;
  assign T3233 = T10320 & T3234;
  assign T3234 = T76[10'h211:10'h211];
  assign T3235 = T68[1'h0:1'h0];
  assign T3236 = T3245 ? counts_531 : counts_530;
  assign T10875 = reset ? 4'h0 : T3237;
  assign T3237 = T3239 ? T52 : T3238;
  assign T3238 = io_resetCounts ? 4'h0 : counts_530;
  assign T3239 = T10320 & T3240;
  assign T3240 = T76[10'h212:10'h212];
  assign T10876 = reset ? 4'h0 : T3241;
  assign T3241 = T3243 ? T52 : T3242;
  assign T3242 = io_resetCounts ? 4'h0 : counts_531;
  assign T3243 = T10320 & T3244;
  assign T3244 = T76[10'h213:10'h213];
  assign T3245 = T68[1'h0:1'h0];
  assign T3246 = T68[1'h1:1'h1];
  assign T3247 = T3268 ? T3258 : T3248;
  assign T3248 = T3257 ? counts_533 : counts_532;
  assign T10877 = reset ? 4'h0 : T3249;
  assign T3249 = T3251 ? T52 : T3250;
  assign T3250 = io_resetCounts ? 4'h0 : counts_532;
  assign T3251 = T10320 & T3252;
  assign T3252 = T76[10'h214:10'h214];
  assign T10878 = reset ? 4'h0 : T3253;
  assign T3253 = T3255 ? T52 : T3254;
  assign T3254 = io_resetCounts ? 4'h0 : counts_533;
  assign T3255 = T10320 & T3256;
  assign T3256 = T76[10'h215:10'h215];
  assign T3257 = T68[1'h0:1'h0];
  assign T3258 = T3267 ? counts_535 : counts_534;
  assign T10879 = reset ? 4'h0 : T3259;
  assign T3259 = T3261 ? T52 : T3260;
  assign T3260 = io_resetCounts ? 4'h0 : counts_534;
  assign T3261 = T10320 & T3262;
  assign T3262 = T76[10'h216:10'h216];
  assign T10880 = reset ? 4'h0 : T3263;
  assign T3263 = T3265 ? T52 : T3264;
  assign T3264 = io_resetCounts ? 4'h0 : counts_535;
  assign T3265 = T10320 & T3266;
  assign T3266 = T76[10'h217:10'h217];
  assign T3267 = T68[1'h0:1'h0];
  assign T3268 = T68[1'h1:1'h1];
  assign T3269 = T68[2'h2:2'h2];
  assign T3270 = T3315 ? T3293 : T3271;
  assign T3271 = T3292 ? T3282 : T3272;
  assign T3272 = T3281 ? counts_537 : counts_536;
  assign T10881 = reset ? 4'h0 : T3273;
  assign T3273 = T3275 ? T52 : T3274;
  assign T3274 = io_resetCounts ? 4'h0 : counts_536;
  assign T3275 = T10320 & T3276;
  assign T3276 = T76[10'h218:10'h218];
  assign T10882 = reset ? 4'h0 : T3277;
  assign T3277 = T3279 ? T52 : T3278;
  assign T3278 = io_resetCounts ? 4'h0 : counts_537;
  assign T3279 = T10320 & T3280;
  assign T3280 = T76[10'h219:10'h219];
  assign T3281 = T68[1'h0:1'h0];
  assign T3282 = T3291 ? counts_539 : counts_538;
  assign T10883 = reset ? 4'h0 : T3283;
  assign T3283 = T3285 ? T52 : T3284;
  assign T3284 = io_resetCounts ? 4'h0 : counts_538;
  assign T3285 = T10320 & T3286;
  assign T3286 = T76[10'h21a:10'h21a];
  assign T10884 = reset ? 4'h0 : T3287;
  assign T3287 = T3289 ? T52 : T3288;
  assign T3288 = io_resetCounts ? 4'h0 : counts_539;
  assign T3289 = T10320 & T3290;
  assign T3290 = T76[10'h21b:10'h21b];
  assign T3291 = T68[1'h0:1'h0];
  assign T3292 = T68[1'h1:1'h1];
  assign T3293 = T3314 ? T3304 : T3294;
  assign T3294 = T3303 ? counts_541 : counts_540;
  assign T10885 = reset ? 4'h0 : T3295;
  assign T3295 = T3297 ? T52 : T3296;
  assign T3296 = io_resetCounts ? 4'h0 : counts_540;
  assign T3297 = T10320 & T3298;
  assign T3298 = T76[10'h21c:10'h21c];
  assign T10886 = reset ? 4'h0 : T3299;
  assign T3299 = T3301 ? T52 : T3300;
  assign T3300 = io_resetCounts ? 4'h0 : counts_541;
  assign T3301 = T10320 & T3302;
  assign T3302 = T76[10'h21d:10'h21d];
  assign T3303 = T68[1'h0:1'h0];
  assign T3304 = T3313 ? counts_543 : counts_542;
  assign T10887 = reset ? 4'h0 : T3305;
  assign T3305 = T3307 ? T52 : T3306;
  assign T3306 = io_resetCounts ? 4'h0 : counts_542;
  assign T3307 = T10320 & T3308;
  assign T3308 = T76[10'h21e:10'h21e];
  assign T10888 = reset ? 4'h0 : T3309;
  assign T3309 = T3311 ? T52 : T3310;
  assign T3310 = io_resetCounts ? 4'h0 : counts_543;
  assign T3311 = T10320 & T3312;
  assign T3312 = T76[10'h21f:10'h21f];
  assign T3313 = T68[1'h0:1'h0];
  assign T3314 = T68[1'h1:1'h1];
  assign T3315 = T68[2'h2:2'h2];
  assign T3316 = T68[2'h3:2'h3];
  assign T3317 = T68[3'h4:3'h4];
  assign T3318 = T3507 ? T3413 : T3319;
  assign T3319 = T3412 ? T3366 : T3320;
  assign T3320 = T3365 ? T3343 : T3321;
  assign T3321 = T3342 ? T3332 : T3322;
  assign T3322 = T3331 ? counts_545 : counts_544;
  assign T10889 = reset ? 4'h0 : T3323;
  assign T3323 = T3325 ? T52 : T3324;
  assign T3324 = io_resetCounts ? 4'h0 : counts_544;
  assign T3325 = T10320 & T3326;
  assign T3326 = T76[10'h220:10'h220];
  assign T10890 = reset ? 4'h0 : T3327;
  assign T3327 = T3329 ? T52 : T3328;
  assign T3328 = io_resetCounts ? 4'h0 : counts_545;
  assign T3329 = T10320 & T3330;
  assign T3330 = T76[10'h221:10'h221];
  assign T3331 = T68[1'h0:1'h0];
  assign T3332 = T3341 ? counts_547 : counts_546;
  assign T10891 = reset ? 4'h0 : T3333;
  assign T3333 = T3335 ? T52 : T3334;
  assign T3334 = io_resetCounts ? 4'h0 : counts_546;
  assign T3335 = T10320 & T3336;
  assign T3336 = T76[10'h222:10'h222];
  assign T10892 = reset ? 4'h0 : T3337;
  assign T3337 = T3339 ? T52 : T3338;
  assign T3338 = io_resetCounts ? 4'h0 : counts_547;
  assign T3339 = T10320 & T3340;
  assign T3340 = T76[10'h223:10'h223];
  assign T3341 = T68[1'h0:1'h0];
  assign T3342 = T68[1'h1:1'h1];
  assign T3343 = T3364 ? T3354 : T3344;
  assign T3344 = T3353 ? counts_549 : counts_548;
  assign T10893 = reset ? 4'h0 : T3345;
  assign T3345 = T3347 ? T52 : T3346;
  assign T3346 = io_resetCounts ? 4'h0 : counts_548;
  assign T3347 = T10320 & T3348;
  assign T3348 = T76[10'h224:10'h224];
  assign T10894 = reset ? 4'h0 : T3349;
  assign T3349 = T3351 ? T52 : T3350;
  assign T3350 = io_resetCounts ? 4'h0 : counts_549;
  assign T3351 = T10320 & T3352;
  assign T3352 = T76[10'h225:10'h225];
  assign T3353 = T68[1'h0:1'h0];
  assign T3354 = T3363 ? counts_551 : counts_550;
  assign T10895 = reset ? 4'h0 : T3355;
  assign T3355 = T3357 ? T52 : T3356;
  assign T3356 = io_resetCounts ? 4'h0 : counts_550;
  assign T3357 = T10320 & T3358;
  assign T3358 = T76[10'h226:10'h226];
  assign T10896 = reset ? 4'h0 : T3359;
  assign T3359 = T3361 ? T52 : T3360;
  assign T3360 = io_resetCounts ? 4'h0 : counts_551;
  assign T3361 = T10320 & T3362;
  assign T3362 = T76[10'h227:10'h227];
  assign T3363 = T68[1'h0:1'h0];
  assign T3364 = T68[1'h1:1'h1];
  assign T3365 = T68[2'h2:2'h2];
  assign T3366 = T3411 ? T3389 : T3367;
  assign T3367 = T3388 ? T3378 : T3368;
  assign T3368 = T3377 ? counts_553 : counts_552;
  assign T10897 = reset ? 4'h0 : T3369;
  assign T3369 = T3371 ? T52 : T3370;
  assign T3370 = io_resetCounts ? 4'h0 : counts_552;
  assign T3371 = T10320 & T3372;
  assign T3372 = T76[10'h228:10'h228];
  assign T10898 = reset ? 4'h0 : T3373;
  assign T3373 = T3375 ? T52 : T3374;
  assign T3374 = io_resetCounts ? 4'h0 : counts_553;
  assign T3375 = T10320 & T3376;
  assign T3376 = T76[10'h229:10'h229];
  assign T3377 = T68[1'h0:1'h0];
  assign T3378 = T3387 ? counts_555 : counts_554;
  assign T10899 = reset ? 4'h0 : T3379;
  assign T3379 = T3381 ? T52 : T3380;
  assign T3380 = io_resetCounts ? 4'h0 : counts_554;
  assign T3381 = T10320 & T3382;
  assign T3382 = T76[10'h22a:10'h22a];
  assign T10900 = reset ? 4'h0 : T3383;
  assign T3383 = T3385 ? T52 : T3384;
  assign T3384 = io_resetCounts ? 4'h0 : counts_555;
  assign T3385 = T10320 & T3386;
  assign T3386 = T76[10'h22b:10'h22b];
  assign T3387 = T68[1'h0:1'h0];
  assign T3388 = T68[1'h1:1'h1];
  assign T3389 = T3410 ? T3400 : T3390;
  assign T3390 = T3399 ? counts_557 : counts_556;
  assign T10901 = reset ? 4'h0 : T3391;
  assign T3391 = T3393 ? T52 : T3392;
  assign T3392 = io_resetCounts ? 4'h0 : counts_556;
  assign T3393 = T10320 & T3394;
  assign T3394 = T76[10'h22c:10'h22c];
  assign T10902 = reset ? 4'h0 : T3395;
  assign T3395 = T3397 ? T52 : T3396;
  assign T3396 = io_resetCounts ? 4'h0 : counts_557;
  assign T3397 = T10320 & T3398;
  assign T3398 = T76[10'h22d:10'h22d];
  assign T3399 = T68[1'h0:1'h0];
  assign T3400 = T3409 ? counts_559 : counts_558;
  assign T10903 = reset ? 4'h0 : T3401;
  assign T3401 = T3403 ? T52 : T3402;
  assign T3402 = io_resetCounts ? 4'h0 : counts_558;
  assign T3403 = T10320 & T3404;
  assign T3404 = T76[10'h22e:10'h22e];
  assign T10904 = reset ? 4'h0 : T3405;
  assign T3405 = T3407 ? T52 : T3406;
  assign T3406 = io_resetCounts ? 4'h0 : counts_559;
  assign T3407 = T10320 & T3408;
  assign T3408 = T76[10'h22f:10'h22f];
  assign T3409 = T68[1'h0:1'h0];
  assign T3410 = T68[1'h1:1'h1];
  assign T3411 = T68[2'h2:2'h2];
  assign T3412 = T68[2'h3:2'h3];
  assign T3413 = T3506 ? T3460 : T3414;
  assign T3414 = T3459 ? T3437 : T3415;
  assign T3415 = T3436 ? T3426 : T3416;
  assign T3416 = T3425 ? counts_561 : counts_560;
  assign T10905 = reset ? 4'h0 : T3417;
  assign T3417 = T3419 ? T52 : T3418;
  assign T3418 = io_resetCounts ? 4'h0 : counts_560;
  assign T3419 = T10320 & T3420;
  assign T3420 = T76[10'h230:10'h230];
  assign T10906 = reset ? 4'h0 : T3421;
  assign T3421 = T3423 ? T52 : T3422;
  assign T3422 = io_resetCounts ? 4'h0 : counts_561;
  assign T3423 = T10320 & T3424;
  assign T3424 = T76[10'h231:10'h231];
  assign T3425 = T68[1'h0:1'h0];
  assign T3426 = T3435 ? counts_563 : counts_562;
  assign T10907 = reset ? 4'h0 : T3427;
  assign T3427 = T3429 ? T52 : T3428;
  assign T3428 = io_resetCounts ? 4'h0 : counts_562;
  assign T3429 = T10320 & T3430;
  assign T3430 = T76[10'h232:10'h232];
  assign T10908 = reset ? 4'h0 : T3431;
  assign T3431 = T3433 ? T52 : T3432;
  assign T3432 = io_resetCounts ? 4'h0 : counts_563;
  assign T3433 = T10320 & T3434;
  assign T3434 = T76[10'h233:10'h233];
  assign T3435 = T68[1'h0:1'h0];
  assign T3436 = T68[1'h1:1'h1];
  assign T3437 = T3458 ? T3448 : T3438;
  assign T3438 = T3447 ? counts_565 : counts_564;
  assign T10909 = reset ? 4'h0 : T3439;
  assign T3439 = T3441 ? T52 : T3440;
  assign T3440 = io_resetCounts ? 4'h0 : counts_564;
  assign T3441 = T10320 & T3442;
  assign T3442 = T76[10'h234:10'h234];
  assign T10910 = reset ? 4'h0 : T3443;
  assign T3443 = T3445 ? T52 : T3444;
  assign T3444 = io_resetCounts ? 4'h0 : counts_565;
  assign T3445 = T10320 & T3446;
  assign T3446 = T76[10'h235:10'h235];
  assign T3447 = T68[1'h0:1'h0];
  assign T3448 = T3457 ? counts_567 : counts_566;
  assign T10911 = reset ? 4'h0 : T3449;
  assign T3449 = T3451 ? T52 : T3450;
  assign T3450 = io_resetCounts ? 4'h0 : counts_566;
  assign T3451 = T10320 & T3452;
  assign T3452 = T76[10'h236:10'h236];
  assign T10912 = reset ? 4'h0 : T3453;
  assign T3453 = T3455 ? T52 : T3454;
  assign T3454 = io_resetCounts ? 4'h0 : counts_567;
  assign T3455 = T10320 & T3456;
  assign T3456 = T76[10'h237:10'h237];
  assign T3457 = T68[1'h0:1'h0];
  assign T3458 = T68[1'h1:1'h1];
  assign T3459 = T68[2'h2:2'h2];
  assign T3460 = T3505 ? T3483 : T3461;
  assign T3461 = T3482 ? T3472 : T3462;
  assign T3462 = T3471 ? counts_569 : counts_568;
  assign T10913 = reset ? 4'h0 : T3463;
  assign T3463 = T3465 ? T52 : T3464;
  assign T3464 = io_resetCounts ? 4'h0 : counts_568;
  assign T3465 = T10320 & T3466;
  assign T3466 = T76[10'h238:10'h238];
  assign T10914 = reset ? 4'h0 : T3467;
  assign T3467 = T3469 ? T52 : T3468;
  assign T3468 = io_resetCounts ? 4'h0 : counts_569;
  assign T3469 = T10320 & T3470;
  assign T3470 = T76[10'h239:10'h239];
  assign T3471 = T68[1'h0:1'h0];
  assign T3472 = T3481 ? counts_571 : counts_570;
  assign T10915 = reset ? 4'h0 : T3473;
  assign T3473 = T3475 ? T52 : T3474;
  assign T3474 = io_resetCounts ? 4'h0 : counts_570;
  assign T3475 = T10320 & T3476;
  assign T3476 = T76[10'h23a:10'h23a];
  assign T10916 = reset ? 4'h0 : T3477;
  assign T3477 = T3479 ? T52 : T3478;
  assign T3478 = io_resetCounts ? 4'h0 : counts_571;
  assign T3479 = T10320 & T3480;
  assign T3480 = T76[10'h23b:10'h23b];
  assign T3481 = T68[1'h0:1'h0];
  assign T3482 = T68[1'h1:1'h1];
  assign T3483 = T3504 ? T3494 : T3484;
  assign T3484 = T3493 ? counts_573 : counts_572;
  assign T10917 = reset ? 4'h0 : T3485;
  assign T3485 = T3487 ? T52 : T3486;
  assign T3486 = io_resetCounts ? 4'h0 : counts_572;
  assign T3487 = T10320 & T3488;
  assign T3488 = T76[10'h23c:10'h23c];
  assign T10918 = reset ? 4'h0 : T3489;
  assign T3489 = T3491 ? T52 : T3490;
  assign T3490 = io_resetCounts ? 4'h0 : counts_573;
  assign T3491 = T10320 & T3492;
  assign T3492 = T76[10'h23d:10'h23d];
  assign T3493 = T68[1'h0:1'h0];
  assign T3494 = T3503 ? counts_575 : counts_574;
  assign T10919 = reset ? 4'h0 : T3495;
  assign T3495 = T3497 ? T52 : T3496;
  assign T3496 = io_resetCounts ? 4'h0 : counts_574;
  assign T3497 = T10320 & T3498;
  assign T3498 = T76[10'h23e:10'h23e];
  assign T10920 = reset ? 4'h0 : T3499;
  assign T3499 = T3501 ? T52 : T3500;
  assign T3500 = io_resetCounts ? 4'h0 : counts_575;
  assign T3501 = T10320 & T3502;
  assign T3502 = T76[10'h23f:10'h23f];
  assign T3503 = T68[1'h0:1'h0];
  assign T3504 = T68[1'h1:1'h1];
  assign T3505 = T68[2'h2:2'h2];
  assign T3506 = T68[2'h3:2'h3];
  assign T3507 = T68[3'h4:3'h4];
  assign T3508 = T68[3'h5:3'h5];
  assign T3509 = T3890 ? T3700 : T3510;
  assign T3510 = T3699 ? T3605 : T3511;
  assign T3511 = T3604 ? T3558 : T3512;
  assign T3512 = T3557 ? T3535 : T3513;
  assign T3513 = T3534 ? T3524 : T3514;
  assign T3514 = T3523 ? counts_577 : counts_576;
  assign T10921 = reset ? 4'h0 : T3515;
  assign T3515 = T3517 ? T52 : T3516;
  assign T3516 = io_resetCounts ? 4'h0 : counts_576;
  assign T3517 = T10320 & T3518;
  assign T3518 = T76[10'h240:10'h240];
  assign T10922 = reset ? 4'h0 : T3519;
  assign T3519 = T3521 ? T52 : T3520;
  assign T3520 = io_resetCounts ? 4'h0 : counts_577;
  assign T3521 = T10320 & T3522;
  assign T3522 = T76[10'h241:10'h241];
  assign T3523 = T68[1'h0:1'h0];
  assign T3524 = T3533 ? counts_579 : counts_578;
  assign T10923 = reset ? 4'h0 : T3525;
  assign T3525 = T3527 ? T52 : T3526;
  assign T3526 = io_resetCounts ? 4'h0 : counts_578;
  assign T3527 = T10320 & T3528;
  assign T3528 = T76[10'h242:10'h242];
  assign T10924 = reset ? 4'h0 : T3529;
  assign T3529 = T3531 ? T52 : T3530;
  assign T3530 = io_resetCounts ? 4'h0 : counts_579;
  assign T3531 = T10320 & T3532;
  assign T3532 = T76[10'h243:10'h243];
  assign T3533 = T68[1'h0:1'h0];
  assign T3534 = T68[1'h1:1'h1];
  assign T3535 = T3556 ? T3546 : T3536;
  assign T3536 = T3545 ? counts_581 : counts_580;
  assign T10925 = reset ? 4'h0 : T3537;
  assign T3537 = T3539 ? T52 : T3538;
  assign T3538 = io_resetCounts ? 4'h0 : counts_580;
  assign T3539 = T10320 & T3540;
  assign T3540 = T76[10'h244:10'h244];
  assign T10926 = reset ? 4'h0 : T3541;
  assign T3541 = T3543 ? T52 : T3542;
  assign T3542 = io_resetCounts ? 4'h0 : counts_581;
  assign T3543 = T10320 & T3544;
  assign T3544 = T76[10'h245:10'h245];
  assign T3545 = T68[1'h0:1'h0];
  assign T3546 = T3555 ? counts_583 : counts_582;
  assign T10927 = reset ? 4'h0 : T3547;
  assign T3547 = T3549 ? T52 : T3548;
  assign T3548 = io_resetCounts ? 4'h0 : counts_582;
  assign T3549 = T10320 & T3550;
  assign T3550 = T76[10'h246:10'h246];
  assign T10928 = reset ? 4'h0 : T3551;
  assign T3551 = T3553 ? T52 : T3552;
  assign T3552 = io_resetCounts ? 4'h0 : counts_583;
  assign T3553 = T10320 & T3554;
  assign T3554 = T76[10'h247:10'h247];
  assign T3555 = T68[1'h0:1'h0];
  assign T3556 = T68[1'h1:1'h1];
  assign T3557 = T68[2'h2:2'h2];
  assign T3558 = T3603 ? T3581 : T3559;
  assign T3559 = T3580 ? T3570 : T3560;
  assign T3560 = T3569 ? counts_585 : counts_584;
  assign T10929 = reset ? 4'h0 : T3561;
  assign T3561 = T3563 ? T52 : T3562;
  assign T3562 = io_resetCounts ? 4'h0 : counts_584;
  assign T3563 = T10320 & T3564;
  assign T3564 = T76[10'h248:10'h248];
  assign T10930 = reset ? 4'h0 : T3565;
  assign T3565 = T3567 ? T52 : T3566;
  assign T3566 = io_resetCounts ? 4'h0 : counts_585;
  assign T3567 = T10320 & T3568;
  assign T3568 = T76[10'h249:10'h249];
  assign T3569 = T68[1'h0:1'h0];
  assign T3570 = T3579 ? counts_587 : counts_586;
  assign T10931 = reset ? 4'h0 : T3571;
  assign T3571 = T3573 ? T52 : T3572;
  assign T3572 = io_resetCounts ? 4'h0 : counts_586;
  assign T3573 = T10320 & T3574;
  assign T3574 = T76[10'h24a:10'h24a];
  assign T10932 = reset ? 4'h0 : T3575;
  assign T3575 = T3577 ? T52 : T3576;
  assign T3576 = io_resetCounts ? 4'h0 : counts_587;
  assign T3577 = T10320 & T3578;
  assign T3578 = T76[10'h24b:10'h24b];
  assign T3579 = T68[1'h0:1'h0];
  assign T3580 = T68[1'h1:1'h1];
  assign T3581 = T3602 ? T3592 : T3582;
  assign T3582 = T3591 ? counts_589 : counts_588;
  assign T10933 = reset ? 4'h0 : T3583;
  assign T3583 = T3585 ? T52 : T3584;
  assign T3584 = io_resetCounts ? 4'h0 : counts_588;
  assign T3585 = T10320 & T3586;
  assign T3586 = T76[10'h24c:10'h24c];
  assign T10934 = reset ? 4'h0 : T3587;
  assign T3587 = T3589 ? T52 : T3588;
  assign T3588 = io_resetCounts ? 4'h0 : counts_589;
  assign T3589 = T10320 & T3590;
  assign T3590 = T76[10'h24d:10'h24d];
  assign T3591 = T68[1'h0:1'h0];
  assign T3592 = T3601 ? counts_591 : counts_590;
  assign T10935 = reset ? 4'h0 : T3593;
  assign T3593 = T3595 ? T52 : T3594;
  assign T3594 = io_resetCounts ? 4'h0 : counts_590;
  assign T3595 = T10320 & T3596;
  assign T3596 = T76[10'h24e:10'h24e];
  assign T10936 = reset ? 4'h0 : T3597;
  assign T3597 = T3599 ? T52 : T3598;
  assign T3598 = io_resetCounts ? 4'h0 : counts_591;
  assign T3599 = T10320 & T3600;
  assign T3600 = T76[10'h24f:10'h24f];
  assign T3601 = T68[1'h0:1'h0];
  assign T3602 = T68[1'h1:1'h1];
  assign T3603 = T68[2'h2:2'h2];
  assign T3604 = T68[2'h3:2'h3];
  assign T3605 = T3698 ? T3652 : T3606;
  assign T3606 = T3651 ? T3629 : T3607;
  assign T3607 = T3628 ? T3618 : T3608;
  assign T3608 = T3617 ? counts_593 : counts_592;
  assign T10937 = reset ? 4'h0 : T3609;
  assign T3609 = T3611 ? T52 : T3610;
  assign T3610 = io_resetCounts ? 4'h0 : counts_592;
  assign T3611 = T10320 & T3612;
  assign T3612 = T76[10'h250:10'h250];
  assign T10938 = reset ? 4'h0 : T3613;
  assign T3613 = T3615 ? T52 : T3614;
  assign T3614 = io_resetCounts ? 4'h0 : counts_593;
  assign T3615 = T10320 & T3616;
  assign T3616 = T76[10'h251:10'h251];
  assign T3617 = T68[1'h0:1'h0];
  assign T3618 = T3627 ? counts_595 : counts_594;
  assign T10939 = reset ? 4'h0 : T3619;
  assign T3619 = T3621 ? T52 : T3620;
  assign T3620 = io_resetCounts ? 4'h0 : counts_594;
  assign T3621 = T10320 & T3622;
  assign T3622 = T76[10'h252:10'h252];
  assign T10940 = reset ? 4'h0 : T3623;
  assign T3623 = T3625 ? T52 : T3624;
  assign T3624 = io_resetCounts ? 4'h0 : counts_595;
  assign T3625 = T10320 & T3626;
  assign T3626 = T76[10'h253:10'h253];
  assign T3627 = T68[1'h0:1'h0];
  assign T3628 = T68[1'h1:1'h1];
  assign T3629 = T3650 ? T3640 : T3630;
  assign T3630 = T3639 ? counts_597 : counts_596;
  assign T10941 = reset ? 4'h0 : T3631;
  assign T3631 = T3633 ? T52 : T3632;
  assign T3632 = io_resetCounts ? 4'h0 : counts_596;
  assign T3633 = T10320 & T3634;
  assign T3634 = T76[10'h254:10'h254];
  assign T10942 = reset ? 4'h0 : T3635;
  assign T3635 = T3637 ? T52 : T3636;
  assign T3636 = io_resetCounts ? 4'h0 : counts_597;
  assign T3637 = T10320 & T3638;
  assign T3638 = T76[10'h255:10'h255];
  assign T3639 = T68[1'h0:1'h0];
  assign T3640 = T3649 ? counts_599 : counts_598;
  assign T10943 = reset ? 4'h0 : T3641;
  assign T3641 = T3643 ? T52 : T3642;
  assign T3642 = io_resetCounts ? 4'h0 : counts_598;
  assign T3643 = T10320 & T3644;
  assign T3644 = T76[10'h256:10'h256];
  assign T10944 = reset ? 4'h0 : T3645;
  assign T3645 = T3647 ? T52 : T3646;
  assign T3646 = io_resetCounts ? 4'h0 : counts_599;
  assign T3647 = T10320 & T3648;
  assign T3648 = T76[10'h257:10'h257];
  assign T3649 = T68[1'h0:1'h0];
  assign T3650 = T68[1'h1:1'h1];
  assign T3651 = T68[2'h2:2'h2];
  assign T3652 = T3697 ? T3675 : T3653;
  assign T3653 = T3674 ? T3664 : T3654;
  assign T3654 = T3663 ? counts_601 : counts_600;
  assign T10945 = reset ? 4'h0 : T3655;
  assign T3655 = T3657 ? T52 : T3656;
  assign T3656 = io_resetCounts ? 4'h0 : counts_600;
  assign T3657 = T10320 & T3658;
  assign T3658 = T76[10'h258:10'h258];
  assign T10946 = reset ? 4'h0 : T3659;
  assign T3659 = T3661 ? T52 : T3660;
  assign T3660 = io_resetCounts ? 4'h0 : counts_601;
  assign T3661 = T10320 & T3662;
  assign T3662 = T76[10'h259:10'h259];
  assign T3663 = T68[1'h0:1'h0];
  assign T3664 = T3673 ? counts_603 : counts_602;
  assign T10947 = reset ? 4'h0 : T3665;
  assign T3665 = T3667 ? T52 : T3666;
  assign T3666 = io_resetCounts ? 4'h0 : counts_602;
  assign T3667 = T10320 & T3668;
  assign T3668 = T76[10'h25a:10'h25a];
  assign T10948 = reset ? 4'h0 : T3669;
  assign T3669 = T3671 ? T52 : T3670;
  assign T3670 = io_resetCounts ? 4'h0 : counts_603;
  assign T3671 = T10320 & T3672;
  assign T3672 = T76[10'h25b:10'h25b];
  assign T3673 = T68[1'h0:1'h0];
  assign T3674 = T68[1'h1:1'h1];
  assign T3675 = T3696 ? T3686 : T3676;
  assign T3676 = T3685 ? counts_605 : counts_604;
  assign T10949 = reset ? 4'h0 : T3677;
  assign T3677 = T3679 ? T52 : T3678;
  assign T3678 = io_resetCounts ? 4'h0 : counts_604;
  assign T3679 = T10320 & T3680;
  assign T3680 = T76[10'h25c:10'h25c];
  assign T10950 = reset ? 4'h0 : T3681;
  assign T3681 = T3683 ? T52 : T3682;
  assign T3682 = io_resetCounts ? 4'h0 : counts_605;
  assign T3683 = T10320 & T3684;
  assign T3684 = T76[10'h25d:10'h25d];
  assign T3685 = T68[1'h0:1'h0];
  assign T3686 = T3695 ? counts_607 : counts_606;
  assign T10951 = reset ? 4'h0 : T3687;
  assign T3687 = T3689 ? T52 : T3688;
  assign T3688 = io_resetCounts ? 4'h0 : counts_606;
  assign T3689 = T10320 & T3690;
  assign T3690 = T76[10'h25e:10'h25e];
  assign T10952 = reset ? 4'h0 : T3691;
  assign T3691 = T3693 ? T52 : T3692;
  assign T3692 = io_resetCounts ? 4'h0 : counts_607;
  assign T3693 = T10320 & T3694;
  assign T3694 = T76[10'h25f:10'h25f];
  assign T3695 = T68[1'h0:1'h0];
  assign T3696 = T68[1'h1:1'h1];
  assign T3697 = T68[2'h2:2'h2];
  assign T3698 = T68[2'h3:2'h3];
  assign T3699 = T68[3'h4:3'h4];
  assign T3700 = T3889 ? T3795 : T3701;
  assign T3701 = T3794 ? T3748 : T3702;
  assign T3702 = T3747 ? T3725 : T3703;
  assign T3703 = T3724 ? T3714 : T3704;
  assign T3704 = T3713 ? counts_609 : counts_608;
  assign T10953 = reset ? 4'h0 : T3705;
  assign T3705 = T3707 ? T52 : T3706;
  assign T3706 = io_resetCounts ? 4'h0 : counts_608;
  assign T3707 = T10320 & T3708;
  assign T3708 = T76[10'h260:10'h260];
  assign T10954 = reset ? 4'h0 : T3709;
  assign T3709 = T3711 ? T52 : T3710;
  assign T3710 = io_resetCounts ? 4'h0 : counts_609;
  assign T3711 = T10320 & T3712;
  assign T3712 = T76[10'h261:10'h261];
  assign T3713 = T68[1'h0:1'h0];
  assign T3714 = T3723 ? counts_611 : counts_610;
  assign T10955 = reset ? 4'h0 : T3715;
  assign T3715 = T3717 ? T52 : T3716;
  assign T3716 = io_resetCounts ? 4'h0 : counts_610;
  assign T3717 = T10320 & T3718;
  assign T3718 = T76[10'h262:10'h262];
  assign T10956 = reset ? 4'h0 : T3719;
  assign T3719 = T3721 ? T52 : T3720;
  assign T3720 = io_resetCounts ? 4'h0 : counts_611;
  assign T3721 = T10320 & T3722;
  assign T3722 = T76[10'h263:10'h263];
  assign T3723 = T68[1'h0:1'h0];
  assign T3724 = T68[1'h1:1'h1];
  assign T3725 = T3746 ? T3736 : T3726;
  assign T3726 = T3735 ? counts_613 : counts_612;
  assign T10957 = reset ? 4'h0 : T3727;
  assign T3727 = T3729 ? T52 : T3728;
  assign T3728 = io_resetCounts ? 4'h0 : counts_612;
  assign T3729 = T10320 & T3730;
  assign T3730 = T76[10'h264:10'h264];
  assign T10958 = reset ? 4'h0 : T3731;
  assign T3731 = T3733 ? T52 : T3732;
  assign T3732 = io_resetCounts ? 4'h0 : counts_613;
  assign T3733 = T10320 & T3734;
  assign T3734 = T76[10'h265:10'h265];
  assign T3735 = T68[1'h0:1'h0];
  assign T3736 = T3745 ? counts_615 : counts_614;
  assign T10959 = reset ? 4'h0 : T3737;
  assign T3737 = T3739 ? T52 : T3738;
  assign T3738 = io_resetCounts ? 4'h0 : counts_614;
  assign T3739 = T10320 & T3740;
  assign T3740 = T76[10'h266:10'h266];
  assign T10960 = reset ? 4'h0 : T3741;
  assign T3741 = T3743 ? T52 : T3742;
  assign T3742 = io_resetCounts ? 4'h0 : counts_615;
  assign T3743 = T10320 & T3744;
  assign T3744 = T76[10'h267:10'h267];
  assign T3745 = T68[1'h0:1'h0];
  assign T3746 = T68[1'h1:1'h1];
  assign T3747 = T68[2'h2:2'h2];
  assign T3748 = T3793 ? T3771 : T3749;
  assign T3749 = T3770 ? T3760 : T3750;
  assign T3750 = T3759 ? counts_617 : counts_616;
  assign T10961 = reset ? 4'h0 : T3751;
  assign T3751 = T3753 ? T52 : T3752;
  assign T3752 = io_resetCounts ? 4'h0 : counts_616;
  assign T3753 = T10320 & T3754;
  assign T3754 = T76[10'h268:10'h268];
  assign T10962 = reset ? 4'h0 : T3755;
  assign T3755 = T3757 ? T52 : T3756;
  assign T3756 = io_resetCounts ? 4'h0 : counts_617;
  assign T3757 = T10320 & T3758;
  assign T3758 = T76[10'h269:10'h269];
  assign T3759 = T68[1'h0:1'h0];
  assign T3760 = T3769 ? counts_619 : counts_618;
  assign T10963 = reset ? 4'h0 : T3761;
  assign T3761 = T3763 ? T52 : T3762;
  assign T3762 = io_resetCounts ? 4'h0 : counts_618;
  assign T3763 = T10320 & T3764;
  assign T3764 = T76[10'h26a:10'h26a];
  assign T10964 = reset ? 4'h0 : T3765;
  assign T3765 = T3767 ? T52 : T3766;
  assign T3766 = io_resetCounts ? 4'h0 : counts_619;
  assign T3767 = T10320 & T3768;
  assign T3768 = T76[10'h26b:10'h26b];
  assign T3769 = T68[1'h0:1'h0];
  assign T3770 = T68[1'h1:1'h1];
  assign T3771 = T3792 ? T3782 : T3772;
  assign T3772 = T3781 ? counts_621 : counts_620;
  assign T10965 = reset ? 4'h0 : T3773;
  assign T3773 = T3775 ? T52 : T3774;
  assign T3774 = io_resetCounts ? 4'h0 : counts_620;
  assign T3775 = T10320 & T3776;
  assign T3776 = T76[10'h26c:10'h26c];
  assign T10966 = reset ? 4'h0 : T3777;
  assign T3777 = T3779 ? T52 : T3778;
  assign T3778 = io_resetCounts ? 4'h0 : counts_621;
  assign T3779 = T10320 & T3780;
  assign T3780 = T76[10'h26d:10'h26d];
  assign T3781 = T68[1'h0:1'h0];
  assign T3782 = T3791 ? counts_623 : counts_622;
  assign T10967 = reset ? 4'h0 : T3783;
  assign T3783 = T3785 ? T52 : T3784;
  assign T3784 = io_resetCounts ? 4'h0 : counts_622;
  assign T3785 = T10320 & T3786;
  assign T3786 = T76[10'h26e:10'h26e];
  assign T10968 = reset ? 4'h0 : T3787;
  assign T3787 = T3789 ? T52 : T3788;
  assign T3788 = io_resetCounts ? 4'h0 : counts_623;
  assign T3789 = T10320 & T3790;
  assign T3790 = T76[10'h26f:10'h26f];
  assign T3791 = T68[1'h0:1'h0];
  assign T3792 = T68[1'h1:1'h1];
  assign T3793 = T68[2'h2:2'h2];
  assign T3794 = T68[2'h3:2'h3];
  assign T3795 = T3888 ? T3842 : T3796;
  assign T3796 = T3841 ? T3819 : T3797;
  assign T3797 = T3818 ? T3808 : T3798;
  assign T3798 = T3807 ? counts_625 : counts_624;
  assign T10969 = reset ? 4'h0 : T3799;
  assign T3799 = T3801 ? T52 : T3800;
  assign T3800 = io_resetCounts ? 4'h0 : counts_624;
  assign T3801 = T10320 & T3802;
  assign T3802 = T76[10'h270:10'h270];
  assign T10970 = reset ? 4'h0 : T3803;
  assign T3803 = T3805 ? T52 : T3804;
  assign T3804 = io_resetCounts ? 4'h0 : counts_625;
  assign T3805 = T10320 & T3806;
  assign T3806 = T76[10'h271:10'h271];
  assign T3807 = T68[1'h0:1'h0];
  assign T3808 = T3817 ? counts_627 : counts_626;
  assign T10971 = reset ? 4'h0 : T3809;
  assign T3809 = T3811 ? T52 : T3810;
  assign T3810 = io_resetCounts ? 4'h0 : counts_626;
  assign T3811 = T10320 & T3812;
  assign T3812 = T76[10'h272:10'h272];
  assign T10972 = reset ? 4'h0 : T3813;
  assign T3813 = T3815 ? T52 : T3814;
  assign T3814 = io_resetCounts ? 4'h0 : counts_627;
  assign T3815 = T10320 & T3816;
  assign T3816 = T76[10'h273:10'h273];
  assign T3817 = T68[1'h0:1'h0];
  assign T3818 = T68[1'h1:1'h1];
  assign T3819 = T3840 ? T3830 : T3820;
  assign T3820 = T3829 ? counts_629 : counts_628;
  assign T10973 = reset ? 4'h0 : T3821;
  assign T3821 = T3823 ? T52 : T3822;
  assign T3822 = io_resetCounts ? 4'h0 : counts_628;
  assign T3823 = T10320 & T3824;
  assign T3824 = T76[10'h274:10'h274];
  assign T10974 = reset ? 4'h0 : T3825;
  assign T3825 = T3827 ? T52 : T3826;
  assign T3826 = io_resetCounts ? 4'h0 : counts_629;
  assign T3827 = T10320 & T3828;
  assign T3828 = T76[10'h275:10'h275];
  assign T3829 = T68[1'h0:1'h0];
  assign T3830 = T3839 ? counts_631 : counts_630;
  assign T10975 = reset ? 4'h0 : T3831;
  assign T3831 = T3833 ? T52 : T3832;
  assign T3832 = io_resetCounts ? 4'h0 : counts_630;
  assign T3833 = T10320 & T3834;
  assign T3834 = T76[10'h276:10'h276];
  assign T10976 = reset ? 4'h0 : T3835;
  assign T3835 = T3837 ? T52 : T3836;
  assign T3836 = io_resetCounts ? 4'h0 : counts_631;
  assign T3837 = T10320 & T3838;
  assign T3838 = T76[10'h277:10'h277];
  assign T3839 = T68[1'h0:1'h0];
  assign T3840 = T68[1'h1:1'h1];
  assign T3841 = T68[2'h2:2'h2];
  assign T3842 = T3887 ? T3865 : T3843;
  assign T3843 = T3864 ? T3854 : T3844;
  assign T3844 = T3853 ? counts_633 : counts_632;
  assign T10977 = reset ? 4'h0 : T3845;
  assign T3845 = T3847 ? T52 : T3846;
  assign T3846 = io_resetCounts ? 4'h0 : counts_632;
  assign T3847 = T10320 & T3848;
  assign T3848 = T76[10'h278:10'h278];
  assign T10978 = reset ? 4'h0 : T3849;
  assign T3849 = T3851 ? T52 : T3850;
  assign T3850 = io_resetCounts ? 4'h0 : counts_633;
  assign T3851 = T10320 & T3852;
  assign T3852 = T76[10'h279:10'h279];
  assign T3853 = T68[1'h0:1'h0];
  assign T3854 = T3863 ? counts_635 : counts_634;
  assign T10979 = reset ? 4'h0 : T3855;
  assign T3855 = T3857 ? T52 : T3856;
  assign T3856 = io_resetCounts ? 4'h0 : counts_634;
  assign T3857 = T10320 & T3858;
  assign T3858 = T76[10'h27a:10'h27a];
  assign T10980 = reset ? 4'h0 : T3859;
  assign T3859 = T3861 ? T52 : T3860;
  assign T3860 = io_resetCounts ? 4'h0 : counts_635;
  assign T3861 = T10320 & T3862;
  assign T3862 = T76[10'h27b:10'h27b];
  assign T3863 = T68[1'h0:1'h0];
  assign T3864 = T68[1'h1:1'h1];
  assign T3865 = T3886 ? T3876 : T3866;
  assign T3866 = T3875 ? counts_637 : counts_636;
  assign T10981 = reset ? 4'h0 : T3867;
  assign T3867 = T3869 ? T52 : T3868;
  assign T3868 = io_resetCounts ? 4'h0 : counts_636;
  assign T3869 = T10320 & T3870;
  assign T3870 = T76[10'h27c:10'h27c];
  assign T10982 = reset ? 4'h0 : T3871;
  assign T3871 = T3873 ? T52 : T3872;
  assign T3872 = io_resetCounts ? 4'h0 : counts_637;
  assign T3873 = T10320 & T3874;
  assign T3874 = T76[10'h27d:10'h27d];
  assign T3875 = T68[1'h0:1'h0];
  assign T3876 = T3885 ? counts_639 : counts_638;
  assign T10983 = reset ? 4'h0 : T3877;
  assign T3877 = T3879 ? T52 : T3878;
  assign T3878 = io_resetCounts ? 4'h0 : counts_638;
  assign T3879 = T10320 & T3880;
  assign T3880 = T76[10'h27e:10'h27e];
  assign T10984 = reset ? 4'h0 : T3881;
  assign T3881 = T3883 ? T52 : T3882;
  assign T3882 = io_resetCounts ? 4'h0 : counts_639;
  assign T3883 = T10320 & T3884;
  assign T3884 = T76[10'h27f:10'h27f];
  assign T3885 = T68[1'h0:1'h0];
  assign T3886 = T68[1'h1:1'h1];
  assign T3887 = T68[2'h2:2'h2];
  assign T3888 = T68[2'h3:2'h3];
  assign T3889 = T68[3'h4:3'h4];
  assign T3890 = T68[3'h5:3'h5];
  assign T3891 = T68[3'h6:3'h6];
  assign T3892 = T4657 ? T4275 : T3893;
  assign T3893 = T4274 ? T4084 : T3894;
  assign T3894 = T4083 ? T3989 : T3895;
  assign T3895 = T3988 ? T3942 : T3896;
  assign T3896 = T3941 ? T3919 : T3897;
  assign T3897 = T3918 ? T3908 : T3898;
  assign T3898 = T3907 ? counts_641 : counts_640;
  assign T10985 = reset ? 4'h0 : T3899;
  assign T3899 = T3901 ? T52 : T3900;
  assign T3900 = io_resetCounts ? 4'h0 : counts_640;
  assign T3901 = T10320 & T3902;
  assign T3902 = T76[10'h280:10'h280];
  assign T10986 = reset ? 4'h0 : T3903;
  assign T3903 = T3905 ? T52 : T3904;
  assign T3904 = io_resetCounts ? 4'h0 : counts_641;
  assign T3905 = T10320 & T3906;
  assign T3906 = T76[10'h281:10'h281];
  assign T3907 = T68[1'h0:1'h0];
  assign T3908 = T3917 ? counts_643 : counts_642;
  assign T10987 = reset ? 4'h0 : T3909;
  assign T3909 = T3911 ? T52 : T3910;
  assign T3910 = io_resetCounts ? 4'h0 : counts_642;
  assign T3911 = T10320 & T3912;
  assign T3912 = T76[10'h282:10'h282];
  assign T10988 = reset ? 4'h0 : T3913;
  assign T3913 = T3915 ? T52 : T3914;
  assign T3914 = io_resetCounts ? 4'h0 : counts_643;
  assign T3915 = T10320 & T3916;
  assign T3916 = T76[10'h283:10'h283];
  assign T3917 = T68[1'h0:1'h0];
  assign T3918 = T68[1'h1:1'h1];
  assign T3919 = T3940 ? T3930 : T3920;
  assign T3920 = T3929 ? counts_645 : counts_644;
  assign T10989 = reset ? 4'h0 : T3921;
  assign T3921 = T3923 ? T52 : T3922;
  assign T3922 = io_resetCounts ? 4'h0 : counts_644;
  assign T3923 = T10320 & T3924;
  assign T3924 = T76[10'h284:10'h284];
  assign T10990 = reset ? 4'h0 : T3925;
  assign T3925 = T3927 ? T52 : T3926;
  assign T3926 = io_resetCounts ? 4'h0 : counts_645;
  assign T3927 = T10320 & T3928;
  assign T3928 = T76[10'h285:10'h285];
  assign T3929 = T68[1'h0:1'h0];
  assign T3930 = T3939 ? counts_647 : counts_646;
  assign T10991 = reset ? 4'h0 : T3931;
  assign T3931 = T3933 ? T52 : T3932;
  assign T3932 = io_resetCounts ? 4'h0 : counts_646;
  assign T3933 = T10320 & T3934;
  assign T3934 = T76[10'h286:10'h286];
  assign T10992 = reset ? 4'h0 : T3935;
  assign T3935 = T3937 ? T52 : T3936;
  assign T3936 = io_resetCounts ? 4'h0 : counts_647;
  assign T3937 = T10320 & T3938;
  assign T3938 = T76[10'h287:10'h287];
  assign T3939 = T68[1'h0:1'h0];
  assign T3940 = T68[1'h1:1'h1];
  assign T3941 = T68[2'h2:2'h2];
  assign T3942 = T3987 ? T3965 : T3943;
  assign T3943 = T3964 ? T3954 : T3944;
  assign T3944 = T3953 ? counts_649 : counts_648;
  assign T10993 = reset ? 4'h0 : T3945;
  assign T3945 = T3947 ? T52 : T3946;
  assign T3946 = io_resetCounts ? 4'h0 : counts_648;
  assign T3947 = T10320 & T3948;
  assign T3948 = T76[10'h288:10'h288];
  assign T10994 = reset ? 4'h0 : T3949;
  assign T3949 = T3951 ? T52 : T3950;
  assign T3950 = io_resetCounts ? 4'h0 : counts_649;
  assign T3951 = T10320 & T3952;
  assign T3952 = T76[10'h289:10'h289];
  assign T3953 = T68[1'h0:1'h0];
  assign T3954 = T3963 ? counts_651 : counts_650;
  assign T10995 = reset ? 4'h0 : T3955;
  assign T3955 = T3957 ? T52 : T3956;
  assign T3956 = io_resetCounts ? 4'h0 : counts_650;
  assign T3957 = T10320 & T3958;
  assign T3958 = T76[10'h28a:10'h28a];
  assign T10996 = reset ? 4'h0 : T3959;
  assign T3959 = T3961 ? T52 : T3960;
  assign T3960 = io_resetCounts ? 4'h0 : counts_651;
  assign T3961 = T10320 & T3962;
  assign T3962 = T76[10'h28b:10'h28b];
  assign T3963 = T68[1'h0:1'h0];
  assign T3964 = T68[1'h1:1'h1];
  assign T3965 = T3986 ? T3976 : T3966;
  assign T3966 = T3975 ? counts_653 : counts_652;
  assign T10997 = reset ? 4'h0 : T3967;
  assign T3967 = T3969 ? T52 : T3968;
  assign T3968 = io_resetCounts ? 4'h0 : counts_652;
  assign T3969 = T10320 & T3970;
  assign T3970 = T76[10'h28c:10'h28c];
  assign T10998 = reset ? 4'h0 : T3971;
  assign T3971 = T3973 ? T52 : T3972;
  assign T3972 = io_resetCounts ? 4'h0 : counts_653;
  assign T3973 = T10320 & T3974;
  assign T3974 = T76[10'h28d:10'h28d];
  assign T3975 = T68[1'h0:1'h0];
  assign T3976 = T3985 ? counts_655 : counts_654;
  assign T10999 = reset ? 4'h0 : T3977;
  assign T3977 = T3979 ? T52 : T3978;
  assign T3978 = io_resetCounts ? 4'h0 : counts_654;
  assign T3979 = T10320 & T3980;
  assign T3980 = T76[10'h28e:10'h28e];
  assign T11000 = reset ? 4'h0 : T3981;
  assign T3981 = T3983 ? T52 : T3982;
  assign T3982 = io_resetCounts ? 4'h0 : counts_655;
  assign T3983 = T10320 & T3984;
  assign T3984 = T76[10'h28f:10'h28f];
  assign T3985 = T68[1'h0:1'h0];
  assign T3986 = T68[1'h1:1'h1];
  assign T3987 = T68[2'h2:2'h2];
  assign T3988 = T68[2'h3:2'h3];
  assign T3989 = T4082 ? T4036 : T3990;
  assign T3990 = T4035 ? T4013 : T3991;
  assign T3991 = T4012 ? T4002 : T3992;
  assign T3992 = T4001 ? counts_657 : counts_656;
  assign T11001 = reset ? 4'h0 : T3993;
  assign T3993 = T3995 ? T52 : T3994;
  assign T3994 = io_resetCounts ? 4'h0 : counts_656;
  assign T3995 = T10320 & T3996;
  assign T3996 = T76[10'h290:10'h290];
  assign T11002 = reset ? 4'h0 : T3997;
  assign T3997 = T3999 ? T52 : T3998;
  assign T3998 = io_resetCounts ? 4'h0 : counts_657;
  assign T3999 = T10320 & T4000;
  assign T4000 = T76[10'h291:10'h291];
  assign T4001 = T68[1'h0:1'h0];
  assign T4002 = T4011 ? counts_659 : counts_658;
  assign T11003 = reset ? 4'h0 : T4003;
  assign T4003 = T4005 ? T52 : T4004;
  assign T4004 = io_resetCounts ? 4'h0 : counts_658;
  assign T4005 = T10320 & T4006;
  assign T4006 = T76[10'h292:10'h292];
  assign T11004 = reset ? 4'h0 : T4007;
  assign T4007 = T4009 ? T52 : T4008;
  assign T4008 = io_resetCounts ? 4'h0 : counts_659;
  assign T4009 = T10320 & T4010;
  assign T4010 = T76[10'h293:10'h293];
  assign T4011 = T68[1'h0:1'h0];
  assign T4012 = T68[1'h1:1'h1];
  assign T4013 = T4034 ? T4024 : T4014;
  assign T4014 = T4023 ? counts_661 : counts_660;
  assign T11005 = reset ? 4'h0 : T4015;
  assign T4015 = T4017 ? T52 : T4016;
  assign T4016 = io_resetCounts ? 4'h0 : counts_660;
  assign T4017 = T10320 & T4018;
  assign T4018 = T76[10'h294:10'h294];
  assign T11006 = reset ? 4'h0 : T4019;
  assign T4019 = T4021 ? T52 : T4020;
  assign T4020 = io_resetCounts ? 4'h0 : counts_661;
  assign T4021 = T10320 & T4022;
  assign T4022 = T76[10'h295:10'h295];
  assign T4023 = T68[1'h0:1'h0];
  assign T4024 = T4033 ? counts_663 : counts_662;
  assign T11007 = reset ? 4'h0 : T4025;
  assign T4025 = T4027 ? T52 : T4026;
  assign T4026 = io_resetCounts ? 4'h0 : counts_662;
  assign T4027 = T10320 & T4028;
  assign T4028 = T76[10'h296:10'h296];
  assign T11008 = reset ? 4'h0 : T4029;
  assign T4029 = T4031 ? T52 : T4030;
  assign T4030 = io_resetCounts ? 4'h0 : counts_663;
  assign T4031 = T10320 & T4032;
  assign T4032 = T76[10'h297:10'h297];
  assign T4033 = T68[1'h0:1'h0];
  assign T4034 = T68[1'h1:1'h1];
  assign T4035 = T68[2'h2:2'h2];
  assign T4036 = T4081 ? T4059 : T4037;
  assign T4037 = T4058 ? T4048 : T4038;
  assign T4038 = T4047 ? counts_665 : counts_664;
  assign T11009 = reset ? 4'h0 : T4039;
  assign T4039 = T4041 ? T52 : T4040;
  assign T4040 = io_resetCounts ? 4'h0 : counts_664;
  assign T4041 = T10320 & T4042;
  assign T4042 = T76[10'h298:10'h298];
  assign T11010 = reset ? 4'h0 : T4043;
  assign T4043 = T4045 ? T52 : T4044;
  assign T4044 = io_resetCounts ? 4'h0 : counts_665;
  assign T4045 = T10320 & T4046;
  assign T4046 = T76[10'h299:10'h299];
  assign T4047 = T68[1'h0:1'h0];
  assign T4048 = T4057 ? counts_667 : counts_666;
  assign T11011 = reset ? 4'h0 : T4049;
  assign T4049 = T4051 ? T52 : T4050;
  assign T4050 = io_resetCounts ? 4'h0 : counts_666;
  assign T4051 = T10320 & T4052;
  assign T4052 = T76[10'h29a:10'h29a];
  assign T11012 = reset ? 4'h0 : T4053;
  assign T4053 = T4055 ? T52 : T4054;
  assign T4054 = io_resetCounts ? 4'h0 : counts_667;
  assign T4055 = T10320 & T4056;
  assign T4056 = T76[10'h29b:10'h29b];
  assign T4057 = T68[1'h0:1'h0];
  assign T4058 = T68[1'h1:1'h1];
  assign T4059 = T4080 ? T4070 : T4060;
  assign T4060 = T4069 ? counts_669 : counts_668;
  assign T11013 = reset ? 4'h0 : T4061;
  assign T4061 = T4063 ? T52 : T4062;
  assign T4062 = io_resetCounts ? 4'h0 : counts_668;
  assign T4063 = T10320 & T4064;
  assign T4064 = T76[10'h29c:10'h29c];
  assign T11014 = reset ? 4'h0 : T4065;
  assign T4065 = T4067 ? T52 : T4066;
  assign T4066 = io_resetCounts ? 4'h0 : counts_669;
  assign T4067 = T10320 & T4068;
  assign T4068 = T76[10'h29d:10'h29d];
  assign T4069 = T68[1'h0:1'h0];
  assign T4070 = T4079 ? counts_671 : counts_670;
  assign T11015 = reset ? 4'h0 : T4071;
  assign T4071 = T4073 ? T52 : T4072;
  assign T4072 = io_resetCounts ? 4'h0 : counts_670;
  assign T4073 = T10320 & T4074;
  assign T4074 = T76[10'h29e:10'h29e];
  assign T11016 = reset ? 4'h0 : T4075;
  assign T4075 = T4077 ? T52 : T4076;
  assign T4076 = io_resetCounts ? 4'h0 : counts_671;
  assign T4077 = T10320 & T4078;
  assign T4078 = T76[10'h29f:10'h29f];
  assign T4079 = T68[1'h0:1'h0];
  assign T4080 = T68[1'h1:1'h1];
  assign T4081 = T68[2'h2:2'h2];
  assign T4082 = T68[2'h3:2'h3];
  assign T4083 = T68[3'h4:3'h4];
  assign T4084 = T4273 ? T4179 : T4085;
  assign T4085 = T4178 ? T4132 : T4086;
  assign T4086 = T4131 ? T4109 : T4087;
  assign T4087 = T4108 ? T4098 : T4088;
  assign T4088 = T4097 ? counts_673 : counts_672;
  assign T11017 = reset ? 4'h0 : T4089;
  assign T4089 = T4091 ? T52 : T4090;
  assign T4090 = io_resetCounts ? 4'h0 : counts_672;
  assign T4091 = T10320 & T4092;
  assign T4092 = T76[10'h2a0:10'h2a0];
  assign T11018 = reset ? 4'h0 : T4093;
  assign T4093 = T4095 ? T52 : T4094;
  assign T4094 = io_resetCounts ? 4'h0 : counts_673;
  assign T4095 = T10320 & T4096;
  assign T4096 = T76[10'h2a1:10'h2a1];
  assign T4097 = T68[1'h0:1'h0];
  assign T4098 = T4107 ? counts_675 : counts_674;
  assign T11019 = reset ? 4'h0 : T4099;
  assign T4099 = T4101 ? T52 : T4100;
  assign T4100 = io_resetCounts ? 4'h0 : counts_674;
  assign T4101 = T10320 & T4102;
  assign T4102 = T76[10'h2a2:10'h2a2];
  assign T11020 = reset ? 4'h0 : T4103;
  assign T4103 = T4105 ? T52 : T4104;
  assign T4104 = io_resetCounts ? 4'h0 : counts_675;
  assign T4105 = T10320 & T4106;
  assign T4106 = T76[10'h2a3:10'h2a3];
  assign T4107 = T68[1'h0:1'h0];
  assign T4108 = T68[1'h1:1'h1];
  assign T4109 = T4130 ? T4120 : T4110;
  assign T4110 = T4119 ? counts_677 : counts_676;
  assign T11021 = reset ? 4'h0 : T4111;
  assign T4111 = T4113 ? T52 : T4112;
  assign T4112 = io_resetCounts ? 4'h0 : counts_676;
  assign T4113 = T10320 & T4114;
  assign T4114 = T76[10'h2a4:10'h2a4];
  assign T11022 = reset ? 4'h0 : T4115;
  assign T4115 = T4117 ? T52 : T4116;
  assign T4116 = io_resetCounts ? 4'h0 : counts_677;
  assign T4117 = T10320 & T4118;
  assign T4118 = T76[10'h2a5:10'h2a5];
  assign T4119 = T68[1'h0:1'h0];
  assign T4120 = T4129 ? counts_679 : counts_678;
  assign T11023 = reset ? 4'h0 : T4121;
  assign T4121 = T4123 ? T52 : T4122;
  assign T4122 = io_resetCounts ? 4'h0 : counts_678;
  assign T4123 = T10320 & T4124;
  assign T4124 = T76[10'h2a6:10'h2a6];
  assign T11024 = reset ? 4'h0 : T4125;
  assign T4125 = T4127 ? T52 : T4126;
  assign T4126 = io_resetCounts ? 4'h0 : counts_679;
  assign T4127 = T10320 & T4128;
  assign T4128 = T76[10'h2a7:10'h2a7];
  assign T4129 = T68[1'h0:1'h0];
  assign T4130 = T68[1'h1:1'h1];
  assign T4131 = T68[2'h2:2'h2];
  assign T4132 = T4177 ? T4155 : T4133;
  assign T4133 = T4154 ? T4144 : T4134;
  assign T4134 = T4143 ? counts_681 : counts_680;
  assign T11025 = reset ? 4'h0 : T4135;
  assign T4135 = T4137 ? T52 : T4136;
  assign T4136 = io_resetCounts ? 4'h0 : counts_680;
  assign T4137 = T10320 & T4138;
  assign T4138 = T76[10'h2a8:10'h2a8];
  assign T11026 = reset ? 4'h0 : T4139;
  assign T4139 = T4141 ? T52 : T4140;
  assign T4140 = io_resetCounts ? 4'h0 : counts_681;
  assign T4141 = T10320 & T4142;
  assign T4142 = T76[10'h2a9:10'h2a9];
  assign T4143 = T68[1'h0:1'h0];
  assign T4144 = T4153 ? counts_683 : counts_682;
  assign T11027 = reset ? 4'h0 : T4145;
  assign T4145 = T4147 ? T52 : T4146;
  assign T4146 = io_resetCounts ? 4'h0 : counts_682;
  assign T4147 = T10320 & T4148;
  assign T4148 = T76[10'h2aa:10'h2aa];
  assign T11028 = reset ? 4'h0 : T4149;
  assign T4149 = T4151 ? T52 : T4150;
  assign T4150 = io_resetCounts ? 4'h0 : counts_683;
  assign T4151 = T10320 & T4152;
  assign T4152 = T76[10'h2ab:10'h2ab];
  assign T4153 = T68[1'h0:1'h0];
  assign T4154 = T68[1'h1:1'h1];
  assign T4155 = T4176 ? T4166 : T4156;
  assign T4156 = T4165 ? counts_685 : counts_684;
  assign T11029 = reset ? 4'h0 : T4157;
  assign T4157 = T4159 ? T52 : T4158;
  assign T4158 = io_resetCounts ? 4'h0 : counts_684;
  assign T4159 = T10320 & T4160;
  assign T4160 = T76[10'h2ac:10'h2ac];
  assign T11030 = reset ? 4'h0 : T4161;
  assign T4161 = T4163 ? T52 : T4162;
  assign T4162 = io_resetCounts ? 4'h0 : counts_685;
  assign T4163 = T10320 & T4164;
  assign T4164 = T76[10'h2ad:10'h2ad];
  assign T4165 = T68[1'h0:1'h0];
  assign T4166 = T4175 ? counts_687 : counts_686;
  assign T11031 = reset ? 4'h0 : T4167;
  assign T4167 = T4169 ? T52 : T4168;
  assign T4168 = io_resetCounts ? 4'h0 : counts_686;
  assign T4169 = T10320 & T4170;
  assign T4170 = T76[10'h2ae:10'h2ae];
  assign T11032 = reset ? 4'h0 : T4171;
  assign T4171 = T4173 ? T52 : T4172;
  assign T4172 = io_resetCounts ? 4'h0 : counts_687;
  assign T4173 = T10320 & T4174;
  assign T4174 = T76[10'h2af:10'h2af];
  assign T4175 = T68[1'h0:1'h0];
  assign T4176 = T68[1'h1:1'h1];
  assign T4177 = T68[2'h2:2'h2];
  assign T4178 = T68[2'h3:2'h3];
  assign T4179 = T4272 ? T4226 : T4180;
  assign T4180 = T4225 ? T4203 : T4181;
  assign T4181 = T4202 ? T4192 : T4182;
  assign T4182 = T4191 ? counts_689 : counts_688;
  assign T11033 = reset ? 4'h0 : T4183;
  assign T4183 = T4185 ? T52 : T4184;
  assign T4184 = io_resetCounts ? 4'h0 : counts_688;
  assign T4185 = T10320 & T4186;
  assign T4186 = T76[10'h2b0:10'h2b0];
  assign T11034 = reset ? 4'h0 : T4187;
  assign T4187 = T4189 ? T52 : T4188;
  assign T4188 = io_resetCounts ? 4'h0 : counts_689;
  assign T4189 = T10320 & T4190;
  assign T4190 = T76[10'h2b1:10'h2b1];
  assign T4191 = T68[1'h0:1'h0];
  assign T4192 = T4201 ? counts_691 : counts_690;
  assign T11035 = reset ? 4'h0 : T4193;
  assign T4193 = T4195 ? T52 : T4194;
  assign T4194 = io_resetCounts ? 4'h0 : counts_690;
  assign T4195 = T10320 & T4196;
  assign T4196 = T76[10'h2b2:10'h2b2];
  assign T11036 = reset ? 4'h0 : T4197;
  assign T4197 = T4199 ? T52 : T4198;
  assign T4198 = io_resetCounts ? 4'h0 : counts_691;
  assign T4199 = T10320 & T4200;
  assign T4200 = T76[10'h2b3:10'h2b3];
  assign T4201 = T68[1'h0:1'h0];
  assign T4202 = T68[1'h1:1'h1];
  assign T4203 = T4224 ? T4214 : T4204;
  assign T4204 = T4213 ? counts_693 : counts_692;
  assign T11037 = reset ? 4'h0 : T4205;
  assign T4205 = T4207 ? T52 : T4206;
  assign T4206 = io_resetCounts ? 4'h0 : counts_692;
  assign T4207 = T10320 & T4208;
  assign T4208 = T76[10'h2b4:10'h2b4];
  assign T11038 = reset ? 4'h0 : T4209;
  assign T4209 = T4211 ? T52 : T4210;
  assign T4210 = io_resetCounts ? 4'h0 : counts_693;
  assign T4211 = T10320 & T4212;
  assign T4212 = T76[10'h2b5:10'h2b5];
  assign T4213 = T68[1'h0:1'h0];
  assign T4214 = T4223 ? counts_695 : counts_694;
  assign T11039 = reset ? 4'h0 : T4215;
  assign T4215 = T4217 ? T52 : T4216;
  assign T4216 = io_resetCounts ? 4'h0 : counts_694;
  assign T4217 = T10320 & T4218;
  assign T4218 = T76[10'h2b6:10'h2b6];
  assign T11040 = reset ? 4'h0 : T4219;
  assign T4219 = T4221 ? T52 : T4220;
  assign T4220 = io_resetCounts ? 4'h0 : counts_695;
  assign T4221 = T10320 & T4222;
  assign T4222 = T76[10'h2b7:10'h2b7];
  assign T4223 = T68[1'h0:1'h0];
  assign T4224 = T68[1'h1:1'h1];
  assign T4225 = T68[2'h2:2'h2];
  assign T4226 = T4271 ? T4249 : T4227;
  assign T4227 = T4248 ? T4238 : T4228;
  assign T4228 = T4237 ? counts_697 : counts_696;
  assign T11041 = reset ? 4'h0 : T4229;
  assign T4229 = T4231 ? T52 : T4230;
  assign T4230 = io_resetCounts ? 4'h0 : counts_696;
  assign T4231 = T10320 & T4232;
  assign T4232 = T76[10'h2b8:10'h2b8];
  assign T11042 = reset ? 4'h0 : T4233;
  assign T4233 = T4235 ? T52 : T4234;
  assign T4234 = io_resetCounts ? 4'h0 : counts_697;
  assign T4235 = T10320 & T4236;
  assign T4236 = T76[10'h2b9:10'h2b9];
  assign T4237 = T68[1'h0:1'h0];
  assign T4238 = T4247 ? counts_699 : counts_698;
  assign T11043 = reset ? 4'h0 : T4239;
  assign T4239 = T4241 ? T52 : T4240;
  assign T4240 = io_resetCounts ? 4'h0 : counts_698;
  assign T4241 = T10320 & T4242;
  assign T4242 = T76[10'h2ba:10'h2ba];
  assign T11044 = reset ? 4'h0 : T4243;
  assign T4243 = T4245 ? T52 : T4244;
  assign T4244 = io_resetCounts ? 4'h0 : counts_699;
  assign T4245 = T10320 & T4246;
  assign T4246 = T76[10'h2bb:10'h2bb];
  assign T4247 = T68[1'h0:1'h0];
  assign T4248 = T68[1'h1:1'h1];
  assign T4249 = T4270 ? T4260 : T4250;
  assign T4250 = T4259 ? counts_701 : counts_700;
  assign T11045 = reset ? 4'h0 : T4251;
  assign T4251 = T4253 ? T52 : T4252;
  assign T4252 = io_resetCounts ? 4'h0 : counts_700;
  assign T4253 = T10320 & T4254;
  assign T4254 = T76[10'h2bc:10'h2bc];
  assign T11046 = reset ? 4'h0 : T4255;
  assign T4255 = T4257 ? T52 : T4256;
  assign T4256 = io_resetCounts ? 4'h0 : counts_701;
  assign T4257 = T10320 & T4258;
  assign T4258 = T76[10'h2bd:10'h2bd];
  assign T4259 = T68[1'h0:1'h0];
  assign T4260 = T4269 ? counts_703 : counts_702;
  assign T11047 = reset ? 4'h0 : T4261;
  assign T4261 = T4263 ? T52 : T4262;
  assign T4262 = io_resetCounts ? 4'h0 : counts_702;
  assign T4263 = T10320 & T4264;
  assign T4264 = T76[10'h2be:10'h2be];
  assign T11048 = reset ? 4'h0 : T4265;
  assign T4265 = T4267 ? T52 : T4266;
  assign T4266 = io_resetCounts ? 4'h0 : counts_703;
  assign T4267 = T10320 & T4268;
  assign T4268 = T76[10'h2bf:10'h2bf];
  assign T4269 = T68[1'h0:1'h0];
  assign T4270 = T68[1'h1:1'h1];
  assign T4271 = T68[2'h2:2'h2];
  assign T4272 = T68[2'h3:2'h3];
  assign T4273 = T68[3'h4:3'h4];
  assign T4274 = T68[3'h5:3'h5];
  assign T4275 = T4656 ? T4466 : T4276;
  assign T4276 = T4465 ? T4371 : T4277;
  assign T4277 = T4370 ? T4324 : T4278;
  assign T4278 = T4323 ? T4301 : T4279;
  assign T4279 = T4300 ? T4290 : T4280;
  assign T4280 = T4289 ? counts_705 : counts_704;
  assign T11049 = reset ? 4'h0 : T4281;
  assign T4281 = T4283 ? T52 : T4282;
  assign T4282 = io_resetCounts ? 4'h0 : counts_704;
  assign T4283 = T10320 & T4284;
  assign T4284 = T76[10'h2c0:10'h2c0];
  assign T11050 = reset ? 4'h0 : T4285;
  assign T4285 = T4287 ? T52 : T4286;
  assign T4286 = io_resetCounts ? 4'h0 : counts_705;
  assign T4287 = T10320 & T4288;
  assign T4288 = T76[10'h2c1:10'h2c1];
  assign T4289 = T68[1'h0:1'h0];
  assign T4290 = T4299 ? counts_707 : counts_706;
  assign T11051 = reset ? 4'h0 : T4291;
  assign T4291 = T4293 ? T52 : T4292;
  assign T4292 = io_resetCounts ? 4'h0 : counts_706;
  assign T4293 = T10320 & T4294;
  assign T4294 = T76[10'h2c2:10'h2c2];
  assign T11052 = reset ? 4'h0 : T4295;
  assign T4295 = T4297 ? T52 : T4296;
  assign T4296 = io_resetCounts ? 4'h0 : counts_707;
  assign T4297 = T10320 & T4298;
  assign T4298 = T76[10'h2c3:10'h2c3];
  assign T4299 = T68[1'h0:1'h0];
  assign T4300 = T68[1'h1:1'h1];
  assign T4301 = T4322 ? T4312 : T4302;
  assign T4302 = T4311 ? counts_709 : counts_708;
  assign T11053 = reset ? 4'h0 : T4303;
  assign T4303 = T4305 ? T52 : T4304;
  assign T4304 = io_resetCounts ? 4'h0 : counts_708;
  assign T4305 = T10320 & T4306;
  assign T4306 = T76[10'h2c4:10'h2c4];
  assign T11054 = reset ? 4'h0 : T4307;
  assign T4307 = T4309 ? T52 : T4308;
  assign T4308 = io_resetCounts ? 4'h0 : counts_709;
  assign T4309 = T10320 & T4310;
  assign T4310 = T76[10'h2c5:10'h2c5];
  assign T4311 = T68[1'h0:1'h0];
  assign T4312 = T4321 ? counts_711 : counts_710;
  assign T11055 = reset ? 4'h0 : T4313;
  assign T4313 = T4315 ? T52 : T4314;
  assign T4314 = io_resetCounts ? 4'h0 : counts_710;
  assign T4315 = T10320 & T4316;
  assign T4316 = T76[10'h2c6:10'h2c6];
  assign T11056 = reset ? 4'h0 : T4317;
  assign T4317 = T4319 ? T52 : T4318;
  assign T4318 = io_resetCounts ? 4'h0 : counts_711;
  assign T4319 = T10320 & T4320;
  assign T4320 = T76[10'h2c7:10'h2c7];
  assign T4321 = T68[1'h0:1'h0];
  assign T4322 = T68[1'h1:1'h1];
  assign T4323 = T68[2'h2:2'h2];
  assign T4324 = T4369 ? T4347 : T4325;
  assign T4325 = T4346 ? T4336 : T4326;
  assign T4326 = T4335 ? counts_713 : counts_712;
  assign T11057 = reset ? 4'h0 : T4327;
  assign T4327 = T4329 ? T52 : T4328;
  assign T4328 = io_resetCounts ? 4'h0 : counts_712;
  assign T4329 = T10320 & T4330;
  assign T4330 = T76[10'h2c8:10'h2c8];
  assign T11058 = reset ? 4'h0 : T4331;
  assign T4331 = T4333 ? T52 : T4332;
  assign T4332 = io_resetCounts ? 4'h0 : counts_713;
  assign T4333 = T10320 & T4334;
  assign T4334 = T76[10'h2c9:10'h2c9];
  assign T4335 = T68[1'h0:1'h0];
  assign T4336 = T4345 ? counts_715 : counts_714;
  assign T11059 = reset ? 4'h0 : T4337;
  assign T4337 = T4339 ? T52 : T4338;
  assign T4338 = io_resetCounts ? 4'h0 : counts_714;
  assign T4339 = T10320 & T4340;
  assign T4340 = T76[10'h2ca:10'h2ca];
  assign T11060 = reset ? 4'h0 : T4341;
  assign T4341 = T4343 ? T52 : T4342;
  assign T4342 = io_resetCounts ? 4'h0 : counts_715;
  assign T4343 = T10320 & T4344;
  assign T4344 = T76[10'h2cb:10'h2cb];
  assign T4345 = T68[1'h0:1'h0];
  assign T4346 = T68[1'h1:1'h1];
  assign T4347 = T4368 ? T4358 : T4348;
  assign T4348 = T4357 ? counts_717 : counts_716;
  assign T11061 = reset ? 4'h0 : T4349;
  assign T4349 = T4351 ? T52 : T4350;
  assign T4350 = io_resetCounts ? 4'h0 : counts_716;
  assign T4351 = T10320 & T4352;
  assign T4352 = T76[10'h2cc:10'h2cc];
  assign T11062 = reset ? 4'h0 : T4353;
  assign T4353 = T4355 ? T52 : T4354;
  assign T4354 = io_resetCounts ? 4'h0 : counts_717;
  assign T4355 = T10320 & T4356;
  assign T4356 = T76[10'h2cd:10'h2cd];
  assign T4357 = T68[1'h0:1'h0];
  assign T4358 = T4367 ? counts_719 : counts_718;
  assign T11063 = reset ? 4'h0 : T4359;
  assign T4359 = T4361 ? T52 : T4360;
  assign T4360 = io_resetCounts ? 4'h0 : counts_718;
  assign T4361 = T10320 & T4362;
  assign T4362 = T76[10'h2ce:10'h2ce];
  assign T11064 = reset ? 4'h0 : T4363;
  assign T4363 = T4365 ? T52 : T4364;
  assign T4364 = io_resetCounts ? 4'h0 : counts_719;
  assign T4365 = T10320 & T4366;
  assign T4366 = T76[10'h2cf:10'h2cf];
  assign T4367 = T68[1'h0:1'h0];
  assign T4368 = T68[1'h1:1'h1];
  assign T4369 = T68[2'h2:2'h2];
  assign T4370 = T68[2'h3:2'h3];
  assign T4371 = T4464 ? T4418 : T4372;
  assign T4372 = T4417 ? T4395 : T4373;
  assign T4373 = T4394 ? T4384 : T4374;
  assign T4374 = T4383 ? counts_721 : counts_720;
  assign T11065 = reset ? 4'h0 : T4375;
  assign T4375 = T4377 ? T52 : T4376;
  assign T4376 = io_resetCounts ? 4'h0 : counts_720;
  assign T4377 = T10320 & T4378;
  assign T4378 = T76[10'h2d0:10'h2d0];
  assign T11066 = reset ? 4'h0 : T4379;
  assign T4379 = T4381 ? T52 : T4380;
  assign T4380 = io_resetCounts ? 4'h0 : counts_721;
  assign T4381 = T10320 & T4382;
  assign T4382 = T76[10'h2d1:10'h2d1];
  assign T4383 = T68[1'h0:1'h0];
  assign T4384 = T4393 ? counts_723 : counts_722;
  assign T11067 = reset ? 4'h0 : T4385;
  assign T4385 = T4387 ? T52 : T4386;
  assign T4386 = io_resetCounts ? 4'h0 : counts_722;
  assign T4387 = T10320 & T4388;
  assign T4388 = T76[10'h2d2:10'h2d2];
  assign T11068 = reset ? 4'h0 : T4389;
  assign T4389 = T4391 ? T52 : T4390;
  assign T4390 = io_resetCounts ? 4'h0 : counts_723;
  assign T4391 = T10320 & T4392;
  assign T4392 = T76[10'h2d3:10'h2d3];
  assign T4393 = T68[1'h0:1'h0];
  assign T4394 = T68[1'h1:1'h1];
  assign T4395 = T4416 ? T4406 : T4396;
  assign T4396 = T4405 ? counts_725 : counts_724;
  assign T11069 = reset ? 4'h0 : T4397;
  assign T4397 = T4399 ? T52 : T4398;
  assign T4398 = io_resetCounts ? 4'h0 : counts_724;
  assign T4399 = T10320 & T4400;
  assign T4400 = T76[10'h2d4:10'h2d4];
  assign T11070 = reset ? 4'h0 : T4401;
  assign T4401 = T4403 ? T52 : T4402;
  assign T4402 = io_resetCounts ? 4'h0 : counts_725;
  assign T4403 = T10320 & T4404;
  assign T4404 = T76[10'h2d5:10'h2d5];
  assign T4405 = T68[1'h0:1'h0];
  assign T4406 = T4415 ? counts_727 : counts_726;
  assign T11071 = reset ? 4'h0 : T4407;
  assign T4407 = T4409 ? T52 : T4408;
  assign T4408 = io_resetCounts ? 4'h0 : counts_726;
  assign T4409 = T10320 & T4410;
  assign T4410 = T76[10'h2d6:10'h2d6];
  assign T11072 = reset ? 4'h0 : T4411;
  assign T4411 = T4413 ? T52 : T4412;
  assign T4412 = io_resetCounts ? 4'h0 : counts_727;
  assign T4413 = T10320 & T4414;
  assign T4414 = T76[10'h2d7:10'h2d7];
  assign T4415 = T68[1'h0:1'h0];
  assign T4416 = T68[1'h1:1'h1];
  assign T4417 = T68[2'h2:2'h2];
  assign T4418 = T4463 ? T4441 : T4419;
  assign T4419 = T4440 ? T4430 : T4420;
  assign T4420 = T4429 ? counts_729 : counts_728;
  assign T11073 = reset ? 4'h0 : T4421;
  assign T4421 = T4423 ? T52 : T4422;
  assign T4422 = io_resetCounts ? 4'h0 : counts_728;
  assign T4423 = T10320 & T4424;
  assign T4424 = T76[10'h2d8:10'h2d8];
  assign T11074 = reset ? 4'h0 : T4425;
  assign T4425 = T4427 ? T52 : T4426;
  assign T4426 = io_resetCounts ? 4'h0 : counts_729;
  assign T4427 = T10320 & T4428;
  assign T4428 = T76[10'h2d9:10'h2d9];
  assign T4429 = T68[1'h0:1'h0];
  assign T4430 = T4439 ? counts_731 : counts_730;
  assign T11075 = reset ? 4'h0 : T4431;
  assign T4431 = T4433 ? T52 : T4432;
  assign T4432 = io_resetCounts ? 4'h0 : counts_730;
  assign T4433 = T10320 & T4434;
  assign T4434 = T76[10'h2da:10'h2da];
  assign T11076 = reset ? 4'h0 : T4435;
  assign T4435 = T4437 ? T52 : T4436;
  assign T4436 = io_resetCounts ? 4'h0 : counts_731;
  assign T4437 = T10320 & T4438;
  assign T4438 = T76[10'h2db:10'h2db];
  assign T4439 = T68[1'h0:1'h0];
  assign T4440 = T68[1'h1:1'h1];
  assign T4441 = T4462 ? T4452 : T4442;
  assign T4442 = T4451 ? counts_733 : counts_732;
  assign T11077 = reset ? 4'h0 : T4443;
  assign T4443 = T4445 ? T52 : T4444;
  assign T4444 = io_resetCounts ? 4'h0 : counts_732;
  assign T4445 = T10320 & T4446;
  assign T4446 = T76[10'h2dc:10'h2dc];
  assign T11078 = reset ? 4'h0 : T4447;
  assign T4447 = T4449 ? T52 : T4448;
  assign T4448 = io_resetCounts ? 4'h0 : counts_733;
  assign T4449 = T10320 & T4450;
  assign T4450 = T76[10'h2dd:10'h2dd];
  assign T4451 = T68[1'h0:1'h0];
  assign T4452 = T4461 ? counts_735 : counts_734;
  assign T11079 = reset ? 4'h0 : T4453;
  assign T4453 = T4455 ? T52 : T4454;
  assign T4454 = io_resetCounts ? 4'h0 : counts_734;
  assign T4455 = T10320 & T4456;
  assign T4456 = T76[10'h2de:10'h2de];
  assign T11080 = reset ? 4'h0 : T4457;
  assign T4457 = T4459 ? T52 : T4458;
  assign T4458 = io_resetCounts ? 4'h0 : counts_735;
  assign T4459 = T10320 & T4460;
  assign T4460 = T76[10'h2df:10'h2df];
  assign T4461 = T68[1'h0:1'h0];
  assign T4462 = T68[1'h1:1'h1];
  assign T4463 = T68[2'h2:2'h2];
  assign T4464 = T68[2'h3:2'h3];
  assign T4465 = T68[3'h4:3'h4];
  assign T4466 = T4655 ? T4561 : T4467;
  assign T4467 = T4560 ? T4514 : T4468;
  assign T4468 = T4513 ? T4491 : T4469;
  assign T4469 = T4490 ? T4480 : T4470;
  assign T4470 = T4479 ? counts_737 : counts_736;
  assign T11081 = reset ? 4'h0 : T4471;
  assign T4471 = T4473 ? T52 : T4472;
  assign T4472 = io_resetCounts ? 4'h0 : counts_736;
  assign T4473 = T10320 & T4474;
  assign T4474 = T76[10'h2e0:10'h2e0];
  assign T11082 = reset ? 4'h0 : T4475;
  assign T4475 = T4477 ? T52 : T4476;
  assign T4476 = io_resetCounts ? 4'h0 : counts_737;
  assign T4477 = T10320 & T4478;
  assign T4478 = T76[10'h2e1:10'h2e1];
  assign T4479 = T68[1'h0:1'h0];
  assign T4480 = T4489 ? counts_739 : counts_738;
  assign T11083 = reset ? 4'h0 : T4481;
  assign T4481 = T4483 ? T52 : T4482;
  assign T4482 = io_resetCounts ? 4'h0 : counts_738;
  assign T4483 = T10320 & T4484;
  assign T4484 = T76[10'h2e2:10'h2e2];
  assign T11084 = reset ? 4'h0 : T4485;
  assign T4485 = T4487 ? T52 : T4486;
  assign T4486 = io_resetCounts ? 4'h0 : counts_739;
  assign T4487 = T10320 & T4488;
  assign T4488 = T76[10'h2e3:10'h2e3];
  assign T4489 = T68[1'h0:1'h0];
  assign T4490 = T68[1'h1:1'h1];
  assign T4491 = T4512 ? T4502 : T4492;
  assign T4492 = T4501 ? counts_741 : counts_740;
  assign T11085 = reset ? 4'h0 : T4493;
  assign T4493 = T4495 ? T52 : T4494;
  assign T4494 = io_resetCounts ? 4'h0 : counts_740;
  assign T4495 = T10320 & T4496;
  assign T4496 = T76[10'h2e4:10'h2e4];
  assign T11086 = reset ? 4'h0 : T4497;
  assign T4497 = T4499 ? T52 : T4498;
  assign T4498 = io_resetCounts ? 4'h0 : counts_741;
  assign T4499 = T10320 & T4500;
  assign T4500 = T76[10'h2e5:10'h2e5];
  assign T4501 = T68[1'h0:1'h0];
  assign T4502 = T4511 ? counts_743 : counts_742;
  assign T11087 = reset ? 4'h0 : T4503;
  assign T4503 = T4505 ? T52 : T4504;
  assign T4504 = io_resetCounts ? 4'h0 : counts_742;
  assign T4505 = T10320 & T4506;
  assign T4506 = T76[10'h2e6:10'h2e6];
  assign T11088 = reset ? 4'h0 : T4507;
  assign T4507 = T4509 ? T52 : T4508;
  assign T4508 = io_resetCounts ? 4'h0 : counts_743;
  assign T4509 = T10320 & T4510;
  assign T4510 = T76[10'h2e7:10'h2e7];
  assign T4511 = T68[1'h0:1'h0];
  assign T4512 = T68[1'h1:1'h1];
  assign T4513 = T68[2'h2:2'h2];
  assign T4514 = T4559 ? T4537 : T4515;
  assign T4515 = T4536 ? T4526 : T4516;
  assign T4516 = T4525 ? counts_745 : counts_744;
  assign T11089 = reset ? 4'h0 : T4517;
  assign T4517 = T4519 ? T52 : T4518;
  assign T4518 = io_resetCounts ? 4'h0 : counts_744;
  assign T4519 = T10320 & T4520;
  assign T4520 = T76[10'h2e8:10'h2e8];
  assign T11090 = reset ? 4'h0 : T4521;
  assign T4521 = T4523 ? T52 : T4522;
  assign T4522 = io_resetCounts ? 4'h0 : counts_745;
  assign T4523 = T10320 & T4524;
  assign T4524 = T76[10'h2e9:10'h2e9];
  assign T4525 = T68[1'h0:1'h0];
  assign T4526 = T4535 ? counts_747 : counts_746;
  assign T11091 = reset ? 4'h0 : T4527;
  assign T4527 = T4529 ? T52 : T4528;
  assign T4528 = io_resetCounts ? 4'h0 : counts_746;
  assign T4529 = T10320 & T4530;
  assign T4530 = T76[10'h2ea:10'h2ea];
  assign T11092 = reset ? 4'h0 : T4531;
  assign T4531 = T4533 ? T52 : T4532;
  assign T4532 = io_resetCounts ? 4'h0 : counts_747;
  assign T4533 = T10320 & T4534;
  assign T4534 = T76[10'h2eb:10'h2eb];
  assign T4535 = T68[1'h0:1'h0];
  assign T4536 = T68[1'h1:1'h1];
  assign T4537 = T4558 ? T4548 : T4538;
  assign T4538 = T4547 ? counts_749 : counts_748;
  assign T11093 = reset ? 4'h0 : T4539;
  assign T4539 = T4541 ? T52 : T4540;
  assign T4540 = io_resetCounts ? 4'h0 : counts_748;
  assign T4541 = T10320 & T4542;
  assign T4542 = T76[10'h2ec:10'h2ec];
  assign T11094 = reset ? 4'h0 : T4543;
  assign T4543 = T4545 ? T52 : T4544;
  assign T4544 = io_resetCounts ? 4'h0 : counts_749;
  assign T4545 = T10320 & T4546;
  assign T4546 = T76[10'h2ed:10'h2ed];
  assign T4547 = T68[1'h0:1'h0];
  assign T4548 = T4557 ? counts_751 : counts_750;
  assign T11095 = reset ? 4'h0 : T4549;
  assign T4549 = T4551 ? T52 : T4550;
  assign T4550 = io_resetCounts ? 4'h0 : counts_750;
  assign T4551 = T10320 & T4552;
  assign T4552 = T76[10'h2ee:10'h2ee];
  assign T11096 = reset ? 4'h0 : T4553;
  assign T4553 = T4555 ? T52 : T4554;
  assign T4554 = io_resetCounts ? 4'h0 : counts_751;
  assign T4555 = T10320 & T4556;
  assign T4556 = T76[10'h2ef:10'h2ef];
  assign T4557 = T68[1'h0:1'h0];
  assign T4558 = T68[1'h1:1'h1];
  assign T4559 = T68[2'h2:2'h2];
  assign T4560 = T68[2'h3:2'h3];
  assign T4561 = T4654 ? T4608 : T4562;
  assign T4562 = T4607 ? T4585 : T4563;
  assign T4563 = T4584 ? T4574 : T4564;
  assign T4564 = T4573 ? counts_753 : counts_752;
  assign T11097 = reset ? 4'h0 : T4565;
  assign T4565 = T4567 ? T52 : T4566;
  assign T4566 = io_resetCounts ? 4'h0 : counts_752;
  assign T4567 = T10320 & T4568;
  assign T4568 = T76[10'h2f0:10'h2f0];
  assign T11098 = reset ? 4'h0 : T4569;
  assign T4569 = T4571 ? T52 : T4570;
  assign T4570 = io_resetCounts ? 4'h0 : counts_753;
  assign T4571 = T10320 & T4572;
  assign T4572 = T76[10'h2f1:10'h2f1];
  assign T4573 = T68[1'h0:1'h0];
  assign T4574 = T4583 ? counts_755 : counts_754;
  assign T11099 = reset ? 4'h0 : T4575;
  assign T4575 = T4577 ? T52 : T4576;
  assign T4576 = io_resetCounts ? 4'h0 : counts_754;
  assign T4577 = T10320 & T4578;
  assign T4578 = T76[10'h2f2:10'h2f2];
  assign T11100 = reset ? 4'h0 : T4579;
  assign T4579 = T4581 ? T52 : T4580;
  assign T4580 = io_resetCounts ? 4'h0 : counts_755;
  assign T4581 = T10320 & T4582;
  assign T4582 = T76[10'h2f3:10'h2f3];
  assign T4583 = T68[1'h0:1'h0];
  assign T4584 = T68[1'h1:1'h1];
  assign T4585 = T4606 ? T4596 : T4586;
  assign T4586 = T4595 ? counts_757 : counts_756;
  assign T11101 = reset ? 4'h0 : T4587;
  assign T4587 = T4589 ? T52 : T4588;
  assign T4588 = io_resetCounts ? 4'h0 : counts_756;
  assign T4589 = T10320 & T4590;
  assign T4590 = T76[10'h2f4:10'h2f4];
  assign T11102 = reset ? 4'h0 : T4591;
  assign T4591 = T4593 ? T52 : T4592;
  assign T4592 = io_resetCounts ? 4'h0 : counts_757;
  assign T4593 = T10320 & T4594;
  assign T4594 = T76[10'h2f5:10'h2f5];
  assign T4595 = T68[1'h0:1'h0];
  assign T4596 = T4605 ? counts_759 : counts_758;
  assign T11103 = reset ? 4'h0 : T4597;
  assign T4597 = T4599 ? T52 : T4598;
  assign T4598 = io_resetCounts ? 4'h0 : counts_758;
  assign T4599 = T10320 & T4600;
  assign T4600 = T76[10'h2f6:10'h2f6];
  assign T11104 = reset ? 4'h0 : T4601;
  assign T4601 = T4603 ? T52 : T4602;
  assign T4602 = io_resetCounts ? 4'h0 : counts_759;
  assign T4603 = T10320 & T4604;
  assign T4604 = T76[10'h2f7:10'h2f7];
  assign T4605 = T68[1'h0:1'h0];
  assign T4606 = T68[1'h1:1'h1];
  assign T4607 = T68[2'h2:2'h2];
  assign T4608 = T4653 ? T4631 : T4609;
  assign T4609 = T4630 ? T4620 : T4610;
  assign T4610 = T4619 ? counts_761 : counts_760;
  assign T11105 = reset ? 4'h0 : T4611;
  assign T4611 = T4613 ? T52 : T4612;
  assign T4612 = io_resetCounts ? 4'h0 : counts_760;
  assign T4613 = T10320 & T4614;
  assign T4614 = T76[10'h2f8:10'h2f8];
  assign T11106 = reset ? 4'h0 : T4615;
  assign T4615 = T4617 ? T52 : T4616;
  assign T4616 = io_resetCounts ? 4'h0 : counts_761;
  assign T4617 = T10320 & T4618;
  assign T4618 = T76[10'h2f9:10'h2f9];
  assign T4619 = T68[1'h0:1'h0];
  assign T4620 = T4629 ? counts_763 : counts_762;
  assign T11107 = reset ? 4'h0 : T4621;
  assign T4621 = T4623 ? T52 : T4622;
  assign T4622 = io_resetCounts ? 4'h0 : counts_762;
  assign T4623 = T10320 & T4624;
  assign T4624 = T76[10'h2fa:10'h2fa];
  assign T11108 = reset ? 4'h0 : T4625;
  assign T4625 = T4627 ? T52 : T4626;
  assign T4626 = io_resetCounts ? 4'h0 : counts_763;
  assign T4627 = T10320 & T4628;
  assign T4628 = T76[10'h2fb:10'h2fb];
  assign T4629 = T68[1'h0:1'h0];
  assign T4630 = T68[1'h1:1'h1];
  assign T4631 = T4652 ? T4642 : T4632;
  assign T4632 = T4641 ? counts_765 : counts_764;
  assign T11109 = reset ? 4'h0 : T4633;
  assign T4633 = T4635 ? T52 : T4634;
  assign T4634 = io_resetCounts ? 4'h0 : counts_764;
  assign T4635 = T10320 & T4636;
  assign T4636 = T76[10'h2fc:10'h2fc];
  assign T11110 = reset ? 4'h0 : T4637;
  assign T4637 = T4639 ? T52 : T4638;
  assign T4638 = io_resetCounts ? 4'h0 : counts_765;
  assign T4639 = T10320 & T4640;
  assign T4640 = T76[10'h2fd:10'h2fd];
  assign T4641 = T68[1'h0:1'h0];
  assign T4642 = T4651 ? counts_767 : counts_766;
  assign T11111 = reset ? 4'h0 : T4643;
  assign T4643 = T4645 ? T52 : T4644;
  assign T4644 = io_resetCounts ? 4'h0 : counts_766;
  assign T4645 = T10320 & T4646;
  assign T4646 = T76[10'h2fe:10'h2fe];
  assign T11112 = reset ? 4'h0 : T4647;
  assign T4647 = T4649 ? T52 : T4648;
  assign T4648 = io_resetCounts ? 4'h0 : counts_767;
  assign T4649 = T10320 & T4650;
  assign T4650 = T76[10'h2ff:10'h2ff];
  assign T4651 = T68[1'h0:1'h0];
  assign T4652 = T68[1'h1:1'h1];
  assign T4653 = T68[2'h2:2'h2];
  assign T4654 = T68[2'h3:2'h3];
  assign T4655 = T68[3'h4:3'h4];
  assign T4656 = T68[3'h5:3'h5];
  assign T4657 = T68[3'h6:3'h6];
  assign T4658 = T68[3'h7:3'h7];
  assign T4659 = T6192 ? T5426 : T4660;
  assign T4660 = T5425 ? T5043 : T4661;
  assign T4661 = T5042 ? T4852 : T4662;
  assign T4662 = T4851 ? T4757 : T4663;
  assign T4663 = T4756 ? T4710 : T4664;
  assign T4664 = T4709 ? T4687 : T4665;
  assign T4665 = T4686 ? T4676 : T4666;
  assign T4666 = T4675 ? counts_769 : counts_768;
  assign T11113 = reset ? 4'h0 : T4667;
  assign T4667 = T4669 ? T52 : T4668;
  assign T4668 = io_resetCounts ? 4'h0 : counts_768;
  assign T4669 = T10320 & T4670;
  assign T4670 = T76[10'h300:10'h300];
  assign T11114 = reset ? 4'h0 : T4671;
  assign T4671 = T4673 ? T52 : T4672;
  assign T4672 = io_resetCounts ? 4'h0 : counts_769;
  assign T4673 = T10320 & T4674;
  assign T4674 = T76[10'h301:10'h301];
  assign T4675 = T68[1'h0:1'h0];
  assign T4676 = T4685 ? counts_771 : counts_770;
  assign T11115 = reset ? 4'h0 : T4677;
  assign T4677 = T4679 ? T52 : T4678;
  assign T4678 = io_resetCounts ? 4'h0 : counts_770;
  assign T4679 = T10320 & T4680;
  assign T4680 = T76[10'h302:10'h302];
  assign T11116 = reset ? 4'h0 : T4681;
  assign T4681 = T4683 ? T52 : T4682;
  assign T4682 = io_resetCounts ? 4'h0 : counts_771;
  assign T4683 = T10320 & T4684;
  assign T4684 = T76[10'h303:10'h303];
  assign T4685 = T68[1'h0:1'h0];
  assign T4686 = T68[1'h1:1'h1];
  assign T4687 = T4708 ? T4698 : T4688;
  assign T4688 = T4697 ? counts_773 : counts_772;
  assign T11117 = reset ? 4'h0 : T4689;
  assign T4689 = T4691 ? T52 : T4690;
  assign T4690 = io_resetCounts ? 4'h0 : counts_772;
  assign T4691 = T10320 & T4692;
  assign T4692 = T76[10'h304:10'h304];
  assign T11118 = reset ? 4'h0 : T4693;
  assign T4693 = T4695 ? T52 : T4694;
  assign T4694 = io_resetCounts ? 4'h0 : counts_773;
  assign T4695 = T10320 & T4696;
  assign T4696 = T76[10'h305:10'h305];
  assign T4697 = T68[1'h0:1'h0];
  assign T4698 = T4707 ? counts_775 : counts_774;
  assign T11119 = reset ? 4'h0 : T4699;
  assign T4699 = T4701 ? T52 : T4700;
  assign T4700 = io_resetCounts ? 4'h0 : counts_774;
  assign T4701 = T10320 & T4702;
  assign T4702 = T76[10'h306:10'h306];
  assign T11120 = reset ? 4'h0 : T4703;
  assign T4703 = T4705 ? T52 : T4704;
  assign T4704 = io_resetCounts ? 4'h0 : counts_775;
  assign T4705 = T10320 & T4706;
  assign T4706 = T76[10'h307:10'h307];
  assign T4707 = T68[1'h0:1'h0];
  assign T4708 = T68[1'h1:1'h1];
  assign T4709 = T68[2'h2:2'h2];
  assign T4710 = T4755 ? T4733 : T4711;
  assign T4711 = T4732 ? T4722 : T4712;
  assign T4712 = T4721 ? counts_777 : counts_776;
  assign T11121 = reset ? 4'h0 : T4713;
  assign T4713 = T4715 ? T52 : T4714;
  assign T4714 = io_resetCounts ? 4'h0 : counts_776;
  assign T4715 = T10320 & T4716;
  assign T4716 = T76[10'h308:10'h308];
  assign T11122 = reset ? 4'h0 : T4717;
  assign T4717 = T4719 ? T52 : T4718;
  assign T4718 = io_resetCounts ? 4'h0 : counts_777;
  assign T4719 = T10320 & T4720;
  assign T4720 = T76[10'h309:10'h309];
  assign T4721 = T68[1'h0:1'h0];
  assign T4722 = T4731 ? counts_779 : counts_778;
  assign T11123 = reset ? 4'h0 : T4723;
  assign T4723 = T4725 ? T52 : T4724;
  assign T4724 = io_resetCounts ? 4'h0 : counts_778;
  assign T4725 = T10320 & T4726;
  assign T4726 = T76[10'h30a:10'h30a];
  assign T11124 = reset ? 4'h0 : T4727;
  assign T4727 = T4729 ? T52 : T4728;
  assign T4728 = io_resetCounts ? 4'h0 : counts_779;
  assign T4729 = T10320 & T4730;
  assign T4730 = T76[10'h30b:10'h30b];
  assign T4731 = T68[1'h0:1'h0];
  assign T4732 = T68[1'h1:1'h1];
  assign T4733 = T4754 ? T4744 : T4734;
  assign T4734 = T4743 ? counts_781 : counts_780;
  assign T11125 = reset ? 4'h0 : T4735;
  assign T4735 = T4737 ? T52 : T4736;
  assign T4736 = io_resetCounts ? 4'h0 : counts_780;
  assign T4737 = T10320 & T4738;
  assign T4738 = T76[10'h30c:10'h30c];
  assign T11126 = reset ? 4'h0 : T4739;
  assign T4739 = T4741 ? T52 : T4740;
  assign T4740 = io_resetCounts ? 4'h0 : counts_781;
  assign T4741 = T10320 & T4742;
  assign T4742 = T76[10'h30d:10'h30d];
  assign T4743 = T68[1'h0:1'h0];
  assign T4744 = T4753 ? counts_783 : counts_782;
  assign T11127 = reset ? 4'h0 : T4745;
  assign T4745 = T4747 ? T52 : T4746;
  assign T4746 = io_resetCounts ? 4'h0 : counts_782;
  assign T4747 = T10320 & T4748;
  assign T4748 = T76[10'h30e:10'h30e];
  assign T11128 = reset ? 4'h0 : T4749;
  assign T4749 = T4751 ? T52 : T4750;
  assign T4750 = io_resetCounts ? 4'h0 : counts_783;
  assign T4751 = T10320 & T4752;
  assign T4752 = T76[10'h30f:10'h30f];
  assign T4753 = T68[1'h0:1'h0];
  assign T4754 = T68[1'h1:1'h1];
  assign T4755 = T68[2'h2:2'h2];
  assign T4756 = T68[2'h3:2'h3];
  assign T4757 = T4850 ? T4804 : T4758;
  assign T4758 = T4803 ? T4781 : T4759;
  assign T4759 = T4780 ? T4770 : T4760;
  assign T4760 = T4769 ? counts_785 : counts_784;
  assign T11129 = reset ? 4'h0 : T4761;
  assign T4761 = T4763 ? T52 : T4762;
  assign T4762 = io_resetCounts ? 4'h0 : counts_784;
  assign T4763 = T10320 & T4764;
  assign T4764 = T76[10'h310:10'h310];
  assign T11130 = reset ? 4'h0 : T4765;
  assign T4765 = T4767 ? T52 : T4766;
  assign T4766 = io_resetCounts ? 4'h0 : counts_785;
  assign T4767 = T10320 & T4768;
  assign T4768 = T76[10'h311:10'h311];
  assign T4769 = T68[1'h0:1'h0];
  assign T4770 = T4779 ? counts_787 : counts_786;
  assign T11131 = reset ? 4'h0 : T4771;
  assign T4771 = T4773 ? T52 : T4772;
  assign T4772 = io_resetCounts ? 4'h0 : counts_786;
  assign T4773 = T10320 & T4774;
  assign T4774 = T76[10'h312:10'h312];
  assign T11132 = reset ? 4'h0 : T4775;
  assign T4775 = T4777 ? T52 : T4776;
  assign T4776 = io_resetCounts ? 4'h0 : counts_787;
  assign T4777 = T10320 & T4778;
  assign T4778 = T76[10'h313:10'h313];
  assign T4779 = T68[1'h0:1'h0];
  assign T4780 = T68[1'h1:1'h1];
  assign T4781 = T4802 ? T4792 : T4782;
  assign T4782 = T4791 ? counts_789 : counts_788;
  assign T11133 = reset ? 4'h0 : T4783;
  assign T4783 = T4785 ? T52 : T4784;
  assign T4784 = io_resetCounts ? 4'h0 : counts_788;
  assign T4785 = T10320 & T4786;
  assign T4786 = T76[10'h314:10'h314];
  assign T11134 = reset ? 4'h0 : T4787;
  assign T4787 = T4789 ? T52 : T4788;
  assign T4788 = io_resetCounts ? 4'h0 : counts_789;
  assign T4789 = T10320 & T4790;
  assign T4790 = T76[10'h315:10'h315];
  assign T4791 = T68[1'h0:1'h0];
  assign T4792 = T4801 ? counts_791 : counts_790;
  assign T11135 = reset ? 4'h0 : T4793;
  assign T4793 = T4795 ? T52 : T4794;
  assign T4794 = io_resetCounts ? 4'h0 : counts_790;
  assign T4795 = T10320 & T4796;
  assign T4796 = T76[10'h316:10'h316];
  assign T11136 = reset ? 4'h0 : T4797;
  assign T4797 = T4799 ? T52 : T4798;
  assign T4798 = io_resetCounts ? 4'h0 : counts_791;
  assign T4799 = T10320 & T4800;
  assign T4800 = T76[10'h317:10'h317];
  assign T4801 = T68[1'h0:1'h0];
  assign T4802 = T68[1'h1:1'h1];
  assign T4803 = T68[2'h2:2'h2];
  assign T4804 = T4849 ? T4827 : T4805;
  assign T4805 = T4826 ? T4816 : T4806;
  assign T4806 = T4815 ? counts_793 : counts_792;
  assign T11137 = reset ? 4'h0 : T4807;
  assign T4807 = T4809 ? T52 : T4808;
  assign T4808 = io_resetCounts ? 4'h0 : counts_792;
  assign T4809 = T10320 & T4810;
  assign T4810 = T76[10'h318:10'h318];
  assign T11138 = reset ? 4'h0 : T4811;
  assign T4811 = T4813 ? T52 : T4812;
  assign T4812 = io_resetCounts ? 4'h0 : counts_793;
  assign T4813 = T10320 & T4814;
  assign T4814 = T76[10'h319:10'h319];
  assign T4815 = T68[1'h0:1'h0];
  assign T4816 = T4825 ? counts_795 : counts_794;
  assign T11139 = reset ? 4'h0 : T4817;
  assign T4817 = T4819 ? T52 : T4818;
  assign T4818 = io_resetCounts ? 4'h0 : counts_794;
  assign T4819 = T10320 & T4820;
  assign T4820 = T76[10'h31a:10'h31a];
  assign T11140 = reset ? 4'h0 : T4821;
  assign T4821 = T4823 ? T52 : T4822;
  assign T4822 = io_resetCounts ? 4'h0 : counts_795;
  assign T4823 = T10320 & T4824;
  assign T4824 = T76[10'h31b:10'h31b];
  assign T4825 = T68[1'h0:1'h0];
  assign T4826 = T68[1'h1:1'h1];
  assign T4827 = T4848 ? T4838 : T4828;
  assign T4828 = T4837 ? counts_797 : counts_796;
  assign T11141 = reset ? 4'h0 : T4829;
  assign T4829 = T4831 ? T52 : T4830;
  assign T4830 = io_resetCounts ? 4'h0 : counts_796;
  assign T4831 = T10320 & T4832;
  assign T4832 = T76[10'h31c:10'h31c];
  assign T11142 = reset ? 4'h0 : T4833;
  assign T4833 = T4835 ? T52 : T4834;
  assign T4834 = io_resetCounts ? 4'h0 : counts_797;
  assign T4835 = T10320 & T4836;
  assign T4836 = T76[10'h31d:10'h31d];
  assign T4837 = T68[1'h0:1'h0];
  assign T4838 = T4847 ? counts_799 : counts_798;
  assign T11143 = reset ? 4'h0 : T4839;
  assign T4839 = T4841 ? T52 : T4840;
  assign T4840 = io_resetCounts ? 4'h0 : counts_798;
  assign T4841 = T10320 & T4842;
  assign T4842 = T76[10'h31e:10'h31e];
  assign T11144 = reset ? 4'h0 : T4843;
  assign T4843 = T4845 ? T52 : T4844;
  assign T4844 = io_resetCounts ? 4'h0 : counts_799;
  assign T4845 = T10320 & T4846;
  assign T4846 = T76[10'h31f:10'h31f];
  assign T4847 = T68[1'h0:1'h0];
  assign T4848 = T68[1'h1:1'h1];
  assign T4849 = T68[2'h2:2'h2];
  assign T4850 = T68[2'h3:2'h3];
  assign T4851 = T68[3'h4:3'h4];
  assign T4852 = T5041 ? T4947 : T4853;
  assign T4853 = T4946 ? T4900 : T4854;
  assign T4854 = T4899 ? T4877 : T4855;
  assign T4855 = T4876 ? T4866 : T4856;
  assign T4856 = T4865 ? counts_801 : counts_800;
  assign T11145 = reset ? 4'h0 : T4857;
  assign T4857 = T4859 ? T52 : T4858;
  assign T4858 = io_resetCounts ? 4'h0 : counts_800;
  assign T4859 = T10320 & T4860;
  assign T4860 = T76[10'h320:10'h320];
  assign T11146 = reset ? 4'h0 : T4861;
  assign T4861 = T4863 ? T52 : T4862;
  assign T4862 = io_resetCounts ? 4'h0 : counts_801;
  assign T4863 = T10320 & T4864;
  assign T4864 = T76[10'h321:10'h321];
  assign T4865 = T68[1'h0:1'h0];
  assign T4866 = T4875 ? counts_803 : counts_802;
  assign T11147 = reset ? 4'h0 : T4867;
  assign T4867 = T4869 ? T52 : T4868;
  assign T4868 = io_resetCounts ? 4'h0 : counts_802;
  assign T4869 = T10320 & T4870;
  assign T4870 = T76[10'h322:10'h322];
  assign T11148 = reset ? 4'h0 : T4871;
  assign T4871 = T4873 ? T52 : T4872;
  assign T4872 = io_resetCounts ? 4'h0 : counts_803;
  assign T4873 = T10320 & T4874;
  assign T4874 = T76[10'h323:10'h323];
  assign T4875 = T68[1'h0:1'h0];
  assign T4876 = T68[1'h1:1'h1];
  assign T4877 = T4898 ? T4888 : T4878;
  assign T4878 = T4887 ? counts_805 : counts_804;
  assign T11149 = reset ? 4'h0 : T4879;
  assign T4879 = T4881 ? T52 : T4880;
  assign T4880 = io_resetCounts ? 4'h0 : counts_804;
  assign T4881 = T10320 & T4882;
  assign T4882 = T76[10'h324:10'h324];
  assign T11150 = reset ? 4'h0 : T4883;
  assign T4883 = T4885 ? T52 : T4884;
  assign T4884 = io_resetCounts ? 4'h0 : counts_805;
  assign T4885 = T10320 & T4886;
  assign T4886 = T76[10'h325:10'h325];
  assign T4887 = T68[1'h0:1'h0];
  assign T4888 = T4897 ? counts_807 : counts_806;
  assign T11151 = reset ? 4'h0 : T4889;
  assign T4889 = T4891 ? T52 : T4890;
  assign T4890 = io_resetCounts ? 4'h0 : counts_806;
  assign T4891 = T10320 & T4892;
  assign T4892 = T76[10'h326:10'h326];
  assign T11152 = reset ? 4'h0 : T4893;
  assign T4893 = T4895 ? T52 : T4894;
  assign T4894 = io_resetCounts ? 4'h0 : counts_807;
  assign T4895 = T10320 & T4896;
  assign T4896 = T76[10'h327:10'h327];
  assign T4897 = T68[1'h0:1'h0];
  assign T4898 = T68[1'h1:1'h1];
  assign T4899 = T68[2'h2:2'h2];
  assign T4900 = T4945 ? T4923 : T4901;
  assign T4901 = T4922 ? T4912 : T4902;
  assign T4902 = T4911 ? counts_809 : counts_808;
  assign T11153 = reset ? 4'h0 : T4903;
  assign T4903 = T4905 ? T52 : T4904;
  assign T4904 = io_resetCounts ? 4'h0 : counts_808;
  assign T4905 = T10320 & T4906;
  assign T4906 = T76[10'h328:10'h328];
  assign T11154 = reset ? 4'h0 : T4907;
  assign T4907 = T4909 ? T52 : T4908;
  assign T4908 = io_resetCounts ? 4'h0 : counts_809;
  assign T4909 = T10320 & T4910;
  assign T4910 = T76[10'h329:10'h329];
  assign T4911 = T68[1'h0:1'h0];
  assign T4912 = T4921 ? counts_811 : counts_810;
  assign T11155 = reset ? 4'h0 : T4913;
  assign T4913 = T4915 ? T52 : T4914;
  assign T4914 = io_resetCounts ? 4'h0 : counts_810;
  assign T4915 = T10320 & T4916;
  assign T4916 = T76[10'h32a:10'h32a];
  assign T11156 = reset ? 4'h0 : T4917;
  assign T4917 = T4919 ? T52 : T4918;
  assign T4918 = io_resetCounts ? 4'h0 : counts_811;
  assign T4919 = T10320 & T4920;
  assign T4920 = T76[10'h32b:10'h32b];
  assign T4921 = T68[1'h0:1'h0];
  assign T4922 = T68[1'h1:1'h1];
  assign T4923 = T4944 ? T4934 : T4924;
  assign T4924 = T4933 ? counts_813 : counts_812;
  assign T11157 = reset ? 4'h0 : T4925;
  assign T4925 = T4927 ? T52 : T4926;
  assign T4926 = io_resetCounts ? 4'h0 : counts_812;
  assign T4927 = T10320 & T4928;
  assign T4928 = T76[10'h32c:10'h32c];
  assign T11158 = reset ? 4'h0 : T4929;
  assign T4929 = T4931 ? T52 : T4930;
  assign T4930 = io_resetCounts ? 4'h0 : counts_813;
  assign T4931 = T10320 & T4932;
  assign T4932 = T76[10'h32d:10'h32d];
  assign T4933 = T68[1'h0:1'h0];
  assign T4934 = T4943 ? counts_815 : counts_814;
  assign T11159 = reset ? 4'h0 : T4935;
  assign T4935 = T4937 ? T52 : T4936;
  assign T4936 = io_resetCounts ? 4'h0 : counts_814;
  assign T4937 = T10320 & T4938;
  assign T4938 = T76[10'h32e:10'h32e];
  assign T11160 = reset ? 4'h0 : T4939;
  assign T4939 = T4941 ? T52 : T4940;
  assign T4940 = io_resetCounts ? 4'h0 : counts_815;
  assign T4941 = T10320 & T4942;
  assign T4942 = T76[10'h32f:10'h32f];
  assign T4943 = T68[1'h0:1'h0];
  assign T4944 = T68[1'h1:1'h1];
  assign T4945 = T68[2'h2:2'h2];
  assign T4946 = T68[2'h3:2'h3];
  assign T4947 = T5040 ? T4994 : T4948;
  assign T4948 = T4993 ? T4971 : T4949;
  assign T4949 = T4970 ? T4960 : T4950;
  assign T4950 = T4959 ? counts_817 : counts_816;
  assign T11161 = reset ? 4'h0 : T4951;
  assign T4951 = T4953 ? T52 : T4952;
  assign T4952 = io_resetCounts ? 4'h0 : counts_816;
  assign T4953 = T10320 & T4954;
  assign T4954 = T76[10'h330:10'h330];
  assign T11162 = reset ? 4'h0 : T4955;
  assign T4955 = T4957 ? T52 : T4956;
  assign T4956 = io_resetCounts ? 4'h0 : counts_817;
  assign T4957 = T10320 & T4958;
  assign T4958 = T76[10'h331:10'h331];
  assign T4959 = T68[1'h0:1'h0];
  assign T4960 = T4969 ? counts_819 : counts_818;
  assign T11163 = reset ? 4'h0 : T4961;
  assign T4961 = T4963 ? T52 : T4962;
  assign T4962 = io_resetCounts ? 4'h0 : counts_818;
  assign T4963 = T10320 & T4964;
  assign T4964 = T76[10'h332:10'h332];
  assign T11164 = reset ? 4'h0 : T4965;
  assign T4965 = T4967 ? T52 : T4966;
  assign T4966 = io_resetCounts ? 4'h0 : counts_819;
  assign T4967 = T10320 & T4968;
  assign T4968 = T76[10'h333:10'h333];
  assign T4969 = T68[1'h0:1'h0];
  assign T4970 = T68[1'h1:1'h1];
  assign T4971 = T4992 ? T4982 : T4972;
  assign T4972 = T4981 ? counts_821 : counts_820;
  assign T11165 = reset ? 4'h0 : T4973;
  assign T4973 = T4975 ? T52 : T4974;
  assign T4974 = io_resetCounts ? 4'h0 : counts_820;
  assign T4975 = T10320 & T4976;
  assign T4976 = T76[10'h334:10'h334];
  assign T11166 = reset ? 4'h0 : T4977;
  assign T4977 = T4979 ? T52 : T4978;
  assign T4978 = io_resetCounts ? 4'h0 : counts_821;
  assign T4979 = T10320 & T4980;
  assign T4980 = T76[10'h335:10'h335];
  assign T4981 = T68[1'h0:1'h0];
  assign T4982 = T4991 ? counts_823 : counts_822;
  assign T11167 = reset ? 4'h0 : T4983;
  assign T4983 = T4985 ? T52 : T4984;
  assign T4984 = io_resetCounts ? 4'h0 : counts_822;
  assign T4985 = T10320 & T4986;
  assign T4986 = T76[10'h336:10'h336];
  assign T11168 = reset ? 4'h0 : T4987;
  assign T4987 = T4989 ? T52 : T4988;
  assign T4988 = io_resetCounts ? 4'h0 : counts_823;
  assign T4989 = T10320 & T4990;
  assign T4990 = T76[10'h337:10'h337];
  assign T4991 = T68[1'h0:1'h0];
  assign T4992 = T68[1'h1:1'h1];
  assign T4993 = T68[2'h2:2'h2];
  assign T4994 = T5039 ? T5017 : T4995;
  assign T4995 = T5016 ? T5006 : T4996;
  assign T4996 = T5005 ? counts_825 : counts_824;
  assign T11169 = reset ? 4'h0 : T4997;
  assign T4997 = T4999 ? T52 : T4998;
  assign T4998 = io_resetCounts ? 4'h0 : counts_824;
  assign T4999 = T10320 & T5000;
  assign T5000 = T76[10'h338:10'h338];
  assign T11170 = reset ? 4'h0 : T5001;
  assign T5001 = T5003 ? T52 : T5002;
  assign T5002 = io_resetCounts ? 4'h0 : counts_825;
  assign T5003 = T10320 & T5004;
  assign T5004 = T76[10'h339:10'h339];
  assign T5005 = T68[1'h0:1'h0];
  assign T5006 = T5015 ? counts_827 : counts_826;
  assign T11171 = reset ? 4'h0 : T5007;
  assign T5007 = T5009 ? T52 : T5008;
  assign T5008 = io_resetCounts ? 4'h0 : counts_826;
  assign T5009 = T10320 & T5010;
  assign T5010 = T76[10'h33a:10'h33a];
  assign T11172 = reset ? 4'h0 : T5011;
  assign T5011 = T5013 ? T52 : T5012;
  assign T5012 = io_resetCounts ? 4'h0 : counts_827;
  assign T5013 = T10320 & T5014;
  assign T5014 = T76[10'h33b:10'h33b];
  assign T5015 = T68[1'h0:1'h0];
  assign T5016 = T68[1'h1:1'h1];
  assign T5017 = T5038 ? T5028 : T5018;
  assign T5018 = T5027 ? counts_829 : counts_828;
  assign T11173 = reset ? 4'h0 : T5019;
  assign T5019 = T5021 ? T52 : T5020;
  assign T5020 = io_resetCounts ? 4'h0 : counts_828;
  assign T5021 = T10320 & T5022;
  assign T5022 = T76[10'h33c:10'h33c];
  assign T11174 = reset ? 4'h0 : T5023;
  assign T5023 = T5025 ? T52 : T5024;
  assign T5024 = io_resetCounts ? 4'h0 : counts_829;
  assign T5025 = T10320 & T5026;
  assign T5026 = T76[10'h33d:10'h33d];
  assign T5027 = T68[1'h0:1'h0];
  assign T5028 = T5037 ? counts_831 : counts_830;
  assign T11175 = reset ? 4'h0 : T5029;
  assign T5029 = T5031 ? T52 : T5030;
  assign T5030 = io_resetCounts ? 4'h0 : counts_830;
  assign T5031 = T10320 & T5032;
  assign T5032 = T76[10'h33e:10'h33e];
  assign T11176 = reset ? 4'h0 : T5033;
  assign T5033 = T5035 ? T52 : T5034;
  assign T5034 = io_resetCounts ? 4'h0 : counts_831;
  assign T5035 = T10320 & T5036;
  assign T5036 = T76[10'h33f:10'h33f];
  assign T5037 = T68[1'h0:1'h0];
  assign T5038 = T68[1'h1:1'h1];
  assign T5039 = T68[2'h2:2'h2];
  assign T5040 = T68[2'h3:2'h3];
  assign T5041 = T68[3'h4:3'h4];
  assign T5042 = T68[3'h5:3'h5];
  assign T5043 = T5424 ? T5234 : T5044;
  assign T5044 = T5233 ? T5139 : T5045;
  assign T5045 = T5138 ? T5092 : T5046;
  assign T5046 = T5091 ? T5069 : T5047;
  assign T5047 = T5068 ? T5058 : T5048;
  assign T5048 = T5057 ? counts_833 : counts_832;
  assign T11177 = reset ? 4'h0 : T5049;
  assign T5049 = T5051 ? T52 : T5050;
  assign T5050 = io_resetCounts ? 4'h0 : counts_832;
  assign T5051 = T10320 & T5052;
  assign T5052 = T76[10'h340:10'h340];
  assign T11178 = reset ? 4'h0 : T5053;
  assign T5053 = T5055 ? T52 : T5054;
  assign T5054 = io_resetCounts ? 4'h0 : counts_833;
  assign T5055 = T10320 & T5056;
  assign T5056 = T76[10'h341:10'h341];
  assign T5057 = T68[1'h0:1'h0];
  assign T5058 = T5067 ? counts_835 : counts_834;
  assign T11179 = reset ? 4'h0 : T5059;
  assign T5059 = T5061 ? T52 : T5060;
  assign T5060 = io_resetCounts ? 4'h0 : counts_834;
  assign T5061 = T10320 & T5062;
  assign T5062 = T76[10'h342:10'h342];
  assign T11180 = reset ? 4'h0 : T5063;
  assign T5063 = T5065 ? T52 : T5064;
  assign T5064 = io_resetCounts ? 4'h0 : counts_835;
  assign T5065 = T10320 & T5066;
  assign T5066 = T76[10'h343:10'h343];
  assign T5067 = T68[1'h0:1'h0];
  assign T5068 = T68[1'h1:1'h1];
  assign T5069 = T5090 ? T5080 : T5070;
  assign T5070 = T5079 ? counts_837 : counts_836;
  assign T11181 = reset ? 4'h0 : T5071;
  assign T5071 = T5073 ? T52 : T5072;
  assign T5072 = io_resetCounts ? 4'h0 : counts_836;
  assign T5073 = T10320 & T5074;
  assign T5074 = T76[10'h344:10'h344];
  assign T11182 = reset ? 4'h0 : T5075;
  assign T5075 = T5077 ? T52 : T5076;
  assign T5076 = io_resetCounts ? 4'h0 : counts_837;
  assign T5077 = T10320 & T5078;
  assign T5078 = T76[10'h345:10'h345];
  assign T5079 = T68[1'h0:1'h0];
  assign T5080 = T5089 ? counts_839 : counts_838;
  assign T11183 = reset ? 4'h0 : T5081;
  assign T5081 = T5083 ? T52 : T5082;
  assign T5082 = io_resetCounts ? 4'h0 : counts_838;
  assign T5083 = T10320 & T5084;
  assign T5084 = T76[10'h346:10'h346];
  assign T11184 = reset ? 4'h0 : T5085;
  assign T5085 = T5087 ? T52 : T5086;
  assign T5086 = io_resetCounts ? 4'h0 : counts_839;
  assign T5087 = T10320 & T5088;
  assign T5088 = T76[10'h347:10'h347];
  assign T5089 = T68[1'h0:1'h0];
  assign T5090 = T68[1'h1:1'h1];
  assign T5091 = T68[2'h2:2'h2];
  assign T5092 = T5137 ? T5115 : T5093;
  assign T5093 = T5114 ? T5104 : T5094;
  assign T5094 = T5103 ? counts_841 : counts_840;
  assign T11185 = reset ? 4'h0 : T5095;
  assign T5095 = T5097 ? T52 : T5096;
  assign T5096 = io_resetCounts ? 4'h0 : counts_840;
  assign T5097 = T10320 & T5098;
  assign T5098 = T76[10'h348:10'h348];
  assign T11186 = reset ? 4'h0 : T5099;
  assign T5099 = T5101 ? T52 : T5100;
  assign T5100 = io_resetCounts ? 4'h0 : counts_841;
  assign T5101 = T10320 & T5102;
  assign T5102 = T76[10'h349:10'h349];
  assign T5103 = T68[1'h0:1'h0];
  assign T5104 = T5113 ? counts_843 : counts_842;
  assign T11187 = reset ? 4'h0 : T5105;
  assign T5105 = T5107 ? T52 : T5106;
  assign T5106 = io_resetCounts ? 4'h0 : counts_842;
  assign T5107 = T10320 & T5108;
  assign T5108 = T76[10'h34a:10'h34a];
  assign T11188 = reset ? 4'h0 : T5109;
  assign T5109 = T5111 ? T52 : T5110;
  assign T5110 = io_resetCounts ? 4'h0 : counts_843;
  assign T5111 = T10320 & T5112;
  assign T5112 = T76[10'h34b:10'h34b];
  assign T5113 = T68[1'h0:1'h0];
  assign T5114 = T68[1'h1:1'h1];
  assign T5115 = T5136 ? T5126 : T5116;
  assign T5116 = T5125 ? counts_845 : counts_844;
  assign T11189 = reset ? 4'h0 : T5117;
  assign T5117 = T5119 ? T52 : T5118;
  assign T5118 = io_resetCounts ? 4'h0 : counts_844;
  assign T5119 = T10320 & T5120;
  assign T5120 = T76[10'h34c:10'h34c];
  assign T11190 = reset ? 4'h0 : T5121;
  assign T5121 = T5123 ? T52 : T5122;
  assign T5122 = io_resetCounts ? 4'h0 : counts_845;
  assign T5123 = T10320 & T5124;
  assign T5124 = T76[10'h34d:10'h34d];
  assign T5125 = T68[1'h0:1'h0];
  assign T5126 = T5135 ? counts_847 : counts_846;
  assign T11191 = reset ? 4'h0 : T5127;
  assign T5127 = T5129 ? T52 : T5128;
  assign T5128 = io_resetCounts ? 4'h0 : counts_846;
  assign T5129 = T10320 & T5130;
  assign T5130 = T76[10'h34e:10'h34e];
  assign T11192 = reset ? 4'h0 : T5131;
  assign T5131 = T5133 ? T52 : T5132;
  assign T5132 = io_resetCounts ? 4'h0 : counts_847;
  assign T5133 = T10320 & T5134;
  assign T5134 = T76[10'h34f:10'h34f];
  assign T5135 = T68[1'h0:1'h0];
  assign T5136 = T68[1'h1:1'h1];
  assign T5137 = T68[2'h2:2'h2];
  assign T5138 = T68[2'h3:2'h3];
  assign T5139 = T5232 ? T5186 : T5140;
  assign T5140 = T5185 ? T5163 : T5141;
  assign T5141 = T5162 ? T5152 : T5142;
  assign T5142 = T5151 ? counts_849 : counts_848;
  assign T11193 = reset ? 4'h0 : T5143;
  assign T5143 = T5145 ? T52 : T5144;
  assign T5144 = io_resetCounts ? 4'h0 : counts_848;
  assign T5145 = T10320 & T5146;
  assign T5146 = T76[10'h350:10'h350];
  assign T11194 = reset ? 4'h0 : T5147;
  assign T5147 = T5149 ? T52 : T5148;
  assign T5148 = io_resetCounts ? 4'h0 : counts_849;
  assign T5149 = T10320 & T5150;
  assign T5150 = T76[10'h351:10'h351];
  assign T5151 = T68[1'h0:1'h0];
  assign T5152 = T5161 ? counts_851 : counts_850;
  assign T11195 = reset ? 4'h0 : T5153;
  assign T5153 = T5155 ? T52 : T5154;
  assign T5154 = io_resetCounts ? 4'h0 : counts_850;
  assign T5155 = T10320 & T5156;
  assign T5156 = T76[10'h352:10'h352];
  assign T11196 = reset ? 4'h0 : T5157;
  assign T5157 = T5159 ? T52 : T5158;
  assign T5158 = io_resetCounts ? 4'h0 : counts_851;
  assign T5159 = T10320 & T5160;
  assign T5160 = T76[10'h353:10'h353];
  assign T5161 = T68[1'h0:1'h0];
  assign T5162 = T68[1'h1:1'h1];
  assign T5163 = T5184 ? T5174 : T5164;
  assign T5164 = T5173 ? counts_853 : counts_852;
  assign T11197 = reset ? 4'h0 : T5165;
  assign T5165 = T5167 ? T52 : T5166;
  assign T5166 = io_resetCounts ? 4'h0 : counts_852;
  assign T5167 = T10320 & T5168;
  assign T5168 = T76[10'h354:10'h354];
  assign T11198 = reset ? 4'h0 : T5169;
  assign T5169 = T5171 ? T52 : T5170;
  assign T5170 = io_resetCounts ? 4'h0 : counts_853;
  assign T5171 = T10320 & T5172;
  assign T5172 = T76[10'h355:10'h355];
  assign T5173 = T68[1'h0:1'h0];
  assign T5174 = T5183 ? counts_855 : counts_854;
  assign T11199 = reset ? 4'h0 : T5175;
  assign T5175 = T5177 ? T52 : T5176;
  assign T5176 = io_resetCounts ? 4'h0 : counts_854;
  assign T5177 = T10320 & T5178;
  assign T5178 = T76[10'h356:10'h356];
  assign T11200 = reset ? 4'h0 : T5179;
  assign T5179 = T5181 ? T52 : T5180;
  assign T5180 = io_resetCounts ? 4'h0 : counts_855;
  assign T5181 = T10320 & T5182;
  assign T5182 = T76[10'h357:10'h357];
  assign T5183 = T68[1'h0:1'h0];
  assign T5184 = T68[1'h1:1'h1];
  assign T5185 = T68[2'h2:2'h2];
  assign T5186 = T5231 ? T5209 : T5187;
  assign T5187 = T5208 ? T5198 : T5188;
  assign T5188 = T5197 ? counts_857 : counts_856;
  assign T11201 = reset ? 4'h0 : T5189;
  assign T5189 = T5191 ? T52 : T5190;
  assign T5190 = io_resetCounts ? 4'h0 : counts_856;
  assign T5191 = T10320 & T5192;
  assign T5192 = T76[10'h358:10'h358];
  assign T11202 = reset ? 4'h0 : T5193;
  assign T5193 = T5195 ? T52 : T5194;
  assign T5194 = io_resetCounts ? 4'h0 : counts_857;
  assign T5195 = T10320 & T5196;
  assign T5196 = T76[10'h359:10'h359];
  assign T5197 = T68[1'h0:1'h0];
  assign T5198 = T5207 ? counts_859 : counts_858;
  assign T11203 = reset ? 4'h0 : T5199;
  assign T5199 = T5201 ? T52 : T5200;
  assign T5200 = io_resetCounts ? 4'h0 : counts_858;
  assign T5201 = T10320 & T5202;
  assign T5202 = T76[10'h35a:10'h35a];
  assign T11204 = reset ? 4'h0 : T5203;
  assign T5203 = T5205 ? T52 : T5204;
  assign T5204 = io_resetCounts ? 4'h0 : counts_859;
  assign T5205 = T10320 & T5206;
  assign T5206 = T76[10'h35b:10'h35b];
  assign T5207 = T68[1'h0:1'h0];
  assign T5208 = T68[1'h1:1'h1];
  assign T5209 = T5230 ? T5220 : T5210;
  assign T5210 = T5219 ? counts_861 : counts_860;
  assign T11205 = reset ? 4'h0 : T5211;
  assign T5211 = T5213 ? T52 : T5212;
  assign T5212 = io_resetCounts ? 4'h0 : counts_860;
  assign T5213 = T10320 & T5214;
  assign T5214 = T76[10'h35c:10'h35c];
  assign T11206 = reset ? 4'h0 : T5215;
  assign T5215 = T5217 ? T52 : T5216;
  assign T5216 = io_resetCounts ? 4'h0 : counts_861;
  assign T5217 = T10320 & T5218;
  assign T5218 = T76[10'h35d:10'h35d];
  assign T5219 = T68[1'h0:1'h0];
  assign T5220 = T5229 ? counts_863 : counts_862;
  assign T11207 = reset ? 4'h0 : T5221;
  assign T5221 = T5223 ? T52 : T5222;
  assign T5222 = io_resetCounts ? 4'h0 : counts_862;
  assign T5223 = T10320 & T5224;
  assign T5224 = T76[10'h35e:10'h35e];
  assign T11208 = reset ? 4'h0 : T5225;
  assign T5225 = T5227 ? T52 : T5226;
  assign T5226 = io_resetCounts ? 4'h0 : counts_863;
  assign T5227 = T10320 & T5228;
  assign T5228 = T76[10'h35f:10'h35f];
  assign T5229 = T68[1'h0:1'h0];
  assign T5230 = T68[1'h1:1'h1];
  assign T5231 = T68[2'h2:2'h2];
  assign T5232 = T68[2'h3:2'h3];
  assign T5233 = T68[3'h4:3'h4];
  assign T5234 = T5423 ? T5329 : T5235;
  assign T5235 = T5328 ? T5282 : T5236;
  assign T5236 = T5281 ? T5259 : T5237;
  assign T5237 = T5258 ? T5248 : T5238;
  assign T5238 = T5247 ? counts_865 : counts_864;
  assign T11209 = reset ? 4'h0 : T5239;
  assign T5239 = T5241 ? T52 : T5240;
  assign T5240 = io_resetCounts ? 4'h0 : counts_864;
  assign T5241 = T10320 & T5242;
  assign T5242 = T76[10'h360:10'h360];
  assign T11210 = reset ? 4'h0 : T5243;
  assign T5243 = T5245 ? T52 : T5244;
  assign T5244 = io_resetCounts ? 4'h0 : counts_865;
  assign T5245 = T10320 & T5246;
  assign T5246 = T76[10'h361:10'h361];
  assign T5247 = T68[1'h0:1'h0];
  assign T5248 = T5257 ? counts_867 : counts_866;
  assign T11211 = reset ? 4'h0 : T5249;
  assign T5249 = T5251 ? T52 : T5250;
  assign T5250 = io_resetCounts ? 4'h0 : counts_866;
  assign T5251 = T10320 & T5252;
  assign T5252 = T76[10'h362:10'h362];
  assign T11212 = reset ? 4'h0 : T5253;
  assign T5253 = T5255 ? T52 : T5254;
  assign T5254 = io_resetCounts ? 4'h0 : counts_867;
  assign T5255 = T10320 & T5256;
  assign T5256 = T76[10'h363:10'h363];
  assign T5257 = T68[1'h0:1'h0];
  assign T5258 = T68[1'h1:1'h1];
  assign T5259 = T5280 ? T5270 : T5260;
  assign T5260 = T5269 ? counts_869 : counts_868;
  assign T11213 = reset ? 4'h0 : T5261;
  assign T5261 = T5263 ? T52 : T5262;
  assign T5262 = io_resetCounts ? 4'h0 : counts_868;
  assign T5263 = T10320 & T5264;
  assign T5264 = T76[10'h364:10'h364];
  assign T11214 = reset ? 4'h0 : T5265;
  assign T5265 = T5267 ? T52 : T5266;
  assign T5266 = io_resetCounts ? 4'h0 : counts_869;
  assign T5267 = T10320 & T5268;
  assign T5268 = T76[10'h365:10'h365];
  assign T5269 = T68[1'h0:1'h0];
  assign T5270 = T5279 ? counts_871 : counts_870;
  assign T11215 = reset ? 4'h0 : T5271;
  assign T5271 = T5273 ? T52 : T5272;
  assign T5272 = io_resetCounts ? 4'h0 : counts_870;
  assign T5273 = T10320 & T5274;
  assign T5274 = T76[10'h366:10'h366];
  assign T11216 = reset ? 4'h0 : T5275;
  assign T5275 = T5277 ? T52 : T5276;
  assign T5276 = io_resetCounts ? 4'h0 : counts_871;
  assign T5277 = T10320 & T5278;
  assign T5278 = T76[10'h367:10'h367];
  assign T5279 = T68[1'h0:1'h0];
  assign T5280 = T68[1'h1:1'h1];
  assign T5281 = T68[2'h2:2'h2];
  assign T5282 = T5327 ? T5305 : T5283;
  assign T5283 = T5304 ? T5294 : T5284;
  assign T5284 = T5293 ? counts_873 : counts_872;
  assign T11217 = reset ? 4'h0 : T5285;
  assign T5285 = T5287 ? T52 : T5286;
  assign T5286 = io_resetCounts ? 4'h0 : counts_872;
  assign T5287 = T10320 & T5288;
  assign T5288 = T76[10'h368:10'h368];
  assign T11218 = reset ? 4'h0 : T5289;
  assign T5289 = T5291 ? T52 : T5290;
  assign T5290 = io_resetCounts ? 4'h0 : counts_873;
  assign T5291 = T10320 & T5292;
  assign T5292 = T76[10'h369:10'h369];
  assign T5293 = T68[1'h0:1'h0];
  assign T5294 = T5303 ? counts_875 : counts_874;
  assign T11219 = reset ? 4'h0 : T5295;
  assign T5295 = T5297 ? T52 : T5296;
  assign T5296 = io_resetCounts ? 4'h0 : counts_874;
  assign T5297 = T10320 & T5298;
  assign T5298 = T76[10'h36a:10'h36a];
  assign T11220 = reset ? 4'h0 : T5299;
  assign T5299 = T5301 ? T52 : T5300;
  assign T5300 = io_resetCounts ? 4'h0 : counts_875;
  assign T5301 = T10320 & T5302;
  assign T5302 = T76[10'h36b:10'h36b];
  assign T5303 = T68[1'h0:1'h0];
  assign T5304 = T68[1'h1:1'h1];
  assign T5305 = T5326 ? T5316 : T5306;
  assign T5306 = T5315 ? counts_877 : counts_876;
  assign T11221 = reset ? 4'h0 : T5307;
  assign T5307 = T5309 ? T52 : T5308;
  assign T5308 = io_resetCounts ? 4'h0 : counts_876;
  assign T5309 = T10320 & T5310;
  assign T5310 = T76[10'h36c:10'h36c];
  assign T11222 = reset ? 4'h0 : T5311;
  assign T5311 = T5313 ? T52 : T5312;
  assign T5312 = io_resetCounts ? 4'h0 : counts_877;
  assign T5313 = T10320 & T5314;
  assign T5314 = T76[10'h36d:10'h36d];
  assign T5315 = T68[1'h0:1'h0];
  assign T5316 = T5325 ? counts_879 : counts_878;
  assign T11223 = reset ? 4'h0 : T5317;
  assign T5317 = T5319 ? T52 : T5318;
  assign T5318 = io_resetCounts ? 4'h0 : counts_878;
  assign T5319 = T10320 & T5320;
  assign T5320 = T76[10'h36e:10'h36e];
  assign T11224 = reset ? 4'h0 : T5321;
  assign T5321 = T5323 ? T52 : T5322;
  assign T5322 = io_resetCounts ? 4'h0 : counts_879;
  assign T5323 = T10320 & T5324;
  assign T5324 = T76[10'h36f:10'h36f];
  assign T5325 = T68[1'h0:1'h0];
  assign T5326 = T68[1'h1:1'h1];
  assign T5327 = T68[2'h2:2'h2];
  assign T5328 = T68[2'h3:2'h3];
  assign T5329 = T5422 ? T5376 : T5330;
  assign T5330 = T5375 ? T5353 : T5331;
  assign T5331 = T5352 ? T5342 : T5332;
  assign T5332 = T5341 ? counts_881 : counts_880;
  assign T11225 = reset ? 4'h0 : T5333;
  assign T5333 = T5335 ? T52 : T5334;
  assign T5334 = io_resetCounts ? 4'h0 : counts_880;
  assign T5335 = T10320 & T5336;
  assign T5336 = T76[10'h370:10'h370];
  assign T11226 = reset ? 4'h0 : T5337;
  assign T5337 = T5339 ? T52 : T5338;
  assign T5338 = io_resetCounts ? 4'h0 : counts_881;
  assign T5339 = T10320 & T5340;
  assign T5340 = T76[10'h371:10'h371];
  assign T5341 = T68[1'h0:1'h0];
  assign T5342 = T5351 ? counts_883 : counts_882;
  assign T11227 = reset ? 4'h0 : T5343;
  assign T5343 = T5345 ? T52 : T5344;
  assign T5344 = io_resetCounts ? 4'h0 : counts_882;
  assign T5345 = T10320 & T5346;
  assign T5346 = T76[10'h372:10'h372];
  assign T11228 = reset ? 4'h0 : T5347;
  assign T5347 = T5349 ? T52 : T5348;
  assign T5348 = io_resetCounts ? 4'h0 : counts_883;
  assign T5349 = T10320 & T5350;
  assign T5350 = T76[10'h373:10'h373];
  assign T5351 = T68[1'h0:1'h0];
  assign T5352 = T68[1'h1:1'h1];
  assign T5353 = T5374 ? T5364 : T5354;
  assign T5354 = T5363 ? counts_885 : counts_884;
  assign T11229 = reset ? 4'h0 : T5355;
  assign T5355 = T5357 ? T52 : T5356;
  assign T5356 = io_resetCounts ? 4'h0 : counts_884;
  assign T5357 = T10320 & T5358;
  assign T5358 = T76[10'h374:10'h374];
  assign T11230 = reset ? 4'h0 : T5359;
  assign T5359 = T5361 ? T52 : T5360;
  assign T5360 = io_resetCounts ? 4'h0 : counts_885;
  assign T5361 = T10320 & T5362;
  assign T5362 = T76[10'h375:10'h375];
  assign T5363 = T68[1'h0:1'h0];
  assign T5364 = T5373 ? counts_887 : counts_886;
  assign T11231 = reset ? 4'h0 : T5365;
  assign T5365 = T5367 ? T52 : T5366;
  assign T5366 = io_resetCounts ? 4'h0 : counts_886;
  assign T5367 = T10320 & T5368;
  assign T5368 = T76[10'h376:10'h376];
  assign T11232 = reset ? 4'h0 : T5369;
  assign T5369 = T5371 ? T52 : T5370;
  assign T5370 = io_resetCounts ? 4'h0 : counts_887;
  assign T5371 = T10320 & T5372;
  assign T5372 = T76[10'h377:10'h377];
  assign T5373 = T68[1'h0:1'h0];
  assign T5374 = T68[1'h1:1'h1];
  assign T5375 = T68[2'h2:2'h2];
  assign T5376 = T5421 ? T5399 : T5377;
  assign T5377 = T5398 ? T5388 : T5378;
  assign T5378 = T5387 ? counts_889 : counts_888;
  assign T11233 = reset ? 4'h0 : T5379;
  assign T5379 = T5381 ? T52 : T5380;
  assign T5380 = io_resetCounts ? 4'h0 : counts_888;
  assign T5381 = T10320 & T5382;
  assign T5382 = T76[10'h378:10'h378];
  assign T11234 = reset ? 4'h0 : T5383;
  assign T5383 = T5385 ? T52 : T5384;
  assign T5384 = io_resetCounts ? 4'h0 : counts_889;
  assign T5385 = T10320 & T5386;
  assign T5386 = T76[10'h379:10'h379];
  assign T5387 = T68[1'h0:1'h0];
  assign T5388 = T5397 ? counts_891 : counts_890;
  assign T11235 = reset ? 4'h0 : T5389;
  assign T5389 = T5391 ? T52 : T5390;
  assign T5390 = io_resetCounts ? 4'h0 : counts_890;
  assign T5391 = T10320 & T5392;
  assign T5392 = T76[10'h37a:10'h37a];
  assign T11236 = reset ? 4'h0 : T5393;
  assign T5393 = T5395 ? T52 : T5394;
  assign T5394 = io_resetCounts ? 4'h0 : counts_891;
  assign T5395 = T10320 & T5396;
  assign T5396 = T76[10'h37b:10'h37b];
  assign T5397 = T68[1'h0:1'h0];
  assign T5398 = T68[1'h1:1'h1];
  assign T5399 = T5420 ? T5410 : T5400;
  assign T5400 = T5409 ? counts_893 : counts_892;
  assign T11237 = reset ? 4'h0 : T5401;
  assign T5401 = T5403 ? T52 : T5402;
  assign T5402 = io_resetCounts ? 4'h0 : counts_892;
  assign T5403 = T10320 & T5404;
  assign T5404 = T76[10'h37c:10'h37c];
  assign T11238 = reset ? 4'h0 : T5405;
  assign T5405 = T5407 ? T52 : T5406;
  assign T5406 = io_resetCounts ? 4'h0 : counts_893;
  assign T5407 = T10320 & T5408;
  assign T5408 = T76[10'h37d:10'h37d];
  assign T5409 = T68[1'h0:1'h0];
  assign T5410 = T5419 ? counts_895 : counts_894;
  assign T11239 = reset ? 4'h0 : T5411;
  assign T5411 = T5413 ? T52 : T5412;
  assign T5412 = io_resetCounts ? 4'h0 : counts_894;
  assign T5413 = T10320 & T5414;
  assign T5414 = T76[10'h37e:10'h37e];
  assign T11240 = reset ? 4'h0 : T5415;
  assign T5415 = T5417 ? T52 : T5416;
  assign T5416 = io_resetCounts ? 4'h0 : counts_895;
  assign T5417 = T10320 & T5418;
  assign T5418 = T76[10'h37f:10'h37f];
  assign T5419 = T68[1'h0:1'h0];
  assign T5420 = T68[1'h1:1'h1];
  assign T5421 = T68[2'h2:2'h2];
  assign T5422 = T68[2'h3:2'h3];
  assign T5423 = T68[3'h4:3'h4];
  assign T5424 = T68[3'h5:3'h5];
  assign T5425 = T68[3'h6:3'h6];
  assign T5426 = T6191 ? T5809 : T5427;
  assign T5427 = T5808 ? T5618 : T5428;
  assign T5428 = T5617 ? T5523 : T5429;
  assign T5429 = T5522 ? T5476 : T5430;
  assign T5430 = T5475 ? T5453 : T5431;
  assign T5431 = T5452 ? T5442 : T5432;
  assign T5432 = T5441 ? counts_897 : counts_896;
  assign T11241 = reset ? 4'h0 : T5433;
  assign T5433 = T5435 ? T52 : T5434;
  assign T5434 = io_resetCounts ? 4'h0 : counts_896;
  assign T5435 = T10320 & T5436;
  assign T5436 = T76[10'h380:10'h380];
  assign T11242 = reset ? 4'h0 : T5437;
  assign T5437 = T5439 ? T52 : T5438;
  assign T5438 = io_resetCounts ? 4'h0 : counts_897;
  assign T5439 = T10320 & T5440;
  assign T5440 = T76[10'h381:10'h381];
  assign T5441 = T68[1'h0:1'h0];
  assign T5442 = T5451 ? counts_899 : counts_898;
  assign T11243 = reset ? 4'h0 : T5443;
  assign T5443 = T5445 ? T52 : T5444;
  assign T5444 = io_resetCounts ? 4'h0 : counts_898;
  assign T5445 = T10320 & T5446;
  assign T5446 = T76[10'h382:10'h382];
  assign T11244 = reset ? 4'h0 : T5447;
  assign T5447 = T5449 ? T52 : T5448;
  assign T5448 = io_resetCounts ? 4'h0 : counts_899;
  assign T5449 = T10320 & T5450;
  assign T5450 = T76[10'h383:10'h383];
  assign T5451 = T68[1'h0:1'h0];
  assign T5452 = T68[1'h1:1'h1];
  assign T5453 = T5474 ? T5464 : T5454;
  assign T5454 = T5463 ? counts_901 : counts_900;
  assign T11245 = reset ? 4'h0 : T5455;
  assign T5455 = T5457 ? T52 : T5456;
  assign T5456 = io_resetCounts ? 4'h0 : counts_900;
  assign T5457 = T10320 & T5458;
  assign T5458 = T76[10'h384:10'h384];
  assign T11246 = reset ? 4'h0 : T5459;
  assign T5459 = T5461 ? T52 : T5460;
  assign T5460 = io_resetCounts ? 4'h0 : counts_901;
  assign T5461 = T10320 & T5462;
  assign T5462 = T76[10'h385:10'h385];
  assign T5463 = T68[1'h0:1'h0];
  assign T5464 = T5473 ? counts_903 : counts_902;
  assign T11247 = reset ? 4'h0 : T5465;
  assign T5465 = T5467 ? T52 : T5466;
  assign T5466 = io_resetCounts ? 4'h0 : counts_902;
  assign T5467 = T10320 & T5468;
  assign T5468 = T76[10'h386:10'h386];
  assign T11248 = reset ? 4'h0 : T5469;
  assign T5469 = T5471 ? T52 : T5470;
  assign T5470 = io_resetCounts ? 4'h0 : counts_903;
  assign T5471 = T10320 & T5472;
  assign T5472 = T76[10'h387:10'h387];
  assign T5473 = T68[1'h0:1'h0];
  assign T5474 = T68[1'h1:1'h1];
  assign T5475 = T68[2'h2:2'h2];
  assign T5476 = T5521 ? T5499 : T5477;
  assign T5477 = T5498 ? T5488 : T5478;
  assign T5478 = T5487 ? counts_905 : counts_904;
  assign T11249 = reset ? 4'h0 : T5479;
  assign T5479 = T5481 ? T52 : T5480;
  assign T5480 = io_resetCounts ? 4'h0 : counts_904;
  assign T5481 = T10320 & T5482;
  assign T5482 = T76[10'h388:10'h388];
  assign T11250 = reset ? 4'h0 : T5483;
  assign T5483 = T5485 ? T52 : T5484;
  assign T5484 = io_resetCounts ? 4'h0 : counts_905;
  assign T5485 = T10320 & T5486;
  assign T5486 = T76[10'h389:10'h389];
  assign T5487 = T68[1'h0:1'h0];
  assign T5488 = T5497 ? counts_907 : counts_906;
  assign T11251 = reset ? 4'h0 : T5489;
  assign T5489 = T5491 ? T52 : T5490;
  assign T5490 = io_resetCounts ? 4'h0 : counts_906;
  assign T5491 = T10320 & T5492;
  assign T5492 = T76[10'h38a:10'h38a];
  assign T11252 = reset ? 4'h0 : T5493;
  assign T5493 = T5495 ? T52 : T5494;
  assign T5494 = io_resetCounts ? 4'h0 : counts_907;
  assign T5495 = T10320 & T5496;
  assign T5496 = T76[10'h38b:10'h38b];
  assign T5497 = T68[1'h0:1'h0];
  assign T5498 = T68[1'h1:1'h1];
  assign T5499 = T5520 ? T5510 : T5500;
  assign T5500 = T5509 ? counts_909 : counts_908;
  assign T11253 = reset ? 4'h0 : T5501;
  assign T5501 = T5503 ? T52 : T5502;
  assign T5502 = io_resetCounts ? 4'h0 : counts_908;
  assign T5503 = T10320 & T5504;
  assign T5504 = T76[10'h38c:10'h38c];
  assign T11254 = reset ? 4'h0 : T5505;
  assign T5505 = T5507 ? T52 : T5506;
  assign T5506 = io_resetCounts ? 4'h0 : counts_909;
  assign T5507 = T10320 & T5508;
  assign T5508 = T76[10'h38d:10'h38d];
  assign T5509 = T68[1'h0:1'h0];
  assign T5510 = T5519 ? counts_911 : counts_910;
  assign T11255 = reset ? 4'h0 : T5511;
  assign T5511 = T5513 ? T52 : T5512;
  assign T5512 = io_resetCounts ? 4'h0 : counts_910;
  assign T5513 = T10320 & T5514;
  assign T5514 = T76[10'h38e:10'h38e];
  assign T11256 = reset ? 4'h0 : T5515;
  assign T5515 = T5517 ? T52 : T5516;
  assign T5516 = io_resetCounts ? 4'h0 : counts_911;
  assign T5517 = T10320 & T5518;
  assign T5518 = T76[10'h38f:10'h38f];
  assign T5519 = T68[1'h0:1'h0];
  assign T5520 = T68[1'h1:1'h1];
  assign T5521 = T68[2'h2:2'h2];
  assign T5522 = T68[2'h3:2'h3];
  assign T5523 = T5616 ? T5570 : T5524;
  assign T5524 = T5569 ? T5547 : T5525;
  assign T5525 = T5546 ? T5536 : T5526;
  assign T5526 = T5535 ? counts_913 : counts_912;
  assign T11257 = reset ? 4'h0 : T5527;
  assign T5527 = T5529 ? T52 : T5528;
  assign T5528 = io_resetCounts ? 4'h0 : counts_912;
  assign T5529 = T10320 & T5530;
  assign T5530 = T76[10'h390:10'h390];
  assign T11258 = reset ? 4'h0 : T5531;
  assign T5531 = T5533 ? T52 : T5532;
  assign T5532 = io_resetCounts ? 4'h0 : counts_913;
  assign T5533 = T10320 & T5534;
  assign T5534 = T76[10'h391:10'h391];
  assign T5535 = T68[1'h0:1'h0];
  assign T5536 = T5545 ? counts_915 : counts_914;
  assign T11259 = reset ? 4'h0 : T5537;
  assign T5537 = T5539 ? T52 : T5538;
  assign T5538 = io_resetCounts ? 4'h0 : counts_914;
  assign T5539 = T10320 & T5540;
  assign T5540 = T76[10'h392:10'h392];
  assign T11260 = reset ? 4'h0 : T5541;
  assign T5541 = T5543 ? T52 : T5542;
  assign T5542 = io_resetCounts ? 4'h0 : counts_915;
  assign T5543 = T10320 & T5544;
  assign T5544 = T76[10'h393:10'h393];
  assign T5545 = T68[1'h0:1'h0];
  assign T5546 = T68[1'h1:1'h1];
  assign T5547 = T5568 ? T5558 : T5548;
  assign T5548 = T5557 ? counts_917 : counts_916;
  assign T11261 = reset ? 4'h0 : T5549;
  assign T5549 = T5551 ? T52 : T5550;
  assign T5550 = io_resetCounts ? 4'h0 : counts_916;
  assign T5551 = T10320 & T5552;
  assign T5552 = T76[10'h394:10'h394];
  assign T11262 = reset ? 4'h0 : T5553;
  assign T5553 = T5555 ? T52 : T5554;
  assign T5554 = io_resetCounts ? 4'h0 : counts_917;
  assign T5555 = T10320 & T5556;
  assign T5556 = T76[10'h395:10'h395];
  assign T5557 = T68[1'h0:1'h0];
  assign T5558 = T5567 ? counts_919 : counts_918;
  assign T11263 = reset ? 4'h0 : T5559;
  assign T5559 = T5561 ? T52 : T5560;
  assign T5560 = io_resetCounts ? 4'h0 : counts_918;
  assign T5561 = T10320 & T5562;
  assign T5562 = T76[10'h396:10'h396];
  assign T11264 = reset ? 4'h0 : T5563;
  assign T5563 = T5565 ? T52 : T5564;
  assign T5564 = io_resetCounts ? 4'h0 : counts_919;
  assign T5565 = T10320 & T5566;
  assign T5566 = T76[10'h397:10'h397];
  assign T5567 = T68[1'h0:1'h0];
  assign T5568 = T68[1'h1:1'h1];
  assign T5569 = T68[2'h2:2'h2];
  assign T5570 = T5615 ? T5593 : T5571;
  assign T5571 = T5592 ? T5582 : T5572;
  assign T5572 = T5581 ? counts_921 : counts_920;
  assign T11265 = reset ? 4'h0 : T5573;
  assign T5573 = T5575 ? T52 : T5574;
  assign T5574 = io_resetCounts ? 4'h0 : counts_920;
  assign T5575 = T10320 & T5576;
  assign T5576 = T76[10'h398:10'h398];
  assign T11266 = reset ? 4'h0 : T5577;
  assign T5577 = T5579 ? T52 : T5578;
  assign T5578 = io_resetCounts ? 4'h0 : counts_921;
  assign T5579 = T10320 & T5580;
  assign T5580 = T76[10'h399:10'h399];
  assign T5581 = T68[1'h0:1'h0];
  assign T5582 = T5591 ? counts_923 : counts_922;
  assign T11267 = reset ? 4'h0 : T5583;
  assign T5583 = T5585 ? T52 : T5584;
  assign T5584 = io_resetCounts ? 4'h0 : counts_922;
  assign T5585 = T10320 & T5586;
  assign T5586 = T76[10'h39a:10'h39a];
  assign T11268 = reset ? 4'h0 : T5587;
  assign T5587 = T5589 ? T52 : T5588;
  assign T5588 = io_resetCounts ? 4'h0 : counts_923;
  assign T5589 = T10320 & T5590;
  assign T5590 = T76[10'h39b:10'h39b];
  assign T5591 = T68[1'h0:1'h0];
  assign T5592 = T68[1'h1:1'h1];
  assign T5593 = T5614 ? T5604 : T5594;
  assign T5594 = T5603 ? counts_925 : counts_924;
  assign T11269 = reset ? 4'h0 : T5595;
  assign T5595 = T5597 ? T52 : T5596;
  assign T5596 = io_resetCounts ? 4'h0 : counts_924;
  assign T5597 = T10320 & T5598;
  assign T5598 = T76[10'h39c:10'h39c];
  assign T11270 = reset ? 4'h0 : T5599;
  assign T5599 = T5601 ? T52 : T5600;
  assign T5600 = io_resetCounts ? 4'h0 : counts_925;
  assign T5601 = T10320 & T5602;
  assign T5602 = T76[10'h39d:10'h39d];
  assign T5603 = T68[1'h0:1'h0];
  assign T5604 = T5613 ? counts_927 : counts_926;
  assign T11271 = reset ? 4'h0 : T5605;
  assign T5605 = T5607 ? T52 : T5606;
  assign T5606 = io_resetCounts ? 4'h0 : counts_926;
  assign T5607 = T10320 & T5608;
  assign T5608 = T76[10'h39e:10'h39e];
  assign T11272 = reset ? 4'h0 : T5609;
  assign T5609 = T5611 ? T52 : T5610;
  assign T5610 = io_resetCounts ? 4'h0 : counts_927;
  assign T5611 = T10320 & T5612;
  assign T5612 = T76[10'h39f:10'h39f];
  assign T5613 = T68[1'h0:1'h0];
  assign T5614 = T68[1'h1:1'h1];
  assign T5615 = T68[2'h2:2'h2];
  assign T5616 = T68[2'h3:2'h3];
  assign T5617 = T68[3'h4:3'h4];
  assign T5618 = T5807 ? T5713 : T5619;
  assign T5619 = T5712 ? T5666 : T5620;
  assign T5620 = T5665 ? T5643 : T5621;
  assign T5621 = T5642 ? T5632 : T5622;
  assign T5622 = T5631 ? counts_929 : counts_928;
  assign T11273 = reset ? 4'h0 : T5623;
  assign T5623 = T5625 ? T52 : T5624;
  assign T5624 = io_resetCounts ? 4'h0 : counts_928;
  assign T5625 = T10320 & T5626;
  assign T5626 = T76[10'h3a0:10'h3a0];
  assign T11274 = reset ? 4'h0 : T5627;
  assign T5627 = T5629 ? T52 : T5628;
  assign T5628 = io_resetCounts ? 4'h0 : counts_929;
  assign T5629 = T10320 & T5630;
  assign T5630 = T76[10'h3a1:10'h3a1];
  assign T5631 = T68[1'h0:1'h0];
  assign T5632 = T5641 ? counts_931 : counts_930;
  assign T11275 = reset ? 4'h0 : T5633;
  assign T5633 = T5635 ? T52 : T5634;
  assign T5634 = io_resetCounts ? 4'h0 : counts_930;
  assign T5635 = T10320 & T5636;
  assign T5636 = T76[10'h3a2:10'h3a2];
  assign T11276 = reset ? 4'h0 : T5637;
  assign T5637 = T5639 ? T52 : T5638;
  assign T5638 = io_resetCounts ? 4'h0 : counts_931;
  assign T5639 = T10320 & T5640;
  assign T5640 = T76[10'h3a3:10'h3a3];
  assign T5641 = T68[1'h0:1'h0];
  assign T5642 = T68[1'h1:1'h1];
  assign T5643 = T5664 ? T5654 : T5644;
  assign T5644 = T5653 ? counts_933 : counts_932;
  assign T11277 = reset ? 4'h0 : T5645;
  assign T5645 = T5647 ? T52 : T5646;
  assign T5646 = io_resetCounts ? 4'h0 : counts_932;
  assign T5647 = T10320 & T5648;
  assign T5648 = T76[10'h3a4:10'h3a4];
  assign T11278 = reset ? 4'h0 : T5649;
  assign T5649 = T5651 ? T52 : T5650;
  assign T5650 = io_resetCounts ? 4'h0 : counts_933;
  assign T5651 = T10320 & T5652;
  assign T5652 = T76[10'h3a5:10'h3a5];
  assign T5653 = T68[1'h0:1'h0];
  assign T5654 = T5663 ? counts_935 : counts_934;
  assign T11279 = reset ? 4'h0 : T5655;
  assign T5655 = T5657 ? T52 : T5656;
  assign T5656 = io_resetCounts ? 4'h0 : counts_934;
  assign T5657 = T10320 & T5658;
  assign T5658 = T76[10'h3a6:10'h3a6];
  assign T11280 = reset ? 4'h0 : T5659;
  assign T5659 = T5661 ? T52 : T5660;
  assign T5660 = io_resetCounts ? 4'h0 : counts_935;
  assign T5661 = T10320 & T5662;
  assign T5662 = T76[10'h3a7:10'h3a7];
  assign T5663 = T68[1'h0:1'h0];
  assign T5664 = T68[1'h1:1'h1];
  assign T5665 = T68[2'h2:2'h2];
  assign T5666 = T5711 ? T5689 : T5667;
  assign T5667 = T5688 ? T5678 : T5668;
  assign T5668 = T5677 ? counts_937 : counts_936;
  assign T11281 = reset ? 4'h0 : T5669;
  assign T5669 = T5671 ? T52 : T5670;
  assign T5670 = io_resetCounts ? 4'h0 : counts_936;
  assign T5671 = T10320 & T5672;
  assign T5672 = T76[10'h3a8:10'h3a8];
  assign T11282 = reset ? 4'h0 : T5673;
  assign T5673 = T5675 ? T52 : T5674;
  assign T5674 = io_resetCounts ? 4'h0 : counts_937;
  assign T5675 = T10320 & T5676;
  assign T5676 = T76[10'h3a9:10'h3a9];
  assign T5677 = T68[1'h0:1'h0];
  assign T5678 = T5687 ? counts_939 : counts_938;
  assign T11283 = reset ? 4'h0 : T5679;
  assign T5679 = T5681 ? T52 : T5680;
  assign T5680 = io_resetCounts ? 4'h0 : counts_938;
  assign T5681 = T10320 & T5682;
  assign T5682 = T76[10'h3aa:10'h3aa];
  assign T11284 = reset ? 4'h0 : T5683;
  assign T5683 = T5685 ? T52 : T5684;
  assign T5684 = io_resetCounts ? 4'h0 : counts_939;
  assign T5685 = T10320 & T5686;
  assign T5686 = T76[10'h3ab:10'h3ab];
  assign T5687 = T68[1'h0:1'h0];
  assign T5688 = T68[1'h1:1'h1];
  assign T5689 = T5710 ? T5700 : T5690;
  assign T5690 = T5699 ? counts_941 : counts_940;
  assign T11285 = reset ? 4'h0 : T5691;
  assign T5691 = T5693 ? T52 : T5692;
  assign T5692 = io_resetCounts ? 4'h0 : counts_940;
  assign T5693 = T10320 & T5694;
  assign T5694 = T76[10'h3ac:10'h3ac];
  assign T11286 = reset ? 4'h0 : T5695;
  assign T5695 = T5697 ? T52 : T5696;
  assign T5696 = io_resetCounts ? 4'h0 : counts_941;
  assign T5697 = T10320 & T5698;
  assign T5698 = T76[10'h3ad:10'h3ad];
  assign T5699 = T68[1'h0:1'h0];
  assign T5700 = T5709 ? counts_943 : counts_942;
  assign T11287 = reset ? 4'h0 : T5701;
  assign T5701 = T5703 ? T52 : T5702;
  assign T5702 = io_resetCounts ? 4'h0 : counts_942;
  assign T5703 = T10320 & T5704;
  assign T5704 = T76[10'h3ae:10'h3ae];
  assign T11288 = reset ? 4'h0 : T5705;
  assign T5705 = T5707 ? T52 : T5706;
  assign T5706 = io_resetCounts ? 4'h0 : counts_943;
  assign T5707 = T10320 & T5708;
  assign T5708 = T76[10'h3af:10'h3af];
  assign T5709 = T68[1'h0:1'h0];
  assign T5710 = T68[1'h1:1'h1];
  assign T5711 = T68[2'h2:2'h2];
  assign T5712 = T68[2'h3:2'h3];
  assign T5713 = T5806 ? T5760 : T5714;
  assign T5714 = T5759 ? T5737 : T5715;
  assign T5715 = T5736 ? T5726 : T5716;
  assign T5716 = T5725 ? counts_945 : counts_944;
  assign T11289 = reset ? 4'h0 : T5717;
  assign T5717 = T5719 ? T52 : T5718;
  assign T5718 = io_resetCounts ? 4'h0 : counts_944;
  assign T5719 = T10320 & T5720;
  assign T5720 = T76[10'h3b0:10'h3b0];
  assign T11290 = reset ? 4'h0 : T5721;
  assign T5721 = T5723 ? T52 : T5722;
  assign T5722 = io_resetCounts ? 4'h0 : counts_945;
  assign T5723 = T10320 & T5724;
  assign T5724 = T76[10'h3b1:10'h3b1];
  assign T5725 = T68[1'h0:1'h0];
  assign T5726 = T5735 ? counts_947 : counts_946;
  assign T11291 = reset ? 4'h0 : T5727;
  assign T5727 = T5729 ? T52 : T5728;
  assign T5728 = io_resetCounts ? 4'h0 : counts_946;
  assign T5729 = T10320 & T5730;
  assign T5730 = T76[10'h3b2:10'h3b2];
  assign T11292 = reset ? 4'h0 : T5731;
  assign T5731 = T5733 ? T52 : T5732;
  assign T5732 = io_resetCounts ? 4'h0 : counts_947;
  assign T5733 = T10320 & T5734;
  assign T5734 = T76[10'h3b3:10'h3b3];
  assign T5735 = T68[1'h0:1'h0];
  assign T5736 = T68[1'h1:1'h1];
  assign T5737 = T5758 ? T5748 : T5738;
  assign T5738 = T5747 ? counts_949 : counts_948;
  assign T11293 = reset ? 4'h0 : T5739;
  assign T5739 = T5741 ? T52 : T5740;
  assign T5740 = io_resetCounts ? 4'h0 : counts_948;
  assign T5741 = T10320 & T5742;
  assign T5742 = T76[10'h3b4:10'h3b4];
  assign T11294 = reset ? 4'h0 : T5743;
  assign T5743 = T5745 ? T52 : T5744;
  assign T5744 = io_resetCounts ? 4'h0 : counts_949;
  assign T5745 = T10320 & T5746;
  assign T5746 = T76[10'h3b5:10'h3b5];
  assign T5747 = T68[1'h0:1'h0];
  assign T5748 = T5757 ? counts_951 : counts_950;
  assign T11295 = reset ? 4'h0 : T5749;
  assign T5749 = T5751 ? T52 : T5750;
  assign T5750 = io_resetCounts ? 4'h0 : counts_950;
  assign T5751 = T10320 & T5752;
  assign T5752 = T76[10'h3b6:10'h3b6];
  assign T11296 = reset ? 4'h0 : T5753;
  assign T5753 = T5755 ? T52 : T5754;
  assign T5754 = io_resetCounts ? 4'h0 : counts_951;
  assign T5755 = T10320 & T5756;
  assign T5756 = T76[10'h3b7:10'h3b7];
  assign T5757 = T68[1'h0:1'h0];
  assign T5758 = T68[1'h1:1'h1];
  assign T5759 = T68[2'h2:2'h2];
  assign T5760 = T5805 ? T5783 : T5761;
  assign T5761 = T5782 ? T5772 : T5762;
  assign T5762 = T5771 ? counts_953 : counts_952;
  assign T11297 = reset ? 4'h0 : T5763;
  assign T5763 = T5765 ? T52 : T5764;
  assign T5764 = io_resetCounts ? 4'h0 : counts_952;
  assign T5765 = T10320 & T5766;
  assign T5766 = T76[10'h3b8:10'h3b8];
  assign T11298 = reset ? 4'h0 : T5767;
  assign T5767 = T5769 ? T52 : T5768;
  assign T5768 = io_resetCounts ? 4'h0 : counts_953;
  assign T5769 = T10320 & T5770;
  assign T5770 = T76[10'h3b9:10'h3b9];
  assign T5771 = T68[1'h0:1'h0];
  assign T5772 = T5781 ? counts_955 : counts_954;
  assign T11299 = reset ? 4'h0 : T5773;
  assign T5773 = T5775 ? T52 : T5774;
  assign T5774 = io_resetCounts ? 4'h0 : counts_954;
  assign T5775 = T10320 & T5776;
  assign T5776 = T76[10'h3ba:10'h3ba];
  assign T11300 = reset ? 4'h0 : T5777;
  assign T5777 = T5779 ? T52 : T5778;
  assign T5778 = io_resetCounts ? 4'h0 : counts_955;
  assign T5779 = T10320 & T5780;
  assign T5780 = T76[10'h3bb:10'h3bb];
  assign T5781 = T68[1'h0:1'h0];
  assign T5782 = T68[1'h1:1'h1];
  assign T5783 = T5804 ? T5794 : T5784;
  assign T5784 = T5793 ? counts_957 : counts_956;
  assign T11301 = reset ? 4'h0 : T5785;
  assign T5785 = T5787 ? T52 : T5786;
  assign T5786 = io_resetCounts ? 4'h0 : counts_956;
  assign T5787 = T10320 & T5788;
  assign T5788 = T76[10'h3bc:10'h3bc];
  assign T11302 = reset ? 4'h0 : T5789;
  assign T5789 = T5791 ? T52 : T5790;
  assign T5790 = io_resetCounts ? 4'h0 : counts_957;
  assign T5791 = T10320 & T5792;
  assign T5792 = T76[10'h3bd:10'h3bd];
  assign T5793 = T68[1'h0:1'h0];
  assign T5794 = T5803 ? counts_959 : counts_958;
  assign T11303 = reset ? 4'h0 : T5795;
  assign T5795 = T5797 ? T52 : T5796;
  assign T5796 = io_resetCounts ? 4'h0 : counts_958;
  assign T5797 = T10320 & T5798;
  assign T5798 = T76[10'h3be:10'h3be];
  assign T11304 = reset ? 4'h0 : T5799;
  assign T5799 = T5801 ? T52 : T5800;
  assign T5800 = io_resetCounts ? 4'h0 : counts_959;
  assign T5801 = T10320 & T5802;
  assign T5802 = T76[10'h3bf:10'h3bf];
  assign T5803 = T68[1'h0:1'h0];
  assign T5804 = T68[1'h1:1'h1];
  assign T5805 = T68[2'h2:2'h2];
  assign T5806 = T68[2'h3:2'h3];
  assign T5807 = T68[3'h4:3'h4];
  assign T5808 = T68[3'h5:3'h5];
  assign T5809 = T6190 ? T6000 : T5810;
  assign T5810 = T5999 ? T5905 : T5811;
  assign T5811 = T5904 ? T5858 : T5812;
  assign T5812 = T5857 ? T5835 : T5813;
  assign T5813 = T5834 ? T5824 : T5814;
  assign T5814 = T5823 ? counts_961 : counts_960;
  assign T11305 = reset ? 4'h0 : T5815;
  assign T5815 = T5817 ? T52 : T5816;
  assign T5816 = io_resetCounts ? 4'h0 : counts_960;
  assign T5817 = T10320 & T5818;
  assign T5818 = T76[10'h3c0:10'h3c0];
  assign T11306 = reset ? 4'h0 : T5819;
  assign T5819 = T5821 ? T52 : T5820;
  assign T5820 = io_resetCounts ? 4'h0 : counts_961;
  assign T5821 = T10320 & T5822;
  assign T5822 = T76[10'h3c1:10'h3c1];
  assign T5823 = T68[1'h0:1'h0];
  assign T5824 = T5833 ? counts_963 : counts_962;
  assign T11307 = reset ? 4'h0 : T5825;
  assign T5825 = T5827 ? T52 : T5826;
  assign T5826 = io_resetCounts ? 4'h0 : counts_962;
  assign T5827 = T10320 & T5828;
  assign T5828 = T76[10'h3c2:10'h3c2];
  assign T11308 = reset ? 4'h0 : T5829;
  assign T5829 = T5831 ? T52 : T5830;
  assign T5830 = io_resetCounts ? 4'h0 : counts_963;
  assign T5831 = T10320 & T5832;
  assign T5832 = T76[10'h3c3:10'h3c3];
  assign T5833 = T68[1'h0:1'h0];
  assign T5834 = T68[1'h1:1'h1];
  assign T5835 = T5856 ? T5846 : T5836;
  assign T5836 = T5845 ? counts_965 : counts_964;
  assign T11309 = reset ? 4'h0 : T5837;
  assign T5837 = T5839 ? T52 : T5838;
  assign T5838 = io_resetCounts ? 4'h0 : counts_964;
  assign T5839 = T10320 & T5840;
  assign T5840 = T76[10'h3c4:10'h3c4];
  assign T11310 = reset ? 4'h0 : T5841;
  assign T5841 = T5843 ? T52 : T5842;
  assign T5842 = io_resetCounts ? 4'h0 : counts_965;
  assign T5843 = T10320 & T5844;
  assign T5844 = T76[10'h3c5:10'h3c5];
  assign T5845 = T68[1'h0:1'h0];
  assign T5846 = T5855 ? counts_967 : counts_966;
  assign T11311 = reset ? 4'h0 : T5847;
  assign T5847 = T5849 ? T52 : T5848;
  assign T5848 = io_resetCounts ? 4'h0 : counts_966;
  assign T5849 = T10320 & T5850;
  assign T5850 = T76[10'h3c6:10'h3c6];
  assign T11312 = reset ? 4'h0 : T5851;
  assign T5851 = T5853 ? T52 : T5852;
  assign T5852 = io_resetCounts ? 4'h0 : counts_967;
  assign T5853 = T10320 & T5854;
  assign T5854 = T76[10'h3c7:10'h3c7];
  assign T5855 = T68[1'h0:1'h0];
  assign T5856 = T68[1'h1:1'h1];
  assign T5857 = T68[2'h2:2'h2];
  assign T5858 = T5903 ? T5881 : T5859;
  assign T5859 = T5880 ? T5870 : T5860;
  assign T5860 = T5869 ? counts_969 : counts_968;
  assign T11313 = reset ? 4'h0 : T5861;
  assign T5861 = T5863 ? T52 : T5862;
  assign T5862 = io_resetCounts ? 4'h0 : counts_968;
  assign T5863 = T10320 & T5864;
  assign T5864 = T76[10'h3c8:10'h3c8];
  assign T11314 = reset ? 4'h0 : T5865;
  assign T5865 = T5867 ? T52 : T5866;
  assign T5866 = io_resetCounts ? 4'h0 : counts_969;
  assign T5867 = T10320 & T5868;
  assign T5868 = T76[10'h3c9:10'h3c9];
  assign T5869 = T68[1'h0:1'h0];
  assign T5870 = T5879 ? counts_971 : counts_970;
  assign T11315 = reset ? 4'h0 : T5871;
  assign T5871 = T5873 ? T52 : T5872;
  assign T5872 = io_resetCounts ? 4'h0 : counts_970;
  assign T5873 = T10320 & T5874;
  assign T5874 = T76[10'h3ca:10'h3ca];
  assign T11316 = reset ? 4'h0 : T5875;
  assign T5875 = T5877 ? T52 : T5876;
  assign T5876 = io_resetCounts ? 4'h0 : counts_971;
  assign T5877 = T10320 & T5878;
  assign T5878 = T76[10'h3cb:10'h3cb];
  assign T5879 = T68[1'h0:1'h0];
  assign T5880 = T68[1'h1:1'h1];
  assign T5881 = T5902 ? T5892 : T5882;
  assign T5882 = T5891 ? counts_973 : counts_972;
  assign T11317 = reset ? 4'h0 : T5883;
  assign T5883 = T5885 ? T52 : T5884;
  assign T5884 = io_resetCounts ? 4'h0 : counts_972;
  assign T5885 = T10320 & T5886;
  assign T5886 = T76[10'h3cc:10'h3cc];
  assign T11318 = reset ? 4'h0 : T5887;
  assign T5887 = T5889 ? T52 : T5888;
  assign T5888 = io_resetCounts ? 4'h0 : counts_973;
  assign T5889 = T10320 & T5890;
  assign T5890 = T76[10'h3cd:10'h3cd];
  assign T5891 = T68[1'h0:1'h0];
  assign T5892 = T5901 ? counts_975 : counts_974;
  assign T11319 = reset ? 4'h0 : T5893;
  assign T5893 = T5895 ? T52 : T5894;
  assign T5894 = io_resetCounts ? 4'h0 : counts_974;
  assign T5895 = T10320 & T5896;
  assign T5896 = T76[10'h3ce:10'h3ce];
  assign T11320 = reset ? 4'h0 : T5897;
  assign T5897 = T5899 ? T52 : T5898;
  assign T5898 = io_resetCounts ? 4'h0 : counts_975;
  assign T5899 = T10320 & T5900;
  assign T5900 = T76[10'h3cf:10'h3cf];
  assign T5901 = T68[1'h0:1'h0];
  assign T5902 = T68[1'h1:1'h1];
  assign T5903 = T68[2'h2:2'h2];
  assign T5904 = T68[2'h3:2'h3];
  assign T5905 = T5998 ? T5952 : T5906;
  assign T5906 = T5951 ? T5929 : T5907;
  assign T5907 = T5928 ? T5918 : T5908;
  assign T5908 = T5917 ? counts_977 : counts_976;
  assign T11321 = reset ? 4'h0 : T5909;
  assign T5909 = T5911 ? T52 : T5910;
  assign T5910 = io_resetCounts ? 4'h0 : counts_976;
  assign T5911 = T10320 & T5912;
  assign T5912 = T76[10'h3d0:10'h3d0];
  assign T11322 = reset ? 4'h0 : T5913;
  assign T5913 = T5915 ? T52 : T5914;
  assign T5914 = io_resetCounts ? 4'h0 : counts_977;
  assign T5915 = T10320 & T5916;
  assign T5916 = T76[10'h3d1:10'h3d1];
  assign T5917 = T68[1'h0:1'h0];
  assign T5918 = T5927 ? counts_979 : counts_978;
  assign T11323 = reset ? 4'h0 : T5919;
  assign T5919 = T5921 ? T52 : T5920;
  assign T5920 = io_resetCounts ? 4'h0 : counts_978;
  assign T5921 = T10320 & T5922;
  assign T5922 = T76[10'h3d2:10'h3d2];
  assign T11324 = reset ? 4'h0 : T5923;
  assign T5923 = T5925 ? T52 : T5924;
  assign T5924 = io_resetCounts ? 4'h0 : counts_979;
  assign T5925 = T10320 & T5926;
  assign T5926 = T76[10'h3d3:10'h3d3];
  assign T5927 = T68[1'h0:1'h0];
  assign T5928 = T68[1'h1:1'h1];
  assign T5929 = T5950 ? T5940 : T5930;
  assign T5930 = T5939 ? counts_981 : counts_980;
  assign T11325 = reset ? 4'h0 : T5931;
  assign T5931 = T5933 ? T52 : T5932;
  assign T5932 = io_resetCounts ? 4'h0 : counts_980;
  assign T5933 = T10320 & T5934;
  assign T5934 = T76[10'h3d4:10'h3d4];
  assign T11326 = reset ? 4'h0 : T5935;
  assign T5935 = T5937 ? T52 : T5936;
  assign T5936 = io_resetCounts ? 4'h0 : counts_981;
  assign T5937 = T10320 & T5938;
  assign T5938 = T76[10'h3d5:10'h3d5];
  assign T5939 = T68[1'h0:1'h0];
  assign T5940 = T5949 ? counts_983 : counts_982;
  assign T11327 = reset ? 4'h0 : T5941;
  assign T5941 = T5943 ? T52 : T5942;
  assign T5942 = io_resetCounts ? 4'h0 : counts_982;
  assign T5943 = T10320 & T5944;
  assign T5944 = T76[10'h3d6:10'h3d6];
  assign T11328 = reset ? 4'h0 : T5945;
  assign T5945 = T5947 ? T52 : T5946;
  assign T5946 = io_resetCounts ? 4'h0 : counts_983;
  assign T5947 = T10320 & T5948;
  assign T5948 = T76[10'h3d7:10'h3d7];
  assign T5949 = T68[1'h0:1'h0];
  assign T5950 = T68[1'h1:1'h1];
  assign T5951 = T68[2'h2:2'h2];
  assign T5952 = T5997 ? T5975 : T5953;
  assign T5953 = T5974 ? T5964 : T5954;
  assign T5954 = T5963 ? counts_985 : counts_984;
  assign T11329 = reset ? 4'h0 : T5955;
  assign T5955 = T5957 ? T52 : T5956;
  assign T5956 = io_resetCounts ? 4'h0 : counts_984;
  assign T5957 = T10320 & T5958;
  assign T5958 = T76[10'h3d8:10'h3d8];
  assign T11330 = reset ? 4'h0 : T5959;
  assign T5959 = T5961 ? T52 : T5960;
  assign T5960 = io_resetCounts ? 4'h0 : counts_985;
  assign T5961 = T10320 & T5962;
  assign T5962 = T76[10'h3d9:10'h3d9];
  assign T5963 = T68[1'h0:1'h0];
  assign T5964 = T5973 ? counts_987 : counts_986;
  assign T11331 = reset ? 4'h0 : T5965;
  assign T5965 = T5967 ? T52 : T5966;
  assign T5966 = io_resetCounts ? 4'h0 : counts_986;
  assign T5967 = T10320 & T5968;
  assign T5968 = T76[10'h3da:10'h3da];
  assign T11332 = reset ? 4'h0 : T5969;
  assign T5969 = T5971 ? T52 : T5970;
  assign T5970 = io_resetCounts ? 4'h0 : counts_987;
  assign T5971 = T10320 & T5972;
  assign T5972 = T76[10'h3db:10'h3db];
  assign T5973 = T68[1'h0:1'h0];
  assign T5974 = T68[1'h1:1'h1];
  assign T5975 = T5996 ? T5986 : T5976;
  assign T5976 = T5985 ? counts_989 : counts_988;
  assign T11333 = reset ? 4'h0 : T5977;
  assign T5977 = T5979 ? T52 : T5978;
  assign T5978 = io_resetCounts ? 4'h0 : counts_988;
  assign T5979 = T10320 & T5980;
  assign T5980 = T76[10'h3dc:10'h3dc];
  assign T11334 = reset ? 4'h0 : T5981;
  assign T5981 = T5983 ? T52 : T5982;
  assign T5982 = io_resetCounts ? 4'h0 : counts_989;
  assign T5983 = T10320 & T5984;
  assign T5984 = T76[10'h3dd:10'h3dd];
  assign T5985 = T68[1'h0:1'h0];
  assign T5986 = T5995 ? counts_991 : counts_990;
  assign T11335 = reset ? 4'h0 : T5987;
  assign T5987 = T5989 ? T52 : T5988;
  assign T5988 = io_resetCounts ? 4'h0 : counts_990;
  assign T5989 = T10320 & T5990;
  assign T5990 = T76[10'h3de:10'h3de];
  assign T11336 = reset ? 4'h0 : T5991;
  assign T5991 = T5993 ? T52 : T5992;
  assign T5992 = io_resetCounts ? 4'h0 : counts_991;
  assign T5993 = T10320 & T5994;
  assign T5994 = T76[10'h3df:10'h3df];
  assign T5995 = T68[1'h0:1'h0];
  assign T5996 = T68[1'h1:1'h1];
  assign T5997 = T68[2'h2:2'h2];
  assign T5998 = T68[2'h3:2'h3];
  assign T5999 = T68[3'h4:3'h4];
  assign T6000 = T6189 ? T6095 : T6001;
  assign T6001 = T6094 ? T6048 : T6002;
  assign T6002 = T6047 ? T6025 : T6003;
  assign T6003 = T6024 ? T6014 : T6004;
  assign T6004 = T6013 ? counts_993 : counts_992;
  assign T11337 = reset ? 4'h0 : T6005;
  assign T6005 = T6007 ? T52 : T6006;
  assign T6006 = io_resetCounts ? 4'h0 : counts_992;
  assign T6007 = T10320 & T6008;
  assign T6008 = T76[10'h3e0:10'h3e0];
  assign T11338 = reset ? 4'h0 : T6009;
  assign T6009 = T6011 ? T52 : T6010;
  assign T6010 = io_resetCounts ? 4'h0 : counts_993;
  assign T6011 = T10320 & T6012;
  assign T6012 = T76[10'h3e1:10'h3e1];
  assign T6013 = T68[1'h0:1'h0];
  assign T6014 = T6023 ? counts_995 : counts_994;
  assign T11339 = reset ? 4'h0 : T6015;
  assign T6015 = T6017 ? T52 : T6016;
  assign T6016 = io_resetCounts ? 4'h0 : counts_994;
  assign T6017 = T10320 & T6018;
  assign T6018 = T76[10'h3e2:10'h3e2];
  assign T11340 = reset ? 4'h0 : T6019;
  assign T6019 = T6021 ? T52 : T6020;
  assign T6020 = io_resetCounts ? 4'h0 : counts_995;
  assign T6021 = T10320 & T6022;
  assign T6022 = T76[10'h3e3:10'h3e3];
  assign T6023 = T68[1'h0:1'h0];
  assign T6024 = T68[1'h1:1'h1];
  assign T6025 = T6046 ? T6036 : T6026;
  assign T6026 = T6035 ? counts_997 : counts_996;
  assign T11341 = reset ? 4'h0 : T6027;
  assign T6027 = T6029 ? T52 : T6028;
  assign T6028 = io_resetCounts ? 4'h0 : counts_996;
  assign T6029 = T10320 & T6030;
  assign T6030 = T76[10'h3e4:10'h3e4];
  assign T11342 = reset ? 4'h0 : T6031;
  assign T6031 = T6033 ? T52 : T6032;
  assign T6032 = io_resetCounts ? 4'h0 : counts_997;
  assign T6033 = T10320 & T6034;
  assign T6034 = T76[10'h3e5:10'h3e5];
  assign T6035 = T68[1'h0:1'h0];
  assign T6036 = T6045 ? counts_999 : counts_998;
  assign T11343 = reset ? 4'h0 : T6037;
  assign T6037 = T6039 ? T52 : T6038;
  assign T6038 = io_resetCounts ? 4'h0 : counts_998;
  assign T6039 = T10320 & T6040;
  assign T6040 = T76[10'h3e6:10'h3e6];
  assign T11344 = reset ? 4'h0 : T6041;
  assign T6041 = T6043 ? T52 : T6042;
  assign T6042 = io_resetCounts ? 4'h0 : counts_999;
  assign T6043 = T10320 & T6044;
  assign T6044 = T76[10'h3e7:10'h3e7];
  assign T6045 = T68[1'h0:1'h0];
  assign T6046 = T68[1'h1:1'h1];
  assign T6047 = T68[2'h2:2'h2];
  assign T6048 = T6093 ? T6071 : T6049;
  assign T6049 = T6070 ? T6060 : T6050;
  assign T6050 = T6059 ? counts_1001 : counts_1000;
  assign T11345 = reset ? 4'h0 : T6051;
  assign T6051 = T6053 ? T52 : T6052;
  assign T6052 = io_resetCounts ? 4'h0 : counts_1000;
  assign T6053 = T10320 & T6054;
  assign T6054 = T76[10'h3e8:10'h3e8];
  assign T11346 = reset ? 4'h0 : T6055;
  assign T6055 = T6057 ? T52 : T6056;
  assign T6056 = io_resetCounts ? 4'h0 : counts_1001;
  assign T6057 = T10320 & T6058;
  assign T6058 = T76[10'h3e9:10'h3e9];
  assign T6059 = T68[1'h0:1'h0];
  assign T6060 = T6069 ? counts_1003 : counts_1002;
  assign T11347 = reset ? 4'h0 : T6061;
  assign T6061 = T6063 ? T52 : T6062;
  assign T6062 = io_resetCounts ? 4'h0 : counts_1002;
  assign T6063 = T10320 & T6064;
  assign T6064 = T76[10'h3ea:10'h3ea];
  assign T11348 = reset ? 4'h0 : T6065;
  assign T6065 = T6067 ? T52 : T6066;
  assign T6066 = io_resetCounts ? 4'h0 : counts_1003;
  assign T6067 = T10320 & T6068;
  assign T6068 = T76[10'h3eb:10'h3eb];
  assign T6069 = T68[1'h0:1'h0];
  assign T6070 = T68[1'h1:1'h1];
  assign T6071 = T6092 ? T6082 : T6072;
  assign T6072 = T6081 ? counts_1005 : counts_1004;
  assign T11349 = reset ? 4'h0 : T6073;
  assign T6073 = T6075 ? T52 : T6074;
  assign T6074 = io_resetCounts ? 4'h0 : counts_1004;
  assign T6075 = T10320 & T6076;
  assign T6076 = T76[10'h3ec:10'h3ec];
  assign T11350 = reset ? 4'h0 : T6077;
  assign T6077 = T6079 ? T52 : T6078;
  assign T6078 = io_resetCounts ? 4'h0 : counts_1005;
  assign T6079 = T10320 & T6080;
  assign T6080 = T76[10'h3ed:10'h3ed];
  assign T6081 = T68[1'h0:1'h0];
  assign T6082 = T6091 ? counts_1007 : counts_1006;
  assign T11351 = reset ? 4'h0 : T6083;
  assign T6083 = T6085 ? T52 : T6084;
  assign T6084 = io_resetCounts ? 4'h0 : counts_1006;
  assign T6085 = T10320 & T6086;
  assign T6086 = T76[10'h3ee:10'h3ee];
  assign T11352 = reset ? 4'h0 : T6087;
  assign T6087 = T6089 ? T52 : T6088;
  assign T6088 = io_resetCounts ? 4'h0 : counts_1007;
  assign T6089 = T10320 & T6090;
  assign T6090 = T76[10'h3ef:10'h3ef];
  assign T6091 = T68[1'h0:1'h0];
  assign T6092 = T68[1'h1:1'h1];
  assign T6093 = T68[2'h2:2'h2];
  assign T6094 = T68[2'h3:2'h3];
  assign T6095 = T6188 ? T6142 : T6096;
  assign T6096 = T6141 ? T6119 : T6097;
  assign T6097 = T6118 ? T6108 : T6098;
  assign T6098 = T6107 ? counts_1009 : counts_1008;
  assign T11353 = reset ? 4'h0 : T6099;
  assign T6099 = T6101 ? T52 : T6100;
  assign T6100 = io_resetCounts ? 4'h0 : counts_1008;
  assign T6101 = T10320 & T6102;
  assign T6102 = T76[10'h3f0:10'h3f0];
  assign T11354 = reset ? 4'h0 : T6103;
  assign T6103 = T6105 ? T52 : T6104;
  assign T6104 = io_resetCounts ? 4'h0 : counts_1009;
  assign T6105 = T10320 & T6106;
  assign T6106 = T76[10'h3f1:10'h3f1];
  assign T6107 = T68[1'h0:1'h0];
  assign T6108 = T6117 ? counts_1011 : counts_1010;
  assign T11355 = reset ? 4'h0 : T6109;
  assign T6109 = T6111 ? T52 : T6110;
  assign T6110 = io_resetCounts ? 4'h0 : counts_1010;
  assign T6111 = T10320 & T6112;
  assign T6112 = T76[10'h3f2:10'h3f2];
  assign T11356 = reset ? 4'h0 : T6113;
  assign T6113 = T6115 ? T52 : T6114;
  assign T6114 = io_resetCounts ? 4'h0 : counts_1011;
  assign T6115 = T10320 & T6116;
  assign T6116 = T76[10'h3f3:10'h3f3];
  assign T6117 = T68[1'h0:1'h0];
  assign T6118 = T68[1'h1:1'h1];
  assign T6119 = T6140 ? T6130 : T6120;
  assign T6120 = T6129 ? counts_1013 : counts_1012;
  assign T11357 = reset ? 4'h0 : T6121;
  assign T6121 = T6123 ? T52 : T6122;
  assign T6122 = io_resetCounts ? 4'h0 : counts_1012;
  assign T6123 = T10320 & T6124;
  assign T6124 = T76[10'h3f4:10'h3f4];
  assign T11358 = reset ? 4'h0 : T6125;
  assign T6125 = T6127 ? T52 : T6126;
  assign T6126 = io_resetCounts ? 4'h0 : counts_1013;
  assign T6127 = T10320 & T6128;
  assign T6128 = T76[10'h3f5:10'h3f5];
  assign T6129 = T68[1'h0:1'h0];
  assign T6130 = T6139 ? counts_1015 : counts_1014;
  assign T11359 = reset ? 4'h0 : T6131;
  assign T6131 = T6133 ? T52 : T6132;
  assign T6132 = io_resetCounts ? 4'h0 : counts_1014;
  assign T6133 = T10320 & T6134;
  assign T6134 = T76[10'h3f6:10'h3f6];
  assign T11360 = reset ? 4'h0 : T6135;
  assign T6135 = T6137 ? T52 : T6136;
  assign T6136 = io_resetCounts ? 4'h0 : counts_1015;
  assign T6137 = T10320 & T6138;
  assign T6138 = T76[10'h3f7:10'h3f7];
  assign T6139 = T68[1'h0:1'h0];
  assign T6140 = T68[1'h1:1'h1];
  assign T6141 = T68[2'h2:2'h2];
  assign T6142 = T6187 ? T6165 : T6143;
  assign T6143 = T6164 ? T6154 : T6144;
  assign T6144 = T6153 ? counts_1017 : counts_1016;
  assign T11361 = reset ? 4'h0 : T6145;
  assign T6145 = T6147 ? T52 : T6146;
  assign T6146 = io_resetCounts ? 4'h0 : counts_1016;
  assign T6147 = T10320 & T6148;
  assign T6148 = T76[10'h3f8:10'h3f8];
  assign T11362 = reset ? 4'h0 : T6149;
  assign T6149 = T6151 ? T52 : T6150;
  assign T6150 = io_resetCounts ? 4'h0 : counts_1017;
  assign T6151 = T10320 & T6152;
  assign T6152 = T76[10'h3f9:10'h3f9];
  assign T6153 = T68[1'h0:1'h0];
  assign T6154 = T6163 ? counts_1019 : counts_1018;
  assign T11363 = reset ? 4'h0 : T6155;
  assign T6155 = T6157 ? T52 : T6156;
  assign T6156 = io_resetCounts ? 4'h0 : counts_1018;
  assign T6157 = T10320 & T6158;
  assign T6158 = T76[10'h3fa:10'h3fa];
  assign T11364 = reset ? 4'h0 : T6159;
  assign T6159 = T6161 ? T52 : T6160;
  assign T6160 = io_resetCounts ? 4'h0 : counts_1019;
  assign T6161 = T10320 & T6162;
  assign T6162 = T76[10'h3fb:10'h3fb];
  assign T6163 = T68[1'h0:1'h0];
  assign T6164 = T68[1'h1:1'h1];
  assign T6165 = T6186 ? T6176 : T6166;
  assign T6166 = T6175 ? counts_1021 : counts_1020;
  assign T11365 = reset ? 4'h0 : T6167;
  assign T6167 = T6169 ? T52 : T6168;
  assign T6168 = io_resetCounts ? 4'h0 : counts_1020;
  assign T6169 = T10320 & T6170;
  assign T6170 = T76[10'h3fc:10'h3fc];
  assign T11366 = reset ? 4'h0 : T6171;
  assign T6171 = T6173 ? T52 : T6172;
  assign T6172 = io_resetCounts ? 4'h0 : counts_1021;
  assign T6173 = T10320 & T6174;
  assign T6174 = T76[10'h3fd:10'h3fd];
  assign T6175 = T68[1'h0:1'h0];
  assign T6176 = T6185 ? counts_1023 : counts_1022;
  assign T11367 = reset ? 4'h0 : T6177;
  assign T6177 = T6179 ? T52 : T6178;
  assign T6178 = io_resetCounts ? 4'h0 : counts_1022;
  assign T6179 = T10320 & T6180;
  assign T6180 = T76[10'h3fe:10'h3fe];
  assign T11368 = reset ? 4'h0 : T6181;
  assign T6181 = T6183 ? T52 : T6182;
  assign T6182 = io_resetCounts ? 4'h0 : counts_1023;
  assign T6183 = T10320 & T6184;
  assign T6184 = T76[10'h3ff:10'h3ff];
  assign T6185 = T68[1'h0:1'h0];
  assign T6186 = T68[1'h1:1'h1];
  assign T6187 = T68[2'h2:2'h2];
  assign T6188 = T68[2'h3:2'h3];
  assign T6189 = T68[3'h4:3'h4];
  assign T6190 = T68[3'h5:3'h5];
  assign T6191 = T68[3'h6:3'h6];
  assign T6192 = T68[3'h7:3'h7];
  assign T6193 = T68[4'h8:4'h8];
  assign T6194 = T68[4'h9:4'h9];
  assign T6195 = T55[2'h3:1'h0];
  assign T6196 = T10320 & T6197;
  assign T6197 = T76[1'h0:1'h0];
  assign T11369 = reset ? 4'h0 : T6198;
  assign T6198 = T6200 ? T52 : T6199;
  assign T6199 = io_resetCounts ? 4'h0 : counts_1;
  assign T6200 = T10320 & T6201;
  assign T6201 = T76[1'h1:1'h1];
  assign T6202 = T6203[1'h0:1'h0];
  assign T6203 = curInfo_hash2;
  assign T6204 = T6205 ? counts_3 : counts_2;
  assign T6205 = T6203[1'h0:1'h0];
  assign T6206 = T6203[1'h1:1'h1];
  assign T6207 = T6212 ? T6210 : T6208;
  assign T6208 = T6209 ? counts_5 : counts_4;
  assign T6209 = T6203[1'h0:1'h0];
  assign T6210 = T6211 ? counts_7 : counts_6;
  assign T6211 = T6203[1'h0:1'h0];
  assign T6212 = T6203[1'h1:1'h1];
  assign T6213 = T6203[2'h2:2'h2];
  assign T6214 = T6227 ? T6221 : T6215;
  assign T6215 = T6220 ? T6218 : T6216;
  assign T6216 = T6217 ? counts_9 : counts_8;
  assign T6217 = T6203[1'h0:1'h0];
  assign T6218 = T6219 ? counts_11 : counts_10;
  assign T6219 = T6203[1'h0:1'h0];
  assign T6220 = T6203[1'h1:1'h1];
  assign T6221 = T6226 ? T6224 : T6222;
  assign T6222 = T6223 ? counts_13 : counts_12;
  assign T6223 = T6203[1'h0:1'h0];
  assign T6224 = T6225 ? counts_15 : counts_14;
  assign T6225 = T6203[1'h0:1'h0];
  assign T6226 = T6203[1'h1:1'h1];
  assign T6227 = T6203[2'h2:2'h2];
  assign T6228 = T6203[2'h3:2'h3];
  assign T6229 = T6258 ? T6244 : T6230;
  assign T6230 = T6243 ? T6237 : T6231;
  assign T6231 = T6236 ? T6234 : T6232;
  assign T6232 = T6233 ? counts_17 : counts_16;
  assign T6233 = T6203[1'h0:1'h0];
  assign T6234 = T6235 ? counts_19 : counts_18;
  assign T6235 = T6203[1'h0:1'h0];
  assign T6236 = T6203[1'h1:1'h1];
  assign T6237 = T6242 ? T6240 : T6238;
  assign T6238 = T6239 ? counts_21 : counts_20;
  assign T6239 = T6203[1'h0:1'h0];
  assign T6240 = T6241 ? counts_23 : counts_22;
  assign T6241 = T6203[1'h0:1'h0];
  assign T6242 = T6203[1'h1:1'h1];
  assign T6243 = T6203[2'h2:2'h2];
  assign T6244 = T6257 ? T6251 : T6245;
  assign T6245 = T6250 ? T6248 : T6246;
  assign T6246 = T6247 ? counts_25 : counts_24;
  assign T6247 = T6203[1'h0:1'h0];
  assign T6248 = T6249 ? counts_27 : counts_26;
  assign T6249 = T6203[1'h0:1'h0];
  assign T6250 = T6203[1'h1:1'h1];
  assign T6251 = T6256 ? T6254 : T6252;
  assign T6252 = T6253 ? counts_29 : counts_28;
  assign T6253 = T6203[1'h0:1'h0];
  assign T6254 = T6255 ? counts_31 : counts_30;
  assign T6255 = T6203[1'h0:1'h0];
  assign T6256 = T6203[1'h1:1'h1];
  assign T6257 = T6203[2'h2:2'h2];
  assign T6258 = T6203[2'h3:2'h3];
  assign T6259 = T6203[3'h4:3'h4];
  assign T6260 = T6321 ? T6291 : T6261;
  assign T6261 = T6290 ? T6276 : T6262;
  assign T6262 = T6275 ? T6269 : T6263;
  assign T6263 = T6268 ? T6266 : T6264;
  assign T6264 = T6265 ? counts_33 : counts_32;
  assign T6265 = T6203[1'h0:1'h0];
  assign T6266 = T6267 ? counts_35 : counts_34;
  assign T6267 = T6203[1'h0:1'h0];
  assign T6268 = T6203[1'h1:1'h1];
  assign T6269 = T6274 ? T6272 : T6270;
  assign T6270 = T6271 ? counts_37 : counts_36;
  assign T6271 = T6203[1'h0:1'h0];
  assign T6272 = T6273 ? counts_39 : counts_38;
  assign T6273 = T6203[1'h0:1'h0];
  assign T6274 = T6203[1'h1:1'h1];
  assign T6275 = T6203[2'h2:2'h2];
  assign T6276 = T6289 ? T6283 : T6277;
  assign T6277 = T6282 ? T6280 : T6278;
  assign T6278 = T6279 ? counts_41 : counts_40;
  assign T6279 = T6203[1'h0:1'h0];
  assign T6280 = T6281 ? counts_43 : counts_42;
  assign T6281 = T6203[1'h0:1'h0];
  assign T6282 = T6203[1'h1:1'h1];
  assign T6283 = T6288 ? T6286 : T6284;
  assign T6284 = T6285 ? counts_45 : counts_44;
  assign T6285 = T6203[1'h0:1'h0];
  assign T6286 = T6287 ? counts_47 : counts_46;
  assign T6287 = T6203[1'h0:1'h0];
  assign T6288 = T6203[1'h1:1'h1];
  assign T6289 = T6203[2'h2:2'h2];
  assign T6290 = T6203[2'h3:2'h3];
  assign T6291 = T6320 ? T6306 : T6292;
  assign T6292 = T6305 ? T6299 : T6293;
  assign T6293 = T6298 ? T6296 : T6294;
  assign T6294 = T6295 ? counts_49 : counts_48;
  assign T6295 = T6203[1'h0:1'h0];
  assign T6296 = T6297 ? counts_51 : counts_50;
  assign T6297 = T6203[1'h0:1'h0];
  assign T6298 = T6203[1'h1:1'h1];
  assign T6299 = T6304 ? T6302 : T6300;
  assign T6300 = T6301 ? counts_53 : counts_52;
  assign T6301 = T6203[1'h0:1'h0];
  assign T6302 = T6303 ? counts_55 : counts_54;
  assign T6303 = T6203[1'h0:1'h0];
  assign T6304 = T6203[1'h1:1'h1];
  assign T6305 = T6203[2'h2:2'h2];
  assign T6306 = T6319 ? T6313 : T6307;
  assign T6307 = T6312 ? T6310 : T6308;
  assign T6308 = T6309 ? counts_57 : counts_56;
  assign T6309 = T6203[1'h0:1'h0];
  assign T6310 = T6311 ? counts_59 : counts_58;
  assign T6311 = T6203[1'h0:1'h0];
  assign T6312 = T6203[1'h1:1'h1];
  assign T6313 = T6318 ? T6316 : T6314;
  assign T6314 = T6315 ? counts_61 : counts_60;
  assign T6315 = T6203[1'h0:1'h0];
  assign T6316 = T6317 ? counts_63 : counts_62;
  assign T6317 = T6203[1'h0:1'h0];
  assign T6318 = T6203[1'h1:1'h1];
  assign T6319 = T6203[2'h2:2'h2];
  assign T6320 = T6203[2'h3:2'h3];
  assign T6321 = T6203[3'h4:3'h4];
  assign T6322 = T6203[3'h5:3'h5];
  assign T6323 = T6448 ? T6386 : T6324;
  assign T6324 = T6385 ? T6355 : T6325;
  assign T6325 = T6354 ? T6340 : T6326;
  assign T6326 = T6339 ? T6333 : T6327;
  assign T6327 = T6332 ? T6330 : T6328;
  assign T6328 = T6329 ? counts_65 : counts_64;
  assign T6329 = T6203[1'h0:1'h0];
  assign T6330 = T6331 ? counts_67 : counts_66;
  assign T6331 = T6203[1'h0:1'h0];
  assign T6332 = T6203[1'h1:1'h1];
  assign T6333 = T6338 ? T6336 : T6334;
  assign T6334 = T6335 ? counts_69 : counts_68;
  assign T6335 = T6203[1'h0:1'h0];
  assign T6336 = T6337 ? counts_71 : counts_70;
  assign T6337 = T6203[1'h0:1'h0];
  assign T6338 = T6203[1'h1:1'h1];
  assign T6339 = T6203[2'h2:2'h2];
  assign T6340 = T6353 ? T6347 : T6341;
  assign T6341 = T6346 ? T6344 : T6342;
  assign T6342 = T6343 ? counts_73 : counts_72;
  assign T6343 = T6203[1'h0:1'h0];
  assign T6344 = T6345 ? counts_75 : counts_74;
  assign T6345 = T6203[1'h0:1'h0];
  assign T6346 = T6203[1'h1:1'h1];
  assign T6347 = T6352 ? T6350 : T6348;
  assign T6348 = T6349 ? counts_77 : counts_76;
  assign T6349 = T6203[1'h0:1'h0];
  assign T6350 = T6351 ? counts_79 : counts_78;
  assign T6351 = T6203[1'h0:1'h0];
  assign T6352 = T6203[1'h1:1'h1];
  assign T6353 = T6203[2'h2:2'h2];
  assign T6354 = T6203[2'h3:2'h3];
  assign T6355 = T6384 ? T6370 : T6356;
  assign T6356 = T6369 ? T6363 : T6357;
  assign T6357 = T6362 ? T6360 : T6358;
  assign T6358 = T6359 ? counts_81 : counts_80;
  assign T6359 = T6203[1'h0:1'h0];
  assign T6360 = T6361 ? counts_83 : counts_82;
  assign T6361 = T6203[1'h0:1'h0];
  assign T6362 = T6203[1'h1:1'h1];
  assign T6363 = T6368 ? T6366 : T6364;
  assign T6364 = T6365 ? counts_85 : counts_84;
  assign T6365 = T6203[1'h0:1'h0];
  assign T6366 = T6367 ? counts_87 : counts_86;
  assign T6367 = T6203[1'h0:1'h0];
  assign T6368 = T6203[1'h1:1'h1];
  assign T6369 = T6203[2'h2:2'h2];
  assign T6370 = T6383 ? T6377 : T6371;
  assign T6371 = T6376 ? T6374 : T6372;
  assign T6372 = T6373 ? counts_89 : counts_88;
  assign T6373 = T6203[1'h0:1'h0];
  assign T6374 = T6375 ? counts_91 : counts_90;
  assign T6375 = T6203[1'h0:1'h0];
  assign T6376 = T6203[1'h1:1'h1];
  assign T6377 = T6382 ? T6380 : T6378;
  assign T6378 = T6379 ? counts_93 : counts_92;
  assign T6379 = T6203[1'h0:1'h0];
  assign T6380 = T6381 ? counts_95 : counts_94;
  assign T6381 = T6203[1'h0:1'h0];
  assign T6382 = T6203[1'h1:1'h1];
  assign T6383 = T6203[2'h2:2'h2];
  assign T6384 = T6203[2'h3:2'h3];
  assign T6385 = T6203[3'h4:3'h4];
  assign T6386 = T6447 ? T6417 : T6387;
  assign T6387 = T6416 ? T6402 : T6388;
  assign T6388 = T6401 ? T6395 : T6389;
  assign T6389 = T6394 ? T6392 : T6390;
  assign T6390 = T6391 ? counts_97 : counts_96;
  assign T6391 = T6203[1'h0:1'h0];
  assign T6392 = T6393 ? counts_99 : counts_98;
  assign T6393 = T6203[1'h0:1'h0];
  assign T6394 = T6203[1'h1:1'h1];
  assign T6395 = T6400 ? T6398 : T6396;
  assign T6396 = T6397 ? counts_101 : counts_100;
  assign T6397 = T6203[1'h0:1'h0];
  assign T6398 = T6399 ? counts_103 : counts_102;
  assign T6399 = T6203[1'h0:1'h0];
  assign T6400 = T6203[1'h1:1'h1];
  assign T6401 = T6203[2'h2:2'h2];
  assign T6402 = T6415 ? T6409 : T6403;
  assign T6403 = T6408 ? T6406 : T6404;
  assign T6404 = T6405 ? counts_105 : counts_104;
  assign T6405 = T6203[1'h0:1'h0];
  assign T6406 = T6407 ? counts_107 : counts_106;
  assign T6407 = T6203[1'h0:1'h0];
  assign T6408 = T6203[1'h1:1'h1];
  assign T6409 = T6414 ? T6412 : T6410;
  assign T6410 = T6411 ? counts_109 : counts_108;
  assign T6411 = T6203[1'h0:1'h0];
  assign T6412 = T6413 ? counts_111 : counts_110;
  assign T6413 = T6203[1'h0:1'h0];
  assign T6414 = T6203[1'h1:1'h1];
  assign T6415 = T6203[2'h2:2'h2];
  assign T6416 = T6203[2'h3:2'h3];
  assign T6417 = T6446 ? T6432 : T6418;
  assign T6418 = T6431 ? T6425 : T6419;
  assign T6419 = T6424 ? T6422 : T6420;
  assign T6420 = T6421 ? counts_113 : counts_112;
  assign T6421 = T6203[1'h0:1'h0];
  assign T6422 = T6423 ? counts_115 : counts_114;
  assign T6423 = T6203[1'h0:1'h0];
  assign T6424 = T6203[1'h1:1'h1];
  assign T6425 = T6430 ? T6428 : T6426;
  assign T6426 = T6427 ? counts_117 : counts_116;
  assign T6427 = T6203[1'h0:1'h0];
  assign T6428 = T6429 ? counts_119 : counts_118;
  assign T6429 = T6203[1'h0:1'h0];
  assign T6430 = T6203[1'h1:1'h1];
  assign T6431 = T6203[2'h2:2'h2];
  assign T6432 = T6445 ? T6439 : T6433;
  assign T6433 = T6438 ? T6436 : T6434;
  assign T6434 = T6435 ? counts_121 : counts_120;
  assign T6435 = T6203[1'h0:1'h0];
  assign T6436 = T6437 ? counts_123 : counts_122;
  assign T6437 = T6203[1'h0:1'h0];
  assign T6438 = T6203[1'h1:1'h1];
  assign T6439 = T6444 ? T6442 : T6440;
  assign T6440 = T6441 ? counts_125 : counts_124;
  assign T6441 = T6203[1'h0:1'h0];
  assign T6442 = T6443 ? counts_127 : counts_126;
  assign T6443 = T6203[1'h0:1'h0];
  assign T6444 = T6203[1'h1:1'h1];
  assign T6445 = T6203[2'h2:2'h2];
  assign T6446 = T6203[2'h3:2'h3];
  assign T6447 = T6203[3'h4:3'h4];
  assign T6448 = T6203[3'h5:3'h5];
  assign T6449 = T6203[3'h6:3'h6];
  assign T6450 = T6703 ? T6577 : T6451;
  assign T6451 = T6576 ? T6514 : T6452;
  assign T6452 = T6513 ? T6483 : T6453;
  assign T6453 = T6482 ? T6468 : T6454;
  assign T6454 = T6467 ? T6461 : T6455;
  assign T6455 = T6460 ? T6458 : T6456;
  assign T6456 = T6457 ? counts_129 : counts_128;
  assign T6457 = T6203[1'h0:1'h0];
  assign T6458 = T6459 ? counts_131 : counts_130;
  assign T6459 = T6203[1'h0:1'h0];
  assign T6460 = T6203[1'h1:1'h1];
  assign T6461 = T6466 ? T6464 : T6462;
  assign T6462 = T6463 ? counts_133 : counts_132;
  assign T6463 = T6203[1'h0:1'h0];
  assign T6464 = T6465 ? counts_135 : counts_134;
  assign T6465 = T6203[1'h0:1'h0];
  assign T6466 = T6203[1'h1:1'h1];
  assign T6467 = T6203[2'h2:2'h2];
  assign T6468 = T6481 ? T6475 : T6469;
  assign T6469 = T6474 ? T6472 : T6470;
  assign T6470 = T6471 ? counts_137 : counts_136;
  assign T6471 = T6203[1'h0:1'h0];
  assign T6472 = T6473 ? counts_139 : counts_138;
  assign T6473 = T6203[1'h0:1'h0];
  assign T6474 = T6203[1'h1:1'h1];
  assign T6475 = T6480 ? T6478 : T6476;
  assign T6476 = T6477 ? counts_141 : counts_140;
  assign T6477 = T6203[1'h0:1'h0];
  assign T6478 = T6479 ? counts_143 : counts_142;
  assign T6479 = T6203[1'h0:1'h0];
  assign T6480 = T6203[1'h1:1'h1];
  assign T6481 = T6203[2'h2:2'h2];
  assign T6482 = T6203[2'h3:2'h3];
  assign T6483 = T6512 ? T6498 : T6484;
  assign T6484 = T6497 ? T6491 : T6485;
  assign T6485 = T6490 ? T6488 : T6486;
  assign T6486 = T6487 ? counts_145 : counts_144;
  assign T6487 = T6203[1'h0:1'h0];
  assign T6488 = T6489 ? counts_147 : counts_146;
  assign T6489 = T6203[1'h0:1'h0];
  assign T6490 = T6203[1'h1:1'h1];
  assign T6491 = T6496 ? T6494 : T6492;
  assign T6492 = T6493 ? counts_149 : counts_148;
  assign T6493 = T6203[1'h0:1'h0];
  assign T6494 = T6495 ? counts_151 : counts_150;
  assign T6495 = T6203[1'h0:1'h0];
  assign T6496 = T6203[1'h1:1'h1];
  assign T6497 = T6203[2'h2:2'h2];
  assign T6498 = T6511 ? T6505 : T6499;
  assign T6499 = T6504 ? T6502 : T6500;
  assign T6500 = T6501 ? counts_153 : counts_152;
  assign T6501 = T6203[1'h0:1'h0];
  assign T6502 = T6503 ? counts_155 : counts_154;
  assign T6503 = T6203[1'h0:1'h0];
  assign T6504 = T6203[1'h1:1'h1];
  assign T6505 = T6510 ? T6508 : T6506;
  assign T6506 = T6507 ? counts_157 : counts_156;
  assign T6507 = T6203[1'h0:1'h0];
  assign T6508 = T6509 ? counts_159 : counts_158;
  assign T6509 = T6203[1'h0:1'h0];
  assign T6510 = T6203[1'h1:1'h1];
  assign T6511 = T6203[2'h2:2'h2];
  assign T6512 = T6203[2'h3:2'h3];
  assign T6513 = T6203[3'h4:3'h4];
  assign T6514 = T6575 ? T6545 : T6515;
  assign T6515 = T6544 ? T6530 : T6516;
  assign T6516 = T6529 ? T6523 : T6517;
  assign T6517 = T6522 ? T6520 : T6518;
  assign T6518 = T6519 ? counts_161 : counts_160;
  assign T6519 = T6203[1'h0:1'h0];
  assign T6520 = T6521 ? counts_163 : counts_162;
  assign T6521 = T6203[1'h0:1'h0];
  assign T6522 = T6203[1'h1:1'h1];
  assign T6523 = T6528 ? T6526 : T6524;
  assign T6524 = T6525 ? counts_165 : counts_164;
  assign T6525 = T6203[1'h0:1'h0];
  assign T6526 = T6527 ? counts_167 : counts_166;
  assign T6527 = T6203[1'h0:1'h0];
  assign T6528 = T6203[1'h1:1'h1];
  assign T6529 = T6203[2'h2:2'h2];
  assign T6530 = T6543 ? T6537 : T6531;
  assign T6531 = T6536 ? T6534 : T6532;
  assign T6532 = T6533 ? counts_169 : counts_168;
  assign T6533 = T6203[1'h0:1'h0];
  assign T6534 = T6535 ? counts_171 : counts_170;
  assign T6535 = T6203[1'h0:1'h0];
  assign T6536 = T6203[1'h1:1'h1];
  assign T6537 = T6542 ? T6540 : T6538;
  assign T6538 = T6539 ? counts_173 : counts_172;
  assign T6539 = T6203[1'h0:1'h0];
  assign T6540 = T6541 ? counts_175 : counts_174;
  assign T6541 = T6203[1'h0:1'h0];
  assign T6542 = T6203[1'h1:1'h1];
  assign T6543 = T6203[2'h2:2'h2];
  assign T6544 = T6203[2'h3:2'h3];
  assign T6545 = T6574 ? T6560 : T6546;
  assign T6546 = T6559 ? T6553 : T6547;
  assign T6547 = T6552 ? T6550 : T6548;
  assign T6548 = T6549 ? counts_177 : counts_176;
  assign T6549 = T6203[1'h0:1'h0];
  assign T6550 = T6551 ? counts_179 : counts_178;
  assign T6551 = T6203[1'h0:1'h0];
  assign T6552 = T6203[1'h1:1'h1];
  assign T6553 = T6558 ? T6556 : T6554;
  assign T6554 = T6555 ? counts_181 : counts_180;
  assign T6555 = T6203[1'h0:1'h0];
  assign T6556 = T6557 ? counts_183 : counts_182;
  assign T6557 = T6203[1'h0:1'h0];
  assign T6558 = T6203[1'h1:1'h1];
  assign T6559 = T6203[2'h2:2'h2];
  assign T6560 = T6573 ? T6567 : T6561;
  assign T6561 = T6566 ? T6564 : T6562;
  assign T6562 = T6563 ? counts_185 : counts_184;
  assign T6563 = T6203[1'h0:1'h0];
  assign T6564 = T6565 ? counts_187 : counts_186;
  assign T6565 = T6203[1'h0:1'h0];
  assign T6566 = T6203[1'h1:1'h1];
  assign T6567 = T6572 ? T6570 : T6568;
  assign T6568 = T6569 ? counts_189 : counts_188;
  assign T6569 = T6203[1'h0:1'h0];
  assign T6570 = T6571 ? counts_191 : counts_190;
  assign T6571 = T6203[1'h0:1'h0];
  assign T6572 = T6203[1'h1:1'h1];
  assign T6573 = T6203[2'h2:2'h2];
  assign T6574 = T6203[2'h3:2'h3];
  assign T6575 = T6203[3'h4:3'h4];
  assign T6576 = T6203[3'h5:3'h5];
  assign T6577 = T6702 ? T6640 : T6578;
  assign T6578 = T6639 ? T6609 : T6579;
  assign T6579 = T6608 ? T6594 : T6580;
  assign T6580 = T6593 ? T6587 : T6581;
  assign T6581 = T6586 ? T6584 : T6582;
  assign T6582 = T6583 ? counts_193 : counts_192;
  assign T6583 = T6203[1'h0:1'h0];
  assign T6584 = T6585 ? counts_195 : counts_194;
  assign T6585 = T6203[1'h0:1'h0];
  assign T6586 = T6203[1'h1:1'h1];
  assign T6587 = T6592 ? T6590 : T6588;
  assign T6588 = T6589 ? counts_197 : counts_196;
  assign T6589 = T6203[1'h0:1'h0];
  assign T6590 = T6591 ? counts_199 : counts_198;
  assign T6591 = T6203[1'h0:1'h0];
  assign T6592 = T6203[1'h1:1'h1];
  assign T6593 = T6203[2'h2:2'h2];
  assign T6594 = T6607 ? T6601 : T6595;
  assign T6595 = T6600 ? T6598 : T6596;
  assign T6596 = T6597 ? counts_201 : counts_200;
  assign T6597 = T6203[1'h0:1'h0];
  assign T6598 = T6599 ? counts_203 : counts_202;
  assign T6599 = T6203[1'h0:1'h0];
  assign T6600 = T6203[1'h1:1'h1];
  assign T6601 = T6606 ? T6604 : T6602;
  assign T6602 = T6603 ? counts_205 : counts_204;
  assign T6603 = T6203[1'h0:1'h0];
  assign T6604 = T6605 ? counts_207 : counts_206;
  assign T6605 = T6203[1'h0:1'h0];
  assign T6606 = T6203[1'h1:1'h1];
  assign T6607 = T6203[2'h2:2'h2];
  assign T6608 = T6203[2'h3:2'h3];
  assign T6609 = T6638 ? T6624 : T6610;
  assign T6610 = T6623 ? T6617 : T6611;
  assign T6611 = T6616 ? T6614 : T6612;
  assign T6612 = T6613 ? counts_209 : counts_208;
  assign T6613 = T6203[1'h0:1'h0];
  assign T6614 = T6615 ? counts_211 : counts_210;
  assign T6615 = T6203[1'h0:1'h0];
  assign T6616 = T6203[1'h1:1'h1];
  assign T6617 = T6622 ? T6620 : T6618;
  assign T6618 = T6619 ? counts_213 : counts_212;
  assign T6619 = T6203[1'h0:1'h0];
  assign T6620 = T6621 ? counts_215 : counts_214;
  assign T6621 = T6203[1'h0:1'h0];
  assign T6622 = T6203[1'h1:1'h1];
  assign T6623 = T6203[2'h2:2'h2];
  assign T6624 = T6637 ? T6631 : T6625;
  assign T6625 = T6630 ? T6628 : T6626;
  assign T6626 = T6627 ? counts_217 : counts_216;
  assign T6627 = T6203[1'h0:1'h0];
  assign T6628 = T6629 ? counts_219 : counts_218;
  assign T6629 = T6203[1'h0:1'h0];
  assign T6630 = T6203[1'h1:1'h1];
  assign T6631 = T6636 ? T6634 : T6632;
  assign T6632 = T6633 ? counts_221 : counts_220;
  assign T6633 = T6203[1'h0:1'h0];
  assign T6634 = T6635 ? counts_223 : counts_222;
  assign T6635 = T6203[1'h0:1'h0];
  assign T6636 = T6203[1'h1:1'h1];
  assign T6637 = T6203[2'h2:2'h2];
  assign T6638 = T6203[2'h3:2'h3];
  assign T6639 = T6203[3'h4:3'h4];
  assign T6640 = T6701 ? T6671 : T6641;
  assign T6641 = T6670 ? T6656 : T6642;
  assign T6642 = T6655 ? T6649 : T6643;
  assign T6643 = T6648 ? T6646 : T6644;
  assign T6644 = T6645 ? counts_225 : counts_224;
  assign T6645 = T6203[1'h0:1'h0];
  assign T6646 = T6647 ? counts_227 : counts_226;
  assign T6647 = T6203[1'h0:1'h0];
  assign T6648 = T6203[1'h1:1'h1];
  assign T6649 = T6654 ? T6652 : T6650;
  assign T6650 = T6651 ? counts_229 : counts_228;
  assign T6651 = T6203[1'h0:1'h0];
  assign T6652 = T6653 ? counts_231 : counts_230;
  assign T6653 = T6203[1'h0:1'h0];
  assign T6654 = T6203[1'h1:1'h1];
  assign T6655 = T6203[2'h2:2'h2];
  assign T6656 = T6669 ? T6663 : T6657;
  assign T6657 = T6662 ? T6660 : T6658;
  assign T6658 = T6659 ? counts_233 : counts_232;
  assign T6659 = T6203[1'h0:1'h0];
  assign T6660 = T6661 ? counts_235 : counts_234;
  assign T6661 = T6203[1'h0:1'h0];
  assign T6662 = T6203[1'h1:1'h1];
  assign T6663 = T6668 ? T6666 : T6664;
  assign T6664 = T6665 ? counts_237 : counts_236;
  assign T6665 = T6203[1'h0:1'h0];
  assign T6666 = T6667 ? counts_239 : counts_238;
  assign T6667 = T6203[1'h0:1'h0];
  assign T6668 = T6203[1'h1:1'h1];
  assign T6669 = T6203[2'h2:2'h2];
  assign T6670 = T6203[2'h3:2'h3];
  assign T6671 = T6700 ? T6686 : T6672;
  assign T6672 = T6685 ? T6679 : T6673;
  assign T6673 = T6678 ? T6676 : T6674;
  assign T6674 = T6675 ? counts_241 : counts_240;
  assign T6675 = T6203[1'h0:1'h0];
  assign T6676 = T6677 ? counts_243 : counts_242;
  assign T6677 = T6203[1'h0:1'h0];
  assign T6678 = T6203[1'h1:1'h1];
  assign T6679 = T6684 ? T6682 : T6680;
  assign T6680 = T6681 ? counts_245 : counts_244;
  assign T6681 = T6203[1'h0:1'h0];
  assign T6682 = T6683 ? counts_247 : counts_246;
  assign T6683 = T6203[1'h0:1'h0];
  assign T6684 = T6203[1'h1:1'h1];
  assign T6685 = T6203[2'h2:2'h2];
  assign T6686 = T6699 ? T6693 : T6687;
  assign T6687 = T6692 ? T6690 : T6688;
  assign T6688 = T6689 ? counts_249 : counts_248;
  assign T6689 = T6203[1'h0:1'h0];
  assign T6690 = T6691 ? counts_251 : counts_250;
  assign T6691 = T6203[1'h0:1'h0];
  assign T6692 = T6203[1'h1:1'h1];
  assign T6693 = T6698 ? T6696 : T6694;
  assign T6694 = T6695 ? counts_253 : counts_252;
  assign T6695 = T6203[1'h0:1'h0];
  assign T6696 = T6697 ? counts_255 : counts_254;
  assign T6697 = T6203[1'h0:1'h0];
  assign T6698 = T6203[1'h1:1'h1];
  assign T6699 = T6203[2'h2:2'h2];
  assign T6700 = T6203[2'h3:2'h3];
  assign T6701 = T6203[3'h4:3'h4];
  assign T6702 = T6203[3'h5:3'h5];
  assign T6703 = T6203[3'h6:3'h6];
  assign T6704 = T6203[3'h7:3'h7];
  assign T6705 = T7214 ? T6960 : T6706;
  assign T6706 = T6959 ? T6833 : T6707;
  assign T6707 = T6832 ? T6770 : T6708;
  assign T6708 = T6769 ? T6739 : T6709;
  assign T6709 = T6738 ? T6724 : T6710;
  assign T6710 = T6723 ? T6717 : T6711;
  assign T6711 = T6716 ? T6714 : T6712;
  assign T6712 = T6713 ? counts_257 : counts_256;
  assign T6713 = T6203[1'h0:1'h0];
  assign T6714 = T6715 ? counts_259 : counts_258;
  assign T6715 = T6203[1'h0:1'h0];
  assign T6716 = T6203[1'h1:1'h1];
  assign T6717 = T6722 ? T6720 : T6718;
  assign T6718 = T6719 ? counts_261 : counts_260;
  assign T6719 = T6203[1'h0:1'h0];
  assign T6720 = T6721 ? counts_263 : counts_262;
  assign T6721 = T6203[1'h0:1'h0];
  assign T6722 = T6203[1'h1:1'h1];
  assign T6723 = T6203[2'h2:2'h2];
  assign T6724 = T6737 ? T6731 : T6725;
  assign T6725 = T6730 ? T6728 : T6726;
  assign T6726 = T6727 ? counts_265 : counts_264;
  assign T6727 = T6203[1'h0:1'h0];
  assign T6728 = T6729 ? counts_267 : counts_266;
  assign T6729 = T6203[1'h0:1'h0];
  assign T6730 = T6203[1'h1:1'h1];
  assign T6731 = T6736 ? T6734 : T6732;
  assign T6732 = T6733 ? counts_269 : counts_268;
  assign T6733 = T6203[1'h0:1'h0];
  assign T6734 = T6735 ? counts_271 : counts_270;
  assign T6735 = T6203[1'h0:1'h0];
  assign T6736 = T6203[1'h1:1'h1];
  assign T6737 = T6203[2'h2:2'h2];
  assign T6738 = T6203[2'h3:2'h3];
  assign T6739 = T6768 ? T6754 : T6740;
  assign T6740 = T6753 ? T6747 : T6741;
  assign T6741 = T6746 ? T6744 : T6742;
  assign T6742 = T6743 ? counts_273 : counts_272;
  assign T6743 = T6203[1'h0:1'h0];
  assign T6744 = T6745 ? counts_275 : counts_274;
  assign T6745 = T6203[1'h0:1'h0];
  assign T6746 = T6203[1'h1:1'h1];
  assign T6747 = T6752 ? T6750 : T6748;
  assign T6748 = T6749 ? counts_277 : counts_276;
  assign T6749 = T6203[1'h0:1'h0];
  assign T6750 = T6751 ? counts_279 : counts_278;
  assign T6751 = T6203[1'h0:1'h0];
  assign T6752 = T6203[1'h1:1'h1];
  assign T6753 = T6203[2'h2:2'h2];
  assign T6754 = T6767 ? T6761 : T6755;
  assign T6755 = T6760 ? T6758 : T6756;
  assign T6756 = T6757 ? counts_281 : counts_280;
  assign T6757 = T6203[1'h0:1'h0];
  assign T6758 = T6759 ? counts_283 : counts_282;
  assign T6759 = T6203[1'h0:1'h0];
  assign T6760 = T6203[1'h1:1'h1];
  assign T6761 = T6766 ? T6764 : T6762;
  assign T6762 = T6763 ? counts_285 : counts_284;
  assign T6763 = T6203[1'h0:1'h0];
  assign T6764 = T6765 ? counts_287 : counts_286;
  assign T6765 = T6203[1'h0:1'h0];
  assign T6766 = T6203[1'h1:1'h1];
  assign T6767 = T6203[2'h2:2'h2];
  assign T6768 = T6203[2'h3:2'h3];
  assign T6769 = T6203[3'h4:3'h4];
  assign T6770 = T6831 ? T6801 : T6771;
  assign T6771 = T6800 ? T6786 : T6772;
  assign T6772 = T6785 ? T6779 : T6773;
  assign T6773 = T6778 ? T6776 : T6774;
  assign T6774 = T6775 ? counts_289 : counts_288;
  assign T6775 = T6203[1'h0:1'h0];
  assign T6776 = T6777 ? counts_291 : counts_290;
  assign T6777 = T6203[1'h0:1'h0];
  assign T6778 = T6203[1'h1:1'h1];
  assign T6779 = T6784 ? T6782 : T6780;
  assign T6780 = T6781 ? counts_293 : counts_292;
  assign T6781 = T6203[1'h0:1'h0];
  assign T6782 = T6783 ? counts_295 : counts_294;
  assign T6783 = T6203[1'h0:1'h0];
  assign T6784 = T6203[1'h1:1'h1];
  assign T6785 = T6203[2'h2:2'h2];
  assign T6786 = T6799 ? T6793 : T6787;
  assign T6787 = T6792 ? T6790 : T6788;
  assign T6788 = T6789 ? counts_297 : counts_296;
  assign T6789 = T6203[1'h0:1'h0];
  assign T6790 = T6791 ? counts_299 : counts_298;
  assign T6791 = T6203[1'h0:1'h0];
  assign T6792 = T6203[1'h1:1'h1];
  assign T6793 = T6798 ? T6796 : T6794;
  assign T6794 = T6795 ? counts_301 : counts_300;
  assign T6795 = T6203[1'h0:1'h0];
  assign T6796 = T6797 ? counts_303 : counts_302;
  assign T6797 = T6203[1'h0:1'h0];
  assign T6798 = T6203[1'h1:1'h1];
  assign T6799 = T6203[2'h2:2'h2];
  assign T6800 = T6203[2'h3:2'h3];
  assign T6801 = T6830 ? T6816 : T6802;
  assign T6802 = T6815 ? T6809 : T6803;
  assign T6803 = T6808 ? T6806 : T6804;
  assign T6804 = T6805 ? counts_305 : counts_304;
  assign T6805 = T6203[1'h0:1'h0];
  assign T6806 = T6807 ? counts_307 : counts_306;
  assign T6807 = T6203[1'h0:1'h0];
  assign T6808 = T6203[1'h1:1'h1];
  assign T6809 = T6814 ? T6812 : T6810;
  assign T6810 = T6811 ? counts_309 : counts_308;
  assign T6811 = T6203[1'h0:1'h0];
  assign T6812 = T6813 ? counts_311 : counts_310;
  assign T6813 = T6203[1'h0:1'h0];
  assign T6814 = T6203[1'h1:1'h1];
  assign T6815 = T6203[2'h2:2'h2];
  assign T6816 = T6829 ? T6823 : T6817;
  assign T6817 = T6822 ? T6820 : T6818;
  assign T6818 = T6819 ? counts_313 : counts_312;
  assign T6819 = T6203[1'h0:1'h0];
  assign T6820 = T6821 ? counts_315 : counts_314;
  assign T6821 = T6203[1'h0:1'h0];
  assign T6822 = T6203[1'h1:1'h1];
  assign T6823 = T6828 ? T6826 : T6824;
  assign T6824 = T6825 ? counts_317 : counts_316;
  assign T6825 = T6203[1'h0:1'h0];
  assign T6826 = T6827 ? counts_319 : counts_318;
  assign T6827 = T6203[1'h0:1'h0];
  assign T6828 = T6203[1'h1:1'h1];
  assign T6829 = T6203[2'h2:2'h2];
  assign T6830 = T6203[2'h3:2'h3];
  assign T6831 = T6203[3'h4:3'h4];
  assign T6832 = T6203[3'h5:3'h5];
  assign T6833 = T6958 ? T6896 : T6834;
  assign T6834 = T6895 ? T6865 : T6835;
  assign T6835 = T6864 ? T6850 : T6836;
  assign T6836 = T6849 ? T6843 : T6837;
  assign T6837 = T6842 ? T6840 : T6838;
  assign T6838 = T6839 ? counts_321 : counts_320;
  assign T6839 = T6203[1'h0:1'h0];
  assign T6840 = T6841 ? counts_323 : counts_322;
  assign T6841 = T6203[1'h0:1'h0];
  assign T6842 = T6203[1'h1:1'h1];
  assign T6843 = T6848 ? T6846 : T6844;
  assign T6844 = T6845 ? counts_325 : counts_324;
  assign T6845 = T6203[1'h0:1'h0];
  assign T6846 = T6847 ? counts_327 : counts_326;
  assign T6847 = T6203[1'h0:1'h0];
  assign T6848 = T6203[1'h1:1'h1];
  assign T6849 = T6203[2'h2:2'h2];
  assign T6850 = T6863 ? T6857 : T6851;
  assign T6851 = T6856 ? T6854 : T6852;
  assign T6852 = T6853 ? counts_329 : counts_328;
  assign T6853 = T6203[1'h0:1'h0];
  assign T6854 = T6855 ? counts_331 : counts_330;
  assign T6855 = T6203[1'h0:1'h0];
  assign T6856 = T6203[1'h1:1'h1];
  assign T6857 = T6862 ? T6860 : T6858;
  assign T6858 = T6859 ? counts_333 : counts_332;
  assign T6859 = T6203[1'h0:1'h0];
  assign T6860 = T6861 ? counts_335 : counts_334;
  assign T6861 = T6203[1'h0:1'h0];
  assign T6862 = T6203[1'h1:1'h1];
  assign T6863 = T6203[2'h2:2'h2];
  assign T6864 = T6203[2'h3:2'h3];
  assign T6865 = T6894 ? T6880 : T6866;
  assign T6866 = T6879 ? T6873 : T6867;
  assign T6867 = T6872 ? T6870 : T6868;
  assign T6868 = T6869 ? counts_337 : counts_336;
  assign T6869 = T6203[1'h0:1'h0];
  assign T6870 = T6871 ? counts_339 : counts_338;
  assign T6871 = T6203[1'h0:1'h0];
  assign T6872 = T6203[1'h1:1'h1];
  assign T6873 = T6878 ? T6876 : T6874;
  assign T6874 = T6875 ? counts_341 : counts_340;
  assign T6875 = T6203[1'h0:1'h0];
  assign T6876 = T6877 ? counts_343 : counts_342;
  assign T6877 = T6203[1'h0:1'h0];
  assign T6878 = T6203[1'h1:1'h1];
  assign T6879 = T6203[2'h2:2'h2];
  assign T6880 = T6893 ? T6887 : T6881;
  assign T6881 = T6886 ? T6884 : T6882;
  assign T6882 = T6883 ? counts_345 : counts_344;
  assign T6883 = T6203[1'h0:1'h0];
  assign T6884 = T6885 ? counts_347 : counts_346;
  assign T6885 = T6203[1'h0:1'h0];
  assign T6886 = T6203[1'h1:1'h1];
  assign T6887 = T6892 ? T6890 : T6888;
  assign T6888 = T6889 ? counts_349 : counts_348;
  assign T6889 = T6203[1'h0:1'h0];
  assign T6890 = T6891 ? counts_351 : counts_350;
  assign T6891 = T6203[1'h0:1'h0];
  assign T6892 = T6203[1'h1:1'h1];
  assign T6893 = T6203[2'h2:2'h2];
  assign T6894 = T6203[2'h3:2'h3];
  assign T6895 = T6203[3'h4:3'h4];
  assign T6896 = T6957 ? T6927 : T6897;
  assign T6897 = T6926 ? T6912 : T6898;
  assign T6898 = T6911 ? T6905 : T6899;
  assign T6899 = T6904 ? T6902 : T6900;
  assign T6900 = T6901 ? counts_353 : counts_352;
  assign T6901 = T6203[1'h0:1'h0];
  assign T6902 = T6903 ? counts_355 : counts_354;
  assign T6903 = T6203[1'h0:1'h0];
  assign T6904 = T6203[1'h1:1'h1];
  assign T6905 = T6910 ? T6908 : T6906;
  assign T6906 = T6907 ? counts_357 : counts_356;
  assign T6907 = T6203[1'h0:1'h0];
  assign T6908 = T6909 ? counts_359 : counts_358;
  assign T6909 = T6203[1'h0:1'h0];
  assign T6910 = T6203[1'h1:1'h1];
  assign T6911 = T6203[2'h2:2'h2];
  assign T6912 = T6925 ? T6919 : T6913;
  assign T6913 = T6918 ? T6916 : T6914;
  assign T6914 = T6915 ? counts_361 : counts_360;
  assign T6915 = T6203[1'h0:1'h0];
  assign T6916 = T6917 ? counts_363 : counts_362;
  assign T6917 = T6203[1'h0:1'h0];
  assign T6918 = T6203[1'h1:1'h1];
  assign T6919 = T6924 ? T6922 : T6920;
  assign T6920 = T6921 ? counts_365 : counts_364;
  assign T6921 = T6203[1'h0:1'h0];
  assign T6922 = T6923 ? counts_367 : counts_366;
  assign T6923 = T6203[1'h0:1'h0];
  assign T6924 = T6203[1'h1:1'h1];
  assign T6925 = T6203[2'h2:2'h2];
  assign T6926 = T6203[2'h3:2'h3];
  assign T6927 = T6956 ? T6942 : T6928;
  assign T6928 = T6941 ? T6935 : T6929;
  assign T6929 = T6934 ? T6932 : T6930;
  assign T6930 = T6931 ? counts_369 : counts_368;
  assign T6931 = T6203[1'h0:1'h0];
  assign T6932 = T6933 ? counts_371 : counts_370;
  assign T6933 = T6203[1'h0:1'h0];
  assign T6934 = T6203[1'h1:1'h1];
  assign T6935 = T6940 ? T6938 : T6936;
  assign T6936 = T6937 ? counts_373 : counts_372;
  assign T6937 = T6203[1'h0:1'h0];
  assign T6938 = T6939 ? counts_375 : counts_374;
  assign T6939 = T6203[1'h0:1'h0];
  assign T6940 = T6203[1'h1:1'h1];
  assign T6941 = T6203[2'h2:2'h2];
  assign T6942 = T6955 ? T6949 : T6943;
  assign T6943 = T6948 ? T6946 : T6944;
  assign T6944 = T6945 ? counts_377 : counts_376;
  assign T6945 = T6203[1'h0:1'h0];
  assign T6946 = T6947 ? counts_379 : counts_378;
  assign T6947 = T6203[1'h0:1'h0];
  assign T6948 = T6203[1'h1:1'h1];
  assign T6949 = T6954 ? T6952 : T6950;
  assign T6950 = T6951 ? counts_381 : counts_380;
  assign T6951 = T6203[1'h0:1'h0];
  assign T6952 = T6953 ? counts_383 : counts_382;
  assign T6953 = T6203[1'h0:1'h0];
  assign T6954 = T6203[1'h1:1'h1];
  assign T6955 = T6203[2'h2:2'h2];
  assign T6956 = T6203[2'h3:2'h3];
  assign T6957 = T6203[3'h4:3'h4];
  assign T6958 = T6203[3'h5:3'h5];
  assign T6959 = T6203[3'h6:3'h6];
  assign T6960 = T7213 ? T7087 : T6961;
  assign T6961 = T7086 ? T7024 : T6962;
  assign T6962 = T7023 ? T6993 : T6963;
  assign T6963 = T6992 ? T6978 : T6964;
  assign T6964 = T6977 ? T6971 : T6965;
  assign T6965 = T6970 ? T6968 : T6966;
  assign T6966 = T6967 ? counts_385 : counts_384;
  assign T6967 = T6203[1'h0:1'h0];
  assign T6968 = T6969 ? counts_387 : counts_386;
  assign T6969 = T6203[1'h0:1'h0];
  assign T6970 = T6203[1'h1:1'h1];
  assign T6971 = T6976 ? T6974 : T6972;
  assign T6972 = T6973 ? counts_389 : counts_388;
  assign T6973 = T6203[1'h0:1'h0];
  assign T6974 = T6975 ? counts_391 : counts_390;
  assign T6975 = T6203[1'h0:1'h0];
  assign T6976 = T6203[1'h1:1'h1];
  assign T6977 = T6203[2'h2:2'h2];
  assign T6978 = T6991 ? T6985 : T6979;
  assign T6979 = T6984 ? T6982 : T6980;
  assign T6980 = T6981 ? counts_393 : counts_392;
  assign T6981 = T6203[1'h0:1'h0];
  assign T6982 = T6983 ? counts_395 : counts_394;
  assign T6983 = T6203[1'h0:1'h0];
  assign T6984 = T6203[1'h1:1'h1];
  assign T6985 = T6990 ? T6988 : T6986;
  assign T6986 = T6987 ? counts_397 : counts_396;
  assign T6987 = T6203[1'h0:1'h0];
  assign T6988 = T6989 ? counts_399 : counts_398;
  assign T6989 = T6203[1'h0:1'h0];
  assign T6990 = T6203[1'h1:1'h1];
  assign T6991 = T6203[2'h2:2'h2];
  assign T6992 = T6203[2'h3:2'h3];
  assign T6993 = T7022 ? T7008 : T6994;
  assign T6994 = T7007 ? T7001 : T6995;
  assign T6995 = T7000 ? T6998 : T6996;
  assign T6996 = T6997 ? counts_401 : counts_400;
  assign T6997 = T6203[1'h0:1'h0];
  assign T6998 = T6999 ? counts_403 : counts_402;
  assign T6999 = T6203[1'h0:1'h0];
  assign T7000 = T6203[1'h1:1'h1];
  assign T7001 = T7006 ? T7004 : T7002;
  assign T7002 = T7003 ? counts_405 : counts_404;
  assign T7003 = T6203[1'h0:1'h0];
  assign T7004 = T7005 ? counts_407 : counts_406;
  assign T7005 = T6203[1'h0:1'h0];
  assign T7006 = T6203[1'h1:1'h1];
  assign T7007 = T6203[2'h2:2'h2];
  assign T7008 = T7021 ? T7015 : T7009;
  assign T7009 = T7014 ? T7012 : T7010;
  assign T7010 = T7011 ? counts_409 : counts_408;
  assign T7011 = T6203[1'h0:1'h0];
  assign T7012 = T7013 ? counts_411 : counts_410;
  assign T7013 = T6203[1'h0:1'h0];
  assign T7014 = T6203[1'h1:1'h1];
  assign T7015 = T7020 ? T7018 : T7016;
  assign T7016 = T7017 ? counts_413 : counts_412;
  assign T7017 = T6203[1'h0:1'h0];
  assign T7018 = T7019 ? counts_415 : counts_414;
  assign T7019 = T6203[1'h0:1'h0];
  assign T7020 = T6203[1'h1:1'h1];
  assign T7021 = T6203[2'h2:2'h2];
  assign T7022 = T6203[2'h3:2'h3];
  assign T7023 = T6203[3'h4:3'h4];
  assign T7024 = T7085 ? T7055 : T7025;
  assign T7025 = T7054 ? T7040 : T7026;
  assign T7026 = T7039 ? T7033 : T7027;
  assign T7027 = T7032 ? T7030 : T7028;
  assign T7028 = T7029 ? counts_417 : counts_416;
  assign T7029 = T6203[1'h0:1'h0];
  assign T7030 = T7031 ? counts_419 : counts_418;
  assign T7031 = T6203[1'h0:1'h0];
  assign T7032 = T6203[1'h1:1'h1];
  assign T7033 = T7038 ? T7036 : T7034;
  assign T7034 = T7035 ? counts_421 : counts_420;
  assign T7035 = T6203[1'h0:1'h0];
  assign T7036 = T7037 ? counts_423 : counts_422;
  assign T7037 = T6203[1'h0:1'h0];
  assign T7038 = T6203[1'h1:1'h1];
  assign T7039 = T6203[2'h2:2'h2];
  assign T7040 = T7053 ? T7047 : T7041;
  assign T7041 = T7046 ? T7044 : T7042;
  assign T7042 = T7043 ? counts_425 : counts_424;
  assign T7043 = T6203[1'h0:1'h0];
  assign T7044 = T7045 ? counts_427 : counts_426;
  assign T7045 = T6203[1'h0:1'h0];
  assign T7046 = T6203[1'h1:1'h1];
  assign T7047 = T7052 ? T7050 : T7048;
  assign T7048 = T7049 ? counts_429 : counts_428;
  assign T7049 = T6203[1'h0:1'h0];
  assign T7050 = T7051 ? counts_431 : counts_430;
  assign T7051 = T6203[1'h0:1'h0];
  assign T7052 = T6203[1'h1:1'h1];
  assign T7053 = T6203[2'h2:2'h2];
  assign T7054 = T6203[2'h3:2'h3];
  assign T7055 = T7084 ? T7070 : T7056;
  assign T7056 = T7069 ? T7063 : T7057;
  assign T7057 = T7062 ? T7060 : T7058;
  assign T7058 = T7059 ? counts_433 : counts_432;
  assign T7059 = T6203[1'h0:1'h0];
  assign T7060 = T7061 ? counts_435 : counts_434;
  assign T7061 = T6203[1'h0:1'h0];
  assign T7062 = T6203[1'h1:1'h1];
  assign T7063 = T7068 ? T7066 : T7064;
  assign T7064 = T7065 ? counts_437 : counts_436;
  assign T7065 = T6203[1'h0:1'h0];
  assign T7066 = T7067 ? counts_439 : counts_438;
  assign T7067 = T6203[1'h0:1'h0];
  assign T7068 = T6203[1'h1:1'h1];
  assign T7069 = T6203[2'h2:2'h2];
  assign T7070 = T7083 ? T7077 : T7071;
  assign T7071 = T7076 ? T7074 : T7072;
  assign T7072 = T7073 ? counts_441 : counts_440;
  assign T7073 = T6203[1'h0:1'h0];
  assign T7074 = T7075 ? counts_443 : counts_442;
  assign T7075 = T6203[1'h0:1'h0];
  assign T7076 = T6203[1'h1:1'h1];
  assign T7077 = T7082 ? T7080 : T7078;
  assign T7078 = T7079 ? counts_445 : counts_444;
  assign T7079 = T6203[1'h0:1'h0];
  assign T7080 = T7081 ? counts_447 : counts_446;
  assign T7081 = T6203[1'h0:1'h0];
  assign T7082 = T6203[1'h1:1'h1];
  assign T7083 = T6203[2'h2:2'h2];
  assign T7084 = T6203[2'h3:2'h3];
  assign T7085 = T6203[3'h4:3'h4];
  assign T7086 = T6203[3'h5:3'h5];
  assign T7087 = T7212 ? T7150 : T7088;
  assign T7088 = T7149 ? T7119 : T7089;
  assign T7089 = T7118 ? T7104 : T7090;
  assign T7090 = T7103 ? T7097 : T7091;
  assign T7091 = T7096 ? T7094 : T7092;
  assign T7092 = T7093 ? counts_449 : counts_448;
  assign T7093 = T6203[1'h0:1'h0];
  assign T7094 = T7095 ? counts_451 : counts_450;
  assign T7095 = T6203[1'h0:1'h0];
  assign T7096 = T6203[1'h1:1'h1];
  assign T7097 = T7102 ? T7100 : T7098;
  assign T7098 = T7099 ? counts_453 : counts_452;
  assign T7099 = T6203[1'h0:1'h0];
  assign T7100 = T7101 ? counts_455 : counts_454;
  assign T7101 = T6203[1'h0:1'h0];
  assign T7102 = T6203[1'h1:1'h1];
  assign T7103 = T6203[2'h2:2'h2];
  assign T7104 = T7117 ? T7111 : T7105;
  assign T7105 = T7110 ? T7108 : T7106;
  assign T7106 = T7107 ? counts_457 : counts_456;
  assign T7107 = T6203[1'h0:1'h0];
  assign T7108 = T7109 ? counts_459 : counts_458;
  assign T7109 = T6203[1'h0:1'h0];
  assign T7110 = T6203[1'h1:1'h1];
  assign T7111 = T7116 ? T7114 : T7112;
  assign T7112 = T7113 ? counts_461 : counts_460;
  assign T7113 = T6203[1'h0:1'h0];
  assign T7114 = T7115 ? counts_463 : counts_462;
  assign T7115 = T6203[1'h0:1'h0];
  assign T7116 = T6203[1'h1:1'h1];
  assign T7117 = T6203[2'h2:2'h2];
  assign T7118 = T6203[2'h3:2'h3];
  assign T7119 = T7148 ? T7134 : T7120;
  assign T7120 = T7133 ? T7127 : T7121;
  assign T7121 = T7126 ? T7124 : T7122;
  assign T7122 = T7123 ? counts_465 : counts_464;
  assign T7123 = T6203[1'h0:1'h0];
  assign T7124 = T7125 ? counts_467 : counts_466;
  assign T7125 = T6203[1'h0:1'h0];
  assign T7126 = T6203[1'h1:1'h1];
  assign T7127 = T7132 ? T7130 : T7128;
  assign T7128 = T7129 ? counts_469 : counts_468;
  assign T7129 = T6203[1'h0:1'h0];
  assign T7130 = T7131 ? counts_471 : counts_470;
  assign T7131 = T6203[1'h0:1'h0];
  assign T7132 = T6203[1'h1:1'h1];
  assign T7133 = T6203[2'h2:2'h2];
  assign T7134 = T7147 ? T7141 : T7135;
  assign T7135 = T7140 ? T7138 : T7136;
  assign T7136 = T7137 ? counts_473 : counts_472;
  assign T7137 = T6203[1'h0:1'h0];
  assign T7138 = T7139 ? counts_475 : counts_474;
  assign T7139 = T6203[1'h0:1'h0];
  assign T7140 = T6203[1'h1:1'h1];
  assign T7141 = T7146 ? T7144 : T7142;
  assign T7142 = T7143 ? counts_477 : counts_476;
  assign T7143 = T6203[1'h0:1'h0];
  assign T7144 = T7145 ? counts_479 : counts_478;
  assign T7145 = T6203[1'h0:1'h0];
  assign T7146 = T6203[1'h1:1'h1];
  assign T7147 = T6203[2'h2:2'h2];
  assign T7148 = T6203[2'h3:2'h3];
  assign T7149 = T6203[3'h4:3'h4];
  assign T7150 = T7211 ? T7181 : T7151;
  assign T7151 = T7180 ? T7166 : T7152;
  assign T7152 = T7165 ? T7159 : T7153;
  assign T7153 = T7158 ? T7156 : T7154;
  assign T7154 = T7155 ? counts_481 : counts_480;
  assign T7155 = T6203[1'h0:1'h0];
  assign T7156 = T7157 ? counts_483 : counts_482;
  assign T7157 = T6203[1'h0:1'h0];
  assign T7158 = T6203[1'h1:1'h1];
  assign T7159 = T7164 ? T7162 : T7160;
  assign T7160 = T7161 ? counts_485 : counts_484;
  assign T7161 = T6203[1'h0:1'h0];
  assign T7162 = T7163 ? counts_487 : counts_486;
  assign T7163 = T6203[1'h0:1'h0];
  assign T7164 = T6203[1'h1:1'h1];
  assign T7165 = T6203[2'h2:2'h2];
  assign T7166 = T7179 ? T7173 : T7167;
  assign T7167 = T7172 ? T7170 : T7168;
  assign T7168 = T7169 ? counts_489 : counts_488;
  assign T7169 = T6203[1'h0:1'h0];
  assign T7170 = T7171 ? counts_491 : counts_490;
  assign T7171 = T6203[1'h0:1'h0];
  assign T7172 = T6203[1'h1:1'h1];
  assign T7173 = T7178 ? T7176 : T7174;
  assign T7174 = T7175 ? counts_493 : counts_492;
  assign T7175 = T6203[1'h0:1'h0];
  assign T7176 = T7177 ? counts_495 : counts_494;
  assign T7177 = T6203[1'h0:1'h0];
  assign T7178 = T6203[1'h1:1'h1];
  assign T7179 = T6203[2'h2:2'h2];
  assign T7180 = T6203[2'h3:2'h3];
  assign T7181 = T7210 ? T7196 : T7182;
  assign T7182 = T7195 ? T7189 : T7183;
  assign T7183 = T7188 ? T7186 : T7184;
  assign T7184 = T7185 ? counts_497 : counts_496;
  assign T7185 = T6203[1'h0:1'h0];
  assign T7186 = T7187 ? counts_499 : counts_498;
  assign T7187 = T6203[1'h0:1'h0];
  assign T7188 = T6203[1'h1:1'h1];
  assign T7189 = T7194 ? T7192 : T7190;
  assign T7190 = T7191 ? counts_501 : counts_500;
  assign T7191 = T6203[1'h0:1'h0];
  assign T7192 = T7193 ? counts_503 : counts_502;
  assign T7193 = T6203[1'h0:1'h0];
  assign T7194 = T6203[1'h1:1'h1];
  assign T7195 = T6203[2'h2:2'h2];
  assign T7196 = T7209 ? T7203 : T7197;
  assign T7197 = T7202 ? T7200 : T7198;
  assign T7198 = T7199 ? counts_505 : counts_504;
  assign T7199 = T6203[1'h0:1'h0];
  assign T7200 = T7201 ? counts_507 : counts_506;
  assign T7201 = T6203[1'h0:1'h0];
  assign T7202 = T6203[1'h1:1'h1];
  assign T7203 = T7208 ? T7206 : T7204;
  assign T7204 = T7205 ? counts_509 : counts_508;
  assign T7205 = T6203[1'h0:1'h0];
  assign T7206 = T7207 ? counts_511 : counts_510;
  assign T7207 = T6203[1'h0:1'h0];
  assign T7208 = T6203[1'h1:1'h1];
  assign T7209 = T6203[2'h2:2'h2];
  assign T7210 = T6203[2'h3:2'h3];
  assign T7211 = T6203[3'h4:3'h4];
  assign T7212 = T6203[3'h5:3'h5];
  assign T7213 = T6203[3'h6:3'h6];
  assign T7214 = T6203[3'h7:3'h7];
  assign T7215 = T6203[4'h8:4'h8];
  assign T7216 = T8237 ? T7727 : T7217;
  assign T7217 = T7726 ? T7472 : T7218;
  assign T7218 = T7471 ? T7345 : T7219;
  assign T7219 = T7344 ? T7282 : T7220;
  assign T7220 = T7281 ? T7251 : T7221;
  assign T7221 = T7250 ? T7236 : T7222;
  assign T7222 = T7235 ? T7229 : T7223;
  assign T7223 = T7228 ? T7226 : T7224;
  assign T7224 = T7225 ? counts_513 : counts_512;
  assign T7225 = T6203[1'h0:1'h0];
  assign T7226 = T7227 ? counts_515 : counts_514;
  assign T7227 = T6203[1'h0:1'h0];
  assign T7228 = T6203[1'h1:1'h1];
  assign T7229 = T7234 ? T7232 : T7230;
  assign T7230 = T7231 ? counts_517 : counts_516;
  assign T7231 = T6203[1'h0:1'h0];
  assign T7232 = T7233 ? counts_519 : counts_518;
  assign T7233 = T6203[1'h0:1'h0];
  assign T7234 = T6203[1'h1:1'h1];
  assign T7235 = T6203[2'h2:2'h2];
  assign T7236 = T7249 ? T7243 : T7237;
  assign T7237 = T7242 ? T7240 : T7238;
  assign T7238 = T7239 ? counts_521 : counts_520;
  assign T7239 = T6203[1'h0:1'h0];
  assign T7240 = T7241 ? counts_523 : counts_522;
  assign T7241 = T6203[1'h0:1'h0];
  assign T7242 = T6203[1'h1:1'h1];
  assign T7243 = T7248 ? T7246 : T7244;
  assign T7244 = T7245 ? counts_525 : counts_524;
  assign T7245 = T6203[1'h0:1'h0];
  assign T7246 = T7247 ? counts_527 : counts_526;
  assign T7247 = T6203[1'h0:1'h0];
  assign T7248 = T6203[1'h1:1'h1];
  assign T7249 = T6203[2'h2:2'h2];
  assign T7250 = T6203[2'h3:2'h3];
  assign T7251 = T7280 ? T7266 : T7252;
  assign T7252 = T7265 ? T7259 : T7253;
  assign T7253 = T7258 ? T7256 : T7254;
  assign T7254 = T7255 ? counts_529 : counts_528;
  assign T7255 = T6203[1'h0:1'h0];
  assign T7256 = T7257 ? counts_531 : counts_530;
  assign T7257 = T6203[1'h0:1'h0];
  assign T7258 = T6203[1'h1:1'h1];
  assign T7259 = T7264 ? T7262 : T7260;
  assign T7260 = T7261 ? counts_533 : counts_532;
  assign T7261 = T6203[1'h0:1'h0];
  assign T7262 = T7263 ? counts_535 : counts_534;
  assign T7263 = T6203[1'h0:1'h0];
  assign T7264 = T6203[1'h1:1'h1];
  assign T7265 = T6203[2'h2:2'h2];
  assign T7266 = T7279 ? T7273 : T7267;
  assign T7267 = T7272 ? T7270 : T7268;
  assign T7268 = T7269 ? counts_537 : counts_536;
  assign T7269 = T6203[1'h0:1'h0];
  assign T7270 = T7271 ? counts_539 : counts_538;
  assign T7271 = T6203[1'h0:1'h0];
  assign T7272 = T6203[1'h1:1'h1];
  assign T7273 = T7278 ? T7276 : T7274;
  assign T7274 = T7275 ? counts_541 : counts_540;
  assign T7275 = T6203[1'h0:1'h0];
  assign T7276 = T7277 ? counts_543 : counts_542;
  assign T7277 = T6203[1'h0:1'h0];
  assign T7278 = T6203[1'h1:1'h1];
  assign T7279 = T6203[2'h2:2'h2];
  assign T7280 = T6203[2'h3:2'h3];
  assign T7281 = T6203[3'h4:3'h4];
  assign T7282 = T7343 ? T7313 : T7283;
  assign T7283 = T7312 ? T7298 : T7284;
  assign T7284 = T7297 ? T7291 : T7285;
  assign T7285 = T7290 ? T7288 : T7286;
  assign T7286 = T7287 ? counts_545 : counts_544;
  assign T7287 = T6203[1'h0:1'h0];
  assign T7288 = T7289 ? counts_547 : counts_546;
  assign T7289 = T6203[1'h0:1'h0];
  assign T7290 = T6203[1'h1:1'h1];
  assign T7291 = T7296 ? T7294 : T7292;
  assign T7292 = T7293 ? counts_549 : counts_548;
  assign T7293 = T6203[1'h0:1'h0];
  assign T7294 = T7295 ? counts_551 : counts_550;
  assign T7295 = T6203[1'h0:1'h0];
  assign T7296 = T6203[1'h1:1'h1];
  assign T7297 = T6203[2'h2:2'h2];
  assign T7298 = T7311 ? T7305 : T7299;
  assign T7299 = T7304 ? T7302 : T7300;
  assign T7300 = T7301 ? counts_553 : counts_552;
  assign T7301 = T6203[1'h0:1'h0];
  assign T7302 = T7303 ? counts_555 : counts_554;
  assign T7303 = T6203[1'h0:1'h0];
  assign T7304 = T6203[1'h1:1'h1];
  assign T7305 = T7310 ? T7308 : T7306;
  assign T7306 = T7307 ? counts_557 : counts_556;
  assign T7307 = T6203[1'h0:1'h0];
  assign T7308 = T7309 ? counts_559 : counts_558;
  assign T7309 = T6203[1'h0:1'h0];
  assign T7310 = T6203[1'h1:1'h1];
  assign T7311 = T6203[2'h2:2'h2];
  assign T7312 = T6203[2'h3:2'h3];
  assign T7313 = T7342 ? T7328 : T7314;
  assign T7314 = T7327 ? T7321 : T7315;
  assign T7315 = T7320 ? T7318 : T7316;
  assign T7316 = T7317 ? counts_561 : counts_560;
  assign T7317 = T6203[1'h0:1'h0];
  assign T7318 = T7319 ? counts_563 : counts_562;
  assign T7319 = T6203[1'h0:1'h0];
  assign T7320 = T6203[1'h1:1'h1];
  assign T7321 = T7326 ? T7324 : T7322;
  assign T7322 = T7323 ? counts_565 : counts_564;
  assign T7323 = T6203[1'h0:1'h0];
  assign T7324 = T7325 ? counts_567 : counts_566;
  assign T7325 = T6203[1'h0:1'h0];
  assign T7326 = T6203[1'h1:1'h1];
  assign T7327 = T6203[2'h2:2'h2];
  assign T7328 = T7341 ? T7335 : T7329;
  assign T7329 = T7334 ? T7332 : T7330;
  assign T7330 = T7331 ? counts_569 : counts_568;
  assign T7331 = T6203[1'h0:1'h0];
  assign T7332 = T7333 ? counts_571 : counts_570;
  assign T7333 = T6203[1'h0:1'h0];
  assign T7334 = T6203[1'h1:1'h1];
  assign T7335 = T7340 ? T7338 : T7336;
  assign T7336 = T7337 ? counts_573 : counts_572;
  assign T7337 = T6203[1'h0:1'h0];
  assign T7338 = T7339 ? counts_575 : counts_574;
  assign T7339 = T6203[1'h0:1'h0];
  assign T7340 = T6203[1'h1:1'h1];
  assign T7341 = T6203[2'h2:2'h2];
  assign T7342 = T6203[2'h3:2'h3];
  assign T7343 = T6203[3'h4:3'h4];
  assign T7344 = T6203[3'h5:3'h5];
  assign T7345 = T7470 ? T7408 : T7346;
  assign T7346 = T7407 ? T7377 : T7347;
  assign T7347 = T7376 ? T7362 : T7348;
  assign T7348 = T7361 ? T7355 : T7349;
  assign T7349 = T7354 ? T7352 : T7350;
  assign T7350 = T7351 ? counts_577 : counts_576;
  assign T7351 = T6203[1'h0:1'h0];
  assign T7352 = T7353 ? counts_579 : counts_578;
  assign T7353 = T6203[1'h0:1'h0];
  assign T7354 = T6203[1'h1:1'h1];
  assign T7355 = T7360 ? T7358 : T7356;
  assign T7356 = T7357 ? counts_581 : counts_580;
  assign T7357 = T6203[1'h0:1'h0];
  assign T7358 = T7359 ? counts_583 : counts_582;
  assign T7359 = T6203[1'h0:1'h0];
  assign T7360 = T6203[1'h1:1'h1];
  assign T7361 = T6203[2'h2:2'h2];
  assign T7362 = T7375 ? T7369 : T7363;
  assign T7363 = T7368 ? T7366 : T7364;
  assign T7364 = T7365 ? counts_585 : counts_584;
  assign T7365 = T6203[1'h0:1'h0];
  assign T7366 = T7367 ? counts_587 : counts_586;
  assign T7367 = T6203[1'h0:1'h0];
  assign T7368 = T6203[1'h1:1'h1];
  assign T7369 = T7374 ? T7372 : T7370;
  assign T7370 = T7371 ? counts_589 : counts_588;
  assign T7371 = T6203[1'h0:1'h0];
  assign T7372 = T7373 ? counts_591 : counts_590;
  assign T7373 = T6203[1'h0:1'h0];
  assign T7374 = T6203[1'h1:1'h1];
  assign T7375 = T6203[2'h2:2'h2];
  assign T7376 = T6203[2'h3:2'h3];
  assign T7377 = T7406 ? T7392 : T7378;
  assign T7378 = T7391 ? T7385 : T7379;
  assign T7379 = T7384 ? T7382 : T7380;
  assign T7380 = T7381 ? counts_593 : counts_592;
  assign T7381 = T6203[1'h0:1'h0];
  assign T7382 = T7383 ? counts_595 : counts_594;
  assign T7383 = T6203[1'h0:1'h0];
  assign T7384 = T6203[1'h1:1'h1];
  assign T7385 = T7390 ? T7388 : T7386;
  assign T7386 = T7387 ? counts_597 : counts_596;
  assign T7387 = T6203[1'h0:1'h0];
  assign T7388 = T7389 ? counts_599 : counts_598;
  assign T7389 = T6203[1'h0:1'h0];
  assign T7390 = T6203[1'h1:1'h1];
  assign T7391 = T6203[2'h2:2'h2];
  assign T7392 = T7405 ? T7399 : T7393;
  assign T7393 = T7398 ? T7396 : T7394;
  assign T7394 = T7395 ? counts_601 : counts_600;
  assign T7395 = T6203[1'h0:1'h0];
  assign T7396 = T7397 ? counts_603 : counts_602;
  assign T7397 = T6203[1'h0:1'h0];
  assign T7398 = T6203[1'h1:1'h1];
  assign T7399 = T7404 ? T7402 : T7400;
  assign T7400 = T7401 ? counts_605 : counts_604;
  assign T7401 = T6203[1'h0:1'h0];
  assign T7402 = T7403 ? counts_607 : counts_606;
  assign T7403 = T6203[1'h0:1'h0];
  assign T7404 = T6203[1'h1:1'h1];
  assign T7405 = T6203[2'h2:2'h2];
  assign T7406 = T6203[2'h3:2'h3];
  assign T7407 = T6203[3'h4:3'h4];
  assign T7408 = T7469 ? T7439 : T7409;
  assign T7409 = T7438 ? T7424 : T7410;
  assign T7410 = T7423 ? T7417 : T7411;
  assign T7411 = T7416 ? T7414 : T7412;
  assign T7412 = T7413 ? counts_609 : counts_608;
  assign T7413 = T6203[1'h0:1'h0];
  assign T7414 = T7415 ? counts_611 : counts_610;
  assign T7415 = T6203[1'h0:1'h0];
  assign T7416 = T6203[1'h1:1'h1];
  assign T7417 = T7422 ? T7420 : T7418;
  assign T7418 = T7419 ? counts_613 : counts_612;
  assign T7419 = T6203[1'h0:1'h0];
  assign T7420 = T7421 ? counts_615 : counts_614;
  assign T7421 = T6203[1'h0:1'h0];
  assign T7422 = T6203[1'h1:1'h1];
  assign T7423 = T6203[2'h2:2'h2];
  assign T7424 = T7437 ? T7431 : T7425;
  assign T7425 = T7430 ? T7428 : T7426;
  assign T7426 = T7427 ? counts_617 : counts_616;
  assign T7427 = T6203[1'h0:1'h0];
  assign T7428 = T7429 ? counts_619 : counts_618;
  assign T7429 = T6203[1'h0:1'h0];
  assign T7430 = T6203[1'h1:1'h1];
  assign T7431 = T7436 ? T7434 : T7432;
  assign T7432 = T7433 ? counts_621 : counts_620;
  assign T7433 = T6203[1'h0:1'h0];
  assign T7434 = T7435 ? counts_623 : counts_622;
  assign T7435 = T6203[1'h0:1'h0];
  assign T7436 = T6203[1'h1:1'h1];
  assign T7437 = T6203[2'h2:2'h2];
  assign T7438 = T6203[2'h3:2'h3];
  assign T7439 = T7468 ? T7454 : T7440;
  assign T7440 = T7453 ? T7447 : T7441;
  assign T7441 = T7446 ? T7444 : T7442;
  assign T7442 = T7443 ? counts_625 : counts_624;
  assign T7443 = T6203[1'h0:1'h0];
  assign T7444 = T7445 ? counts_627 : counts_626;
  assign T7445 = T6203[1'h0:1'h0];
  assign T7446 = T6203[1'h1:1'h1];
  assign T7447 = T7452 ? T7450 : T7448;
  assign T7448 = T7449 ? counts_629 : counts_628;
  assign T7449 = T6203[1'h0:1'h0];
  assign T7450 = T7451 ? counts_631 : counts_630;
  assign T7451 = T6203[1'h0:1'h0];
  assign T7452 = T6203[1'h1:1'h1];
  assign T7453 = T6203[2'h2:2'h2];
  assign T7454 = T7467 ? T7461 : T7455;
  assign T7455 = T7460 ? T7458 : T7456;
  assign T7456 = T7457 ? counts_633 : counts_632;
  assign T7457 = T6203[1'h0:1'h0];
  assign T7458 = T7459 ? counts_635 : counts_634;
  assign T7459 = T6203[1'h0:1'h0];
  assign T7460 = T6203[1'h1:1'h1];
  assign T7461 = T7466 ? T7464 : T7462;
  assign T7462 = T7463 ? counts_637 : counts_636;
  assign T7463 = T6203[1'h0:1'h0];
  assign T7464 = T7465 ? counts_639 : counts_638;
  assign T7465 = T6203[1'h0:1'h0];
  assign T7466 = T6203[1'h1:1'h1];
  assign T7467 = T6203[2'h2:2'h2];
  assign T7468 = T6203[2'h3:2'h3];
  assign T7469 = T6203[3'h4:3'h4];
  assign T7470 = T6203[3'h5:3'h5];
  assign T7471 = T6203[3'h6:3'h6];
  assign T7472 = T7725 ? T7599 : T7473;
  assign T7473 = T7598 ? T7536 : T7474;
  assign T7474 = T7535 ? T7505 : T7475;
  assign T7475 = T7504 ? T7490 : T7476;
  assign T7476 = T7489 ? T7483 : T7477;
  assign T7477 = T7482 ? T7480 : T7478;
  assign T7478 = T7479 ? counts_641 : counts_640;
  assign T7479 = T6203[1'h0:1'h0];
  assign T7480 = T7481 ? counts_643 : counts_642;
  assign T7481 = T6203[1'h0:1'h0];
  assign T7482 = T6203[1'h1:1'h1];
  assign T7483 = T7488 ? T7486 : T7484;
  assign T7484 = T7485 ? counts_645 : counts_644;
  assign T7485 = T6203[1'h0:1'h0];
  assign T7486 = T7487 ? counts_647 : counts_646;
  assign T7487 = T6203[1'h0:1'h0];
  assign T7488 = T6203[1'h1:1'h1];
  assign T7489 = T6203[2'h2:2'h2];
  assign T7490 = T7503 ? T7497 : T7491;
  assign T7491 = T7496 ? T7494 : T7492;
  assign T7492 = T7493 ? counts_649 : counts_648;
  assign T7493 = T6203[1'h0:1'h0];
  assign T7494 = T7495 ? counts_651 : counts_650;
  assign T7495 = T6203[1'h0:1'h0];
  assign T7496 = T6203[1'h1:1'h1];
  assign T7497 = T7502 ? T7500 : T7498;
  assign T7498 = T7499 ? counts_653 : counts_652;
  assign T7499 = T6203[1'h0:1'h0];
  assign T7500 = T7501 ? counts_655 : counts_654;
  assign T7501 = T6203[1'h0:1'h0];
  assign T7502 = T6203[1'h1:1'h1];
  assign T7503 = T6203[2'h2:2'h2];
  assign T7504 = T6203[2'h3:2'h3];
  assign T7505 = T7534 ? T7520 : T7506;
  assign T7506 = T7519 ? T7513 : T7507;
  assign T7507 = T7512 ? T7510 : T7508;
  assign T7508 = T7509 ? counts_657 : counts_656;
  assign T7509 = T6203[1'h0:1'h0];
  assign T7510 = T7511 ? counts_659 : counts_658;
  assign T7511 = T6203[1'h0:1'h0];
  assign T7512 = T6203[1'h1:1'h1];
  assign T7513 = T7518 ? T7516 : T7514;
  assign T7514 = T7515 ? counts_661 : counts_660;
  assign T7515 = T6203[1'h0:1'h0];
  assign T7516 = T7517 ? counts_663 : counts_662;
  assign T7517 = T6203[1'h0:1'h0];
  assign T7518 = T6203[1'h1:1'h1];
  assign T7519 = T6203[2'h2:2'h2];
  assign T7520 = T7533 ? T7527 : T7521;
  assign T7521 = T7526 ? T7524 : T7522;
  assign T7522 = T7523 ? counts_665 : counts_664;
  assign T7523 = T6203[1'h0:1'h0];
  assign T7524 = T7525 ? counts_667 : counts_666;
  assign T7525 = T6203[1'h0:1'h0];
  assign T7526 = T6203[1'h1:1'h1];
  assign T7527 = T7532 ? T7530 : T7528;
  assign T7528 = T7529 ? counts_669 : counts_668;
  assign T7529 = T6203[1'h0:1'h0];
  assign T7530 = T7531 ? counts_671 : counts_670;
  assign T7531 = T6203[1'h0:1'h0];
  assign T7532 = T6203[1'h1:1'h1];
  assign T7533 = T6203[2'h2:2'h2];
  assign T7534 = T6203[2'h3:2'h3];
  assign T7535 = T6203[3'h4:3'h4];
  assign T7536 = T7597 ? T7567 : T7537;
  assign T7537 = T7566 ? T7552 : T7538;
  assign T7538 = T7551 ? T7545 : T7539;
  assign T7539 = T7544 ? T7542 : T7540;
  assign T7540 = T7541 ? counts_673 : counts_672;
  assign T7541 = T6203[1'h0:1'h0];
  assign T7542 = T7543 ? counts_675 : counts_674;
  assign T7543 = T6203[1'h0:1'h0];
  assign T7544 = T6203[1'h1:1'h1];
  assign T7545 = T7550 ? T7548 : T7546;
  assign T7546 = T7547 ? counts_677 : counts_676;
  assign T7547 = T6203[1'h0:1'h0];
  assign T7548 = T7549 ? counts_679 : counts_678;
  assign T7549 = T6203[1'h0:1'h0];
  assign T7550 = T6203[1'h1:1'h1];
  assign T7551 = T6203[2'h2:2'h2];
  assign T7552 = T7565 ? T7559 : T7553;
  assign T7553 = T7558 ? T7556 : T7554;
  assign T7554 = T7555 ? counts_681 : counts_680;
  assign T7555 = T6203[1'h0:1'h0];
  assign T7556 = T7557 ? counts_683 : counts_682;
  assign T7557 = T6203[1'h0:1'h0];
  assign T7558 = T6203[1'h1:1'h1];
  assign T7559 = T7564 ? T7562 : T7560;
  assign T7560 = T7561 ? counts_685 : counts_684;
  assign T7561 = T6203[1'h0:1'h0];
  assign T7562 = T7563 ? counts_687 : counts_686;
  assign T7563 = T6203[1'h0:1'h0];
  assign T7564 = T6203[1'h1:1'h1];
  assign T7565 = T6203[2'h2:2'h2];
  assign T7566 = T6203[2'h3:2'h3];
  assign T7567 = T7596 ? T7582 : T7568;
  assign T7568 = T7581 ? T7575 : T7569;
  assign T7569 = T7574 ? T7572 : T7570;
  assign T7570 = T7571 ? counts_689 : counts_688;
  assign T7571 = T6203[1'h0:1'h0];
  assign T7572 = T7573 ? counts_691 : counts_690;
  assign T7573 = T6203[1'h0:1'h0];
  assign T7574 = T6203[1'h1:1'h1];
  assign T7575 = T7580 ? T7578 : T7576;
  assign T7576 = T7577 ? counts_693 : counts_692;
  assign T7577 = T6203[1'h0:1'h0];
  assign T7578 = T7579 ? counts_695 : counts_694;
  assign T7579 = T6203[1'h0:1'h0];
  assign T7580 = T6203[1'h1:1'h1];
  assign T7581 = T6203[2'h2:2'h2];
  assign T7582 = T7595 ? T7589 : T7583;
  assign T7583 = T7588 ? T7586 : T7584;
  assign T7584 = T7585 ? counts_697 : counts_696;
  assign T7585 = T6203[1'h0:1'h0];
  assign T7586 = T7587 ? counts_699 : counts_698;
  assign T7587 = T6203[1'h0:1'h0];
  assign T7588 = T6203[1'h1:1'h1];
  assign T7589 = T7594 ? T7592 : T7590;
  assign T7590 = T7591 ? counts_701 : counts_700;
  assign T7591 = T6203[1'h0:1'h0];
  assign T7592 = T7593 ? counts_703 : counts_702;
  assign T7593 = T6203[1'h0:1'h0];
  assign T7594 = T6203[1'h1:1'h1];
  assign T7595 = T6203[2'h2:2'h2];
  assign T7596 = T6203[2'h3:2'h3];
  assign T7597 = T6203[3'h4:3'h4];
  assign T7598 = T6203[3'h5:3'h5];
  assign T7599 = T7724 ? T7662 : T7600;
  assign T7600 = T7661 ? T7631 : T7601;
  assign T7601 = T7630 ? T7616 : T7602;
  assign T7602 = T7615 ? T7609 : T7603;
  assign T7603 = T7608 ? T7606 : T7604;
  assign T7604 = T7605 ? counts_705 : counts_704;
  assign T7605 = T6203[1'h0:1'h0];
  assign T7606 = T7607 ? counts_707 : counts_706;
  assign T7607 = T6203[1'h0:1'h0];
  assign T7608 = T6203[1'h1:1'h1];
  assign T7609 = T7614 ? T7612 : T7610;
  assign T7610 = T7611 ? counts_709 : counts_708;
  assign T7611 = T6203[1'h0:1'h0];
  assign T7612 = T7613 ? counts_711 : counts_710;
  assign T7613 = T6203[1'h0:1'h0];
  assign T7614 = T6203[1'h1:1'h1];
  assign T7615 = T6203[2'h2:2'h2];
  assign T7616 = T7629 ? T7623 : T7617;
  assign T7617 = T7622 ? T7620 : T7618;
  assign T7618 = T7619 ? counts_713 : counts_712;
  assign T7619 = T6203[1'h0:1'h0];
  assign T7620 = T7621 ? counts_715 : counts_714;
  assign T7621 = T6203[1'h0:1'h0];
  assign T7622 = T6203[1'h1:1'h1];
  assign T7623 = T7628 ? T7626 : T7624;
  assign T7624 = T7625 ? counts_717 : counts_716;
  assign T7625 = T6203[1'h0:1'h0];
  assign T7626 = T7627 ? counts_719 : counts_718;
  assign T7627 = T6203[1'h0:1'h0];
  assign T7628 = T6203[1'h1:1'h1];
  assign T7629 = T6203[2'h2:2'h2];
  assign T7630 = T6203[2'h3:2'h3];
  assign T7631 = T7660 ? T7646 : T7632;
  assign T7632 = T7645 ? T7639 : T7633;
  assign T7633 = T7638 ? T7636 : T7634;
  assign T7634 = T7635 ? counts_721 : counts_720;
  assign T7635 = T6203[1'h0:1'h0];
  assign T7636 = T7637 ? counts_723 : counts_722;
  assign T7637 = T6203[1'h0:1'h0];
  assign T7638 = T6203[1'h1:1'h1];
  assign T7639 = T7644 ? T7642 : T7640;
  assign T7640 = T7641 ? counts_725 : counts_724;
  assign T7641 = T6203[1'h0:1'h0];
  assign T7642 = T7643 ? counts_727 : counts_726;
  assign T7643 = T6203[1'h0:1'h0];
  assign T7644 = T6203[1'h1:1'h1];
  assign T7645 = T6203[2'h2:2'h2];
  assign T7646 = T7659 ? T7653 : T7647;
  assign T7647 = T7652 ? T7650 : T7648;
  assign T7648 = T7649 ? counts_729 : counts_728;
  assign T7649 = T6203[1'h0:1'h0];
  assign T7650 = T7651 ? counts_731 : counts_730;
  assign T7651 = T6203[1'h0:1'h0];
  assign T7652 = T6203[1'h1:1'h1];
  assign T7653 = T7658 ? T7656 : T7654;
  assign T7654 = T7655 ? counts_733 : counts_732;
  assign T7655 = T6203[1'h0:1'h0];
  assign T7656 = T7657 ? counts_735 : counts_734;
  assign T7657 = T6203[1'h0:1'h0];
  assign T7658 = T6203[1'h1:1'h1];
  assign T7659 = T6203[2'h2:2'h2];
  assign T7660 = T6203[2'h3:2'h3];
  assign T7661 = T6203[3'h4:3'h4];
  assign T7662 = T7723 ? T7693 : T7663;
  assign T7663 = T7692 ? T7678 : T7664;
  assign T7664 = T7677 ? T7671 : T7665;
  assign T7665 = T7670 ? T7668 : T7666;
  assign T7666 = T7667 ? counts_737 : counts_736;
  assign T7667 = T6203[1'h0:1'h0];
  assign T7668 = T7669 ? counts_739 : counts_738;
  assign T7669 = T6203[1'h0:1'h0];
  assign T7670 = T6203[1'h1:1'h1];
  assign T7671 = T7676 ? T7674 : T7672;
  assign T7672 = T7673 ? counts_741 : counts_740;
  assign T7673 = T6203[1'h0:1'h0];
  assign T7674 = T7675 ? counts_743 : counts_742;
  assign T7675 = T6203[1'h0:1'h0];
  assign T7676 = T6203[1'h1:1'h1];
  assign T7677 = T6203[2'h2:2'h2];
  assign T7678 = T7691 ? T7685 : T7679;
  assign T7679 = T7684 ? T7682 : T7680;
  assign T7680 = T7681 ? counts_745 : counts_744;
  assign T7681 = T6203[1'h0:1'h0];
  assign T7682 = T7683 ? counts_747 : counts_746;
  assign T7683 = T6203[1'h0:1'h0];
  assign T7684 = T6203[1'h1:1'h1];
  assign T7685 = T7690 ? T7688 : T7686;
  assign T7686 = T7687 ? counts_749 : counts_748;
  assign T7687 = T6203[1'h0:1'h0];
  assign T7688 = T7689 ? counts_751 : counts_750;
  assign T7689 = T6203[1'h0:1'h0];
  assign T7690 = T6203[1'h1:1'h1];
  assign T7691 = T6203[2'h2:2'h2];
  assign T7692 = T6203[2'h3:2'h3];
  assign T7693 = T7722 ? T7708 : T7694;
  assign T7694 = T7707 ? T7701 : T7695;
  assign T7695 = T7700 ? T7698 : T7696;
  assign T7696 = T7697 ? counts_753 : counts_752;
  assign T7697 = T6203[1'h0:1'h0];
  assign T7698 = T7699 ? counts_755 : counts_754;
  assign T7699 = T6203[1'h0:1'h0];
  assign T7700 = T6203[1'h1:1'h1];
  assign T7701 = T7706 ? T7704 : T7702;
  assign T7702 = T7703 ? counts_757 : counts_756;
  assign T7703 = T6203[1'h0:1'h0];
  assign T7704 = T7705 ? counts_759 : counts_758;
  assign T7705 = T6203[1'h0:1'h0];
  assign T7706 = T6203[1'h1:1'h1];
  assign T7707 = T6203[2'h2:2'h2];
  assign T7708 = T7721 ? T7715 : T7709;
  assign T7709 = T7714 ? T7712 : T7710;
  assign T7710 = T7711 ? counts_761 : counts_760;
  assign T7711 = T6203[1'h0:1'h0];
  assign T7712 = T7713 ? counts_763 : counts_762;
  assign T7713 = T6203[1'h0:1'h0];
  assign T7714 = T6203[1'h1:1'h1];
  assign T7715 = T7720 ? T7718 : T7716;
  assign T7716 = T7717 ? counts_765 : counts_764;
  assign T7717 = T6203[1'h0:1'h0];
  assign T7718 = T7719 ? counts_767 : counts_766;
  assign T7719 = T6203[1'h0:1'h0];
  assign T7720 = T6203[1'h1:1'h1];
  assign T7721 = T6203[2'h2:2'h2];
  assign T7722 = T6203[2'h3:2'h3];
  assign T7723 = T6203[3'h4:3'h4];
  assign T7724 = T6203[3'h5:3'h5];
  assign T7725 = T6203[3'h6:3'h6];
  assign T7726 = T6203[3'h7:3'h7];
  assign T7727 = T8236 ? T7982 : T7728;
  assign T7728 = T7981 ? T7855 : T7729;
  assign T7729 = T7854 ? T7792 : T7730;
  assign T7730 = T7791 ? T7761 : T7731;
  assign T7731 = T7760 ? T7746 : T7732;
  assign T7732 = T7745 ? T7739 : T7733;
  assign T7733 = T7738 ? T7736 : T7734;
  assign T7734 = T7735 ? counts_769 : counts_768;
  assign T7735 = T6203[1'h0:1'h0];
  assign T7736 = T7737 ? counts_771 : counts_770;
  assign T7737 = T6203[1'h0:1'h0];
  assign T7738 = T6203[1'h1:1'h1];
  assign T7739 = T7744 ? T7742 : T7740;
  assign T7740 = T7741 ? counts_773 : counts_772;
  assign T7741 = T6203[1'h0:1'h0];
  assign T7742 = T7743 ? counts_775 : counts_774;
  assign T7743 = T6203[1'h0:1'h0];
  assign T7744 = T6203[1'h1:1'h1];
  assign T7745 = T6203[2'h2:2'h2];
  assign T7746 = T7759 ? T7753 : T7747;
  assign T7747 = T7752 ? T7750 : T7748;
  assign T7748 = T7749 ? counts_777 : counts_776;
  assign T7749 = T6203[1'h0:1'h0];
  assign T7750 = T7751 ? counts_779 : counts_778;
  assign T7751 = T6203[1'h0:1'h0];
  assign T7752 = T6203[1'h1:1'h1];
  assign T7753 = T7758 ? T7756 : T7754;
  assign T7754 = T7755 ? counts_781 : counts_780;
  assign T7755 = T6203[1'h0:1'h0];
  assign T7756 = T7757 ? counts_783 : counts_782;
  assign T7757 = T6203[1'h0:1'h0];
  assign T7758 = T6203[1'h1:1'h1];
  assign T7759 = T6203[2'h2:2'h2];
  assign T7760 = T6203[2'h3:2'h3];
  assign T7761 = T7790 ? T7776 : T7762;
  assign T7762 = T7775 ? T7769 : T7763;
  assign T7763 = T7768 ? T7766 : T7764;
  assign T7764 = T7765 ? counts_785 : counts_784;
  assign T7765 = T6203[1'h0:1'h0];
  assign T7766 = T7767 ? counts_787 : counts_786;
  assign T7767 = T6203[1'h0:1'h0];
  assign T7768 = T6203[1'h1:1'h1];
  assign T7769 = T7774 ? T7772 : T7770;
  assign T7770 = T7771 ? counts_789 : counts_788;
  assign T7771 = T6203[1'h0:1'h0];
  assign T7772 = T7773 ? counts_791 : counts_790;
  assign T7773 = T6203[1'h0:1'h0];
  assign T7774 = T6203[1'h1:1'h1];
  assign T7775 = T6203[2'h2:2'h2];
  assign T7776 = T7789 ? T7783 : T7777;
  assign T7777 = T7782 ? T7780 : T7778;
  assign T7778 = T7779 ? counts_793 : counts_792;
  assign T7779 = T6203[1'h0:1'h0];
  assign T7780 = T7781 ? counts_795 : counts_794;
  assign T7781 = T6203[1'h0:1'h0];
  assign T7782 = T6203[1'h1:1'h1];
  assign T7783 = T7788 ? T7786 : T7784;
  assign T7784 = T7785 ? counts_797 : counts_796;
  assign T7785 = T6203[1'h0:1'h0];
  assign T7786 = T7787 ? counts_799 : counts_798;
  assign T7787 = T6203[1'h0:1'h0];
  assign T7788 = T6203[1'h1:1'h1];
  assign T7789 = T6203[2'h2:2'h2];
  assign T7790 = T6203[2'h3:2'h3];
  assign T7791 = T6203[3'h4:3'h4];
  assign T7792 = T7853 ? T7823 : T7793;
  assign T7793 = T7822 ? T7808 : T7794;
  assign T7794 = T7807 ? T7801 : T7795;
  assign T7795 = T7800 ? T7798 : T7796;
  assign T7796 = T7797 ? counts_801 : counts_800;
  assign T7797 = T6203[1'h0:1'h0];
  assign T7798 = T7799 ? counts_803 : counts_802;
  assign T7799 = T6203[1'h0:1'h0];
  assign T7800 = T6203[1'h1:1'h1];
  assign T7801 = T7806 ? T7804 : T7802;
  assign T7802 = T7803 ? counts_805 : counts_804;
  assign T7803 = T6203[1'h0:1'h0];
  assign T7804 = T7805 ? counts_807 : counts_806;
  assign T7805 = T6203[1'h0:1'h0];
  assign T7806 = T6203[1'h1:1'h1];
  assign T7807 = T6203[2'h2:2'h2];
  assign T7808 = T7821 ? T7815 : T7809;
  assign T7809 = T7814 ? T7812 : T7810;
  assign T7810 = T7811 ? counts_809 : counts_808;
  assign T7811 = T6203[1'h0:1'h0];
  assign T7812 = T7813 ? counts_811 : counts_810;
  assign T7813 = T6203[1'h0:1'h0];
  assign T7814 = T6203[1'h1:1'h1];
  assign T7815 = T7820 ? T7818 : T7816;
  assign T7816 = T7817 ? counts_813 : counts_812;
  assign T7817 = T6203[1'h0:1'h0];
  assign T7818 = T7819 ? counts_815 : counts_814;
  assign T7819 = T6203[1'h0:1'h0];
  assign T7820 = T6203[1'h1:1'h1];
  assign T7821 = T6203[2'h2:2'h2];
  assign T7822 = T6203[2'h3:2'h3];
  assign T7823 = T7852 ? T7838 : T7824;
  assign T7824 = T7837 ? T7831 : T7825;
  assign T7825 = T7830 ? T7828 : T7826;
  assign T7826 = T7827 ? counts_817 : counts_816;
  assign T7827 = T6203[1'h0:1'h0];
  assign T7828 = T7829 ? counts_819 : counts_818;
  assign T7829 = T6203[1'h0:1'h0];
  assign T7830 = T6203[1'h1:1'h1];
  assign T7831 = T7836 ? T7834 : T7832;
  assign T7832 = T7833 ? counts_821 : counts_820;
  assign T7833 = T6203[1'h0:1'h0];
  assign T7834 = T7835 ? counts_823 : counts_822;
  assign T7835 = T6203[1'h0:1'h0];
  assign T7836 = T6203[1'h1:1'h1];
  assign T7837 = T6203[2'h2:2'h2];
  assign T7838 = T7851 ? T7845 : T7839;
  assign T7839 = T7844 ? T7842 : T7840;
  assign T7840 = T7841 ? counts_825 : counts_824;
  assign T7841 = T6203[1'h0:1'h0];
  assign T7842 = T7843 ? counts_827 : counts_826;
  assign T7843 = T6203[1'h0:1'h0];
  assign T7844 = T6203[1'h1:1'h1];
  assign T7845 = T7850 ? T7848 : T7846;
  assign T7846 = T7847 ? counts_829 : counts_828;
  assign T7847 = T6203[1'h0:1'h0];
  assign T7848 = T7849 ? counts_831 : counts_830;
  assign T7849 = T6203[1'h0:1'h0];
  assign T7850 = T6203[1'h1:1'h1];
  assign T7851 = T6203[2'h2:2'h2];
  assign T7852 = T6203[2'h3:2'h3];
  assign T7853 = T6203[3'h4:3'h4];
  assign T7854 = T6203[3'h5:3'h5];
  assign T7855 = T7980 ? T7918 : T7856;
  assign T7856 = T7917 ? T7887 : T7857;
  assign T7857 = T7886 ? T7872 : T7858;
  assign T7858 = T7871 ? T7865 : T7859;
  assign T7859 = T7864 ? T7862 : T7860;
  assign T7860 = T7861 ? counts_833 : counts_832;
  assign T7861 = T6203[1'h0:1'h0];
  assign T7862 = T7863 ? counts_835 : counts_834;
  assign T7863 = T6203[1'h0:1'h0];
  assign T7864 = T6203[1'h1:1'h1];
  assign T7865 = T7870 ? T7868 : T7866;
  assign T7866 = T7867 ? counts_837 : counts_836;
  assign T7867 = T6203[1'h0:1'h0];
  assign T7868 = T7869 ? counts_839 : counts_838;
  assign T7869 = T6203[1'h0:1'h0];
  assign T7870 = T6203[1'h1:1'h1];
  assign T7871 = T6203[2'h2:2'h2];
  assign T7872 = T7885 ? T7879 : T7873;
  assign T7873 = T7878 ? T7876 : T7874;
  assign T7874 = T7875 ? counts_841 : counts_840;
  assign T7875 = T6203[1'h0:1'h0];
  assign T7876 = T7877 ? counts_843 : counts_842;
  assign T7877 = T6203[1'h0:1'h0];
  assign T7878 = T6203[1'h1:1'h1];
  assign T7879 = T7884 ? T7882 : T7880;
  assign T7880 = T7881 ? counts_845 : counts_844;
  assign T7881 = T6203[1'h0:1'h0];
  assign T7882 = T7883 ? counts_847 : counts_846;
  assign T7883 = T6203[1'h0:1'h0];
  assign T7884 = T6203[1'h1:1'h1];
  assign T7885 = T6203[2'h2:2'h2];
  assign T7886 = T6203[2'h3:2'h3];
  assign T7887 = T7916 ? T7902 : T7888;
  assign T7888 = T7901 ? T7895 : T7889;
  assign T7889 = T7894 ? T7892 : T7890;
  assign T7890 = T7891 ? counts_849 : counts_848;
  assign T7891 = T6203[1'h0:1'h0];
  assign T7892 = T7893 ? counts_851 : counts_850;
  assign T7893 = T6203[1'h0:1'h0];
  assign T7894 = T6203[1'h1:1'h1];
  assign T7895 = T7900 ? T7898 : T7896;
  assign T7896 = T7897 ? counts_853 : counts_852;
  assign T7897 = T6203[1'h0:1'h0];
  assign T7898 = T7899 ? counts_855 : counts_854;
  assign T7899 = T6203[1'h0:1'h0];
  assign T7900 = T6203[1'h1:1'h1];
  assign T7901 = T6203[2'h2:2'h2];
  assign T7902 = T7915 ? T7909 : T7903;
  assign T7903 = T7908 ? T7906 : T7904;
  assign T7904 = T7905 ? counts_857 : counts_856;
  assign T7905 = T6203[1'h0:1'h0];
  assign T7906 = T7907 ? counts_859 : counts_858;
  assign T7907 = T6203[1'h0:1'h0];
  assign T7908 = T6203[1'h1:1'h1];
  assign T7909 = T7914 ? T7912 : T7910;
  assign T7910 = T7911 ? counts_861 : counts_860;
  assign T7911 = T6203[1'h0:1'h0];
  assign T7912 = T7913 ? counts_863 : counts_862;
  assign T7913 = T6203[1'h0:1'h0];
  assign T7914 = T6203[1'h1:1'h1];
  assign T7915 = T6203[2'h2:2'h2];
  assign T7916 = T6203[2'h3:2'h3];
  assign T7917 = T6203[3'h4:3'h4];
  assign T7918 = T7979 ? T7949 : T7919;
  assign T7919 = T7948 ? T7934 : T7920;
  assign T7920 = T7933 ? T7927 : T7921;
  assign T7921 = T7926 ? T7924 : T7922;
  assign T7922 = T7923 ? counts_865 : counts_864;
  assign T7923 = T6203[1'h0:1'h0];
  assign T7924 = T7925 ? counts_867 : counts_866;
  assign T7925 = T6203[1'h0:1'h0];
  assign T7926 = T6203[1'h1:1'h1];
  assign T7927 = T7932 ? T7930 : T7928;
  assign T7928 = T7929 ? counts_869 : counts_868;
  assign T7929 = T6203[1'h0:1'h0];
  assign T7930 = T7931 ? counts_871 : counts_870;
  assign T7931 = T6203[1'h0:1'h0];
  assign T7932 = T6203[1'h1:1'h1];
  assign T7933 = T6203[2'h2:2'h2];
  assign T7934 = T7947 ? T7941 : T7935;
  assign T7935 = T7940 ? T7938 : T7936;
  assign T7936 = T7937 ? counts_873 : counts_872;
  assign T7937 = T6203[1'h0:1'h0];
  assign T7938 = T7939 ? counts_875 : counts_874;
  assign T7939 = T6203[1'h0:1'h0];
  assign T7940 = T6203[1'h1:1'h1];
  assign T7941 = T7946 ? T7944 : T7942;
  assign T7942 = T7943 ? counts_877 : counts_876;
  assign T7943 = T6203[1'h0:1'h0];
  assign T7944 = T7945 ? counts_879 : counts_878;
  assign T7945 = T6203[1'h0:1'h0];
  assign T7946 = T6203[1'h1:1'h1];
  assign T7947 = T6203[2'h2:2'h2];
  assign T7948 = T6203[2'h3:2'h3];
  assign T7949 = T7978 ? T7964 : T7950;
  assign T7950 = T7963 ? T7957 : T7951;
  assign T7951 = T7956 ? T7954 : T7952;
  assign T7952 = T7953 ? counts_881 : counts_880;
  assign T7953 = T6203[1'h0:1'h0];
  assign T7954 = T7955 ? counts_883 : counts_882;
  assign T7955 = T6203[1'h0:1'h0];
  assign T7956 = T6203[1'h1:1'h1];
  assign T7957 = T7962 ? T7960 : T7958;
  assign T7958 = T7959 ? counts_885 : counts_884;
  assign T7959 = T6203[1'h0:1'h0];
  assign T7960 = T7961 ? counts_887 : counts_886;
  assign T7961 = T6203[1'h0:1'h0];
  assign T7962 = T6203[1'h1:1'h1];
  assign T7963 = T6203[2'h2:2'h2];
  assign T7964 = T7977 ? T7971 : T7965;
  assign T7965 = T7970 ? T7968 : T7966;
  assign T7966 = T7967 ? counts_889 : counts_888;
  assign T7967 = T6203[1'h0:1'h0];
  assign T7968 = T7969 ? counts_891 : counts_890;
  assign T7969 = T6203[1'h0:1'h0];
  assign T7970 = T6203[1'h1:1'h1];
  assign T7971 = T7976 ? T7974 : T7972;
  assign T7972 = T7973 ? counts_893 : counts_892;
  assign T7973 = T6203[1'h0:1'h0];
  assign T7974 = T7975 ? counts_895 : counts_894;
  assign T7975 = T6203[1'h0:1'h0];
  assign T7976 = T6203[1'h1:1'h1];
  assign T7977 = T6203[2'h2:2'h2];
  assign T7978 = T6203[2'h3:2'h3];
  assign T7979 = T6203[3'h4:3'h4];
  assign T7980 = T6203[3'h5:3'h5];
  assign T7981 = T6203[3'h6:3'h6];
  assign T7982 = T8235 ? T8109 : T7983;
  assign T7983 = T8108 ? T8046 : T7984;
  assign T7984 = T8045 ? T8015 : T7985;
  assign T7985 = T8014 ? T8000 : T7986;
  assign T7986 = T7999 ? T7993 : T7987;
  assign T7987 = T7992 ? T7990 : T7988;
  assign T7988 = T7989 ? counts_897 : counts_896;
  assign T7989 = T6203[1'h0:1'h0];
  assign T7990 = T7991 ? counts_899 : counts_898;
  assign T7991 = T6203[1'h0:1'h0];
  assign T7992 = T6203[1'h1:1'h1];
  assign T7993 = T7998 ? T7996 : T7994;
  assign T7994 = T7995 ? counts_901 : counts_900;
  assign T7995 = T6203[1'h0:1'h0];
  assign T7996 = T7997 ? counts_903 : counts_902;
  assign T7997 = T6203[1'h0:1'h0];
  assign T7998 = T6203[1'h1:1'h1];
  assign T7999 = T6203[2'h2:2'h2];
  assign T8000 = T8013 ? T8007 : T8001;
  assign T8001 = T8006 ? T8004 : T8002;
  assign T8002 = T8003 ? counts_905 : counts_904;
  assign T8003 = T6203[1'h0:1'h0];
  assign T8004 = T8005 ? counts_907 : counts_906;
  assign T8005 = T6203[1'h0:1'h0];
  assign T8006 = T6203[1'h1:1'h1];
  assign T8007 = T8012 ? T8010 : T8008;
  assign T8008 = T8009 ? counts_909 : counts_908;
  assign T8009 = T6203[1'h0:1'h0];
  assign T8010 = T8011 ? counts_911 : counts_910;
  assign T8011 = T6203[1'h0:1'h0];
  assign T8012 = T6203[1'h1:1'h1];
  assign T8013 = T6203[2'h2:2'h2];
  assign T8014 = T6203[2'h3:2'h3];
  assign T8015 = T8044 ? T8030 : T8016;
  assign T8016 = T8029 ? T8023 : T8017;
  assign T8017 = T8022 ? T8020 : T8018;
  assign T8018 = T8019 ? counts_913 : counts_912;
  assign T8019 = T6203[1'h0:1'h0];
  assign T8020 = T8021 ? counts_915 : counts_914;
  assign T8021 = T6203[1'h0:1'h0];
  assign T8022 = T6203[1'h1:1'h1];
  assign T8023 = T8028 ? T8026 : T8024;
  assign T8024 = T8025 ? counts_917 : counts_916;
  assign T8025 = T6203[1'h0:1'h0];
  assign T8026 = T8027 ? counts_919 : counts_918;
  assign T8027 = T6203[1'h0:1'h0];
  assign T8028 = T6203[1'h1:1'h1];
  assign T8029 = T6203[2'h2:2'h2];
  assign T8030 = T8043 ? T8037 : T8031;
  assign T8031 = T8036 ? T8034 : T8032;
  assign T8032 = T8033 ? counts_921 : counts_920;
  assign T8033 = T6203[1'h0:1'h0];
  assign T8034 = T8035 ? counts_923 : counts_922;
  assign T8035 = T6203[1'h0:1'h0];
  assign T8036 = T6203[1'h1:1'h1];
  assign T8037 = T8042 ? T8040 : T8038;
  assign T8038 = T8039 ? counts_925 : counts_924;
  assign T8039 = T6203[1'h0:1'h0];
  assign T8040 = T8041 ? counts_927 : counts_926;
  assign T8041 = T6203[1'h0:1'h0];
  assign T8042 = T6203[1'h1:1'h1];
  assign T8043 = T6203[2'h2:2'h2];
  assign T8044 = T6203[2'h3:2'h3];
  assign T8045 = T6203[3'h4:3'h4];
  assign T8046 = T8107 ? T8077 : T8047;
  assign T8047 = T8076 ? T8062 : T8048;
  assign T8048 = T8061 ? T8055 : T8049;
  assign T8049 = T8054 ? T8052 : T8050;
  assign T8050 = T8051 ? counts_929 : counts_928;
  assign T8051 = T6203[1'h0:1'h0];
  assign T8052 = T8053 ? counts_931 : counts_930;
  assign T8053 = T6203[1'h0:1'h0];
  assign T8054 = T6203[1'h1:1'h1];
  assign T8055 = T8060 ? T8058 : T8056;
  assign T8056 = T8057 ? counts_933 : counts_932;
  assign T8057 = T6203[1'h0:1'h0];
  assign T8058 = T8059 ? counts_935 : counts_934;
  assign T8059 = T6203[1'h0:1'h0];
  assign T8060 = T6203[1'h1:1'h1];
  assign T8061 = T6203[2'h2:2'h2];
  assign T8062 = T8075 ? T8069 : T8063;
  assign T8063 = T8068 ? T8066 : T8064;
  assign T8064 = T8065 ? counts_937 : counts_936;
  assign T8065 = T6203[1'h0:1'h0];
  assign T8066 = T8067 ? counts_939 : counts_938;
  assign T8067 = T6203[1'h0:1'h0];
  assign T8068 = T6203[1'h1:1'h1];
  assign T8069 = T8074 ? T8072 : T8070;
  assign T8070 = T8071 ? counts_941 : counts_940;
  assign T8071 = T6203[1'h0:1'h0];
  assign T8072 = T8073 ? counts_943 : counts_942;
  assign T8073 = T6203[1'h0:1'h0];
  assign T8074 = T6203[1'h1:1'h1];
  assign T8075 = T6203[2'h2:2'h2];
  assign T8076 = T6203[2'h3:2'h3];
  assign T8077 = T8106 ? T8092 : T8078;
  assign T8078 = T8091 ? T8085 : T8079;
  assign T8079 = T8084 ? T8082 : T8080;
  assign T8080 = T8081 ? counts_945 : counts_944;
  assign T8081 = T6203[1'h0:1'h0];
  assign T8082 = T8083 ? counts_947 : counts_946;
  assign T8083 = T6203[1'h0:1'h0];
  assign T8084 = T6203[1'h1:1'h1];
  assign T8085 = T8090 ? T8088 : T8086;
  assign T8086 = T8087 ? counts_949 : counts_948;
  assign T8087 = T6203[1'h0:1'h0];
  assign T8088 = T8089 ? counts_951 : counts_950;
  assign T8089 = T6203[1'h0:1'h0];
  assign T8090 = T6203[1'h1:1'h1];
  assign T8091 = T6203[2'h2:2'h2];
  assign T8092 = T8105 ? T8099 : T8093;
  assign T8093 = T8098 ? T8096 : T8094;
  assign T8094 = T8095 ? counts_953 : counts_952;
  assign T8095 = T6203[1'h0:1'h0];
  assign T8096 = T8097 ? counts_955 : counts_954;
  assign T8097 = T6203[1'h0:1'h0];
  assign T8098 = T6203[1'h1:1'h1];
  assign T8099 = T8104 ? T8102 : T8100;
  assign T8100 = T8101 ? counts_957 : counts_956;
  assign T8101 = T6203[1'h0:1'h0];
  assign T8102 = T8103 ? counts_959 : counts_958;
  assign T8103 = T6203[1'h0:1'h0];
  assign T8104 = T6203[1'h1:1'h1];
  assign T8105 = T6203[2'h2:2'h2];
  assign T8106 = T6203[2'h3:2'h3];
  assign T8107 = T6203[3'h4:3'h4];
  assign T8108 = T6203[3'h5:3'h5];
  assign T8109 = T8234 ? T8172 : T8110;
  assign T8110 = T8171 ? T8141 : T8111;
  assign T8111 = T8140 ? T8126 : T8112;
  assign T8112 = T8125 ? T8119 : T8113;
  assign T8113 = T8118 ? T8116 : T8114;
  assign T8114 = T8115 ? counts_961 : counts_960;
  assign T8115 = T6203[1'h0:1'h0];
  assign T8116 = T8117 ? counts_963 : counts_962;
  assign T8117 = T6203[1'h0:1'h0];
  assign T8118 = T6203[1'h1:1'h1];
  assign T8119 = T8124 ? T8122 : T8120;
  assign T8120 = T8121 ? counts_965 : counts_964;
  assign T8121 = T6203[1'h0:1'h0];
  assign T8122 = T8123 ? counts_967 : counts_966;
  assign T8123 = T6203[1'h0:1'h0];
  assign T8124 = T6203[1'h1:1'h1];
  assign T8125 = T6203[2'h2:2'h2];
  assign T8126 = T8139 ? T8133 : T8127;
  assign T8127 = T8132 ? T8130 : T8128;
  assign T8128 = T8129 ? counts_969 : counts_968;
  assign T8129 = T6203[1'h0:1'h0];
  assign T8130 = T8131 ? counts_971 : counts_970;
  assign T8131 = T6203[1'h0:1'h0];
  assign T8132 = T6203[1'h1:1'h1];
  assign T8133 = T8138 ? T8136 : T8134;
  assign T8134 = T8135 ? counts_973 : counts_972;
  assign T8135 = T6203[1'h0:1'h0];
  assign T8136 = T8137 ? counts_975 : counts_974;
  assign T8137 = T6203[1'h0:1'h0];
  assign T8138 = T6203[1'h1:1'h1];
  assign T8139 = T6203[2'h2:2'h2];
  assign T8140 = T6203[2'h3:2'h3];
  assign T8141 = T8170 ? T8156 : T8142;
  assign T8142 = T8155 ? T8149 : T8143;
  assign T8143 = T8148 ? T8146 : T8144;
  assign T8144 = T8145 ? counts_977 : counts_976;
  assign T8145 = T6203[1'h0:1'h0];
  assign T8146 = T8147 ? counts_979 : counts_978;
  assign T8147 = T6203[1'h0:1'h0];
  assign T8148 = T6203[1'h1:1'h1];
  assign T8149 = T8154 ? T8152 : T8150;
  assign T8150 = T8151 ? counts_981 : counts_980;
  assign T8151 = T6203[1'h0:1'h0];
  assign T8152 = T8153 ? counts_983 : counts_982;
  assign T8153 = T6203[1'h0:1'h0];
  assign T8154 = T6203[1'h1:1'h1];
  assign T8155 = T6203[2'h2:2'h2];
  assign T8156 = T8169 ? T8163 : T8157;
  assign T8157 = T8162 ? T8160 : T8158;
  assign T8158 = T8159 ? counts_985 : counts_984;
  assign T8159 = T6203[1'h0:1'h0];
  assign T8160 = T8161 ? counts_987 : counts_986;
  assign T8161 = T6203[1'h0:1'h0];
  assign T8162 = T6203[1'h1:1'h1];
  assign T8163 = T8168 ? T8166 : T8164;
  assign T8164 = T8165 ? counts_989 : counts_988;
  assign T8165 = T6203[1'h0:1'h0];
  assign T8166 = T8167 ? counts_991 : counts_990;
  assign T8167 = T6203[1'h0:1'h0];
  assign T8168 = T6203[1'h1:1'h1];
  assign T8169 = T6203[2'h2:2'h2];
  assign T8170 = T6203[2'h3:2'h3];
  assign T8171 = T6203[3'h4:3'h4];
  assign T8172 = T8233 ? T8203 : T8173;
  assign T8173 = T8202 ? T8188 : T8174;
  assign T8174 = T8187 ? T8181 : T8175;
  assign T8175 = T8180 ? T8178 : T8176;
  assign T8176 = T8177 ? counts_993 : counts_992;
  assign T8177 = T6203[1'h0:1'h0];
  assign T8178 = T8179 ? counts_995 : counts_994;
  assign T8179 = T6203[1'h0:1'h0];
  assign T8180 = T6203[1'h1:1'h1];
  assign T8181 = T8186 ? T8184 : T8182;
  assign T8182 = T8183 ? counts_997 : counts_996;
  assign T8183 = T6203[1'h0:1'h0];
  assign T8184 = T8185 ? counts_999 : counts_998;
  assign T8185 = T6203[1'h0:1'h0];
  assign T8186 = T6203[1'h1:1'h1];
  assign T8187 = T6203[2'h2:2'h2];
  assign T8188 = T8201 ? T8195 : T8189;
  assign T8189 = T8194 ? T8192 : T8190;
  assign T8190 = T8191 ? counts_1001 : counts_1000;
  assign T8191 = T6203[1'h0:1'h0];
  assign T8192 = T8193 ? counts_1003 : counts_1002;
  assign T8193 = T6203[1'h0:1'h0];
  assign T8194 = T6203[1'h1:1'h1];
  assign T8195 = T8200 ? T8198 : T8196;
  assign T8196 = T8197 ? counts_1005 : counts_1004;
  assign T8197 = T6203[1'h0:1'h0];
  assign T8198 = T8199 ? counts_1007 : counts_1006;
  assign T8199 = T6203[1'h0:1'h0];
  assign T8200 = T6203[1'h1:1'h1];
  assign T8201 = T6203[2'h2:2'h2];
  assign T8202 = T6203[2'h3:2'h3];
  assign T8203 = T8232 ? T8218 : T8204;
  assign T8204 = T8217 ? T8211 : T8205;
  assign T8205 = T8210 ? T8208 : T8206;
  assign T8206 = T8207 ? counts_1009 : counts_1008;
  assign T8207 = T6203[1'h0:1'h0];
  assign T8208 = T8209 ? counts_1011 : counts_1010;
  assign T8209 = T6203[1'h0:1'h0];
  assign T8210 = T6203[1'h1:1'h1];
  assign T8211 = T8216 ? T8214 : T8212;
  assign T8212 = T8213 ? counts_1013 : counts_1012;
  assign T8213 = T6203[1'h0:1'h0];
  assign T8214 = T8215 ? counts_1015 : counts_1014;
  assign T8215 = T6203[1'h0:1'h0];
  assign T8216 = T6203[1'h1:1'h1];
  assign T8217 = T6203[2'h2:2'h2];
  assign T8218 = T8231 ? T8225 : T8219;
  assign T8219 = T8224 ? T8222 : T8220;
  assign T8220 = T8221 ? counts_1017 : counts_1016;
  assign T8221 = T6203[1'h0:1'h0];
  assign T8222 = T8223 ? counts_1019 : counts_1018;
  assign T8223 = T6203[1'h0:1'h0];
  assign T8224 = T6203[1'h1:1'h1];
  assign T8225 = T8230 ? T8228 : T8226;
  assign T8226 = T8227 ? counts_1021 : counts_1020;
  assign T8227 = T6203[1'h0:1'h0];
  assign T8228 = T8229 ? counts_1023 : counts_1022;
  assign T8229 = T6203[1'h0:1'h0];
  assign T8230 = T6203[1'h1:1'h1];
  assign T8231 = T6203[2'h2:2'h2];
  assign T8232 = T6203[2'h3:2'h3];
  assign T8233 = T6203[3'h4:3'h4];
  assign T8234 = T6203[3'h5:3'h5];
  assign T8235 = T6203[3'h6:3'h6];
  assign T8236 = T6203[3'h7:3'h7];
  assign T8237 = T6203[4'h8:4'h8];
  assign T8238 = T6203[4'h9:4'h9];
  assign T11370 = reset ? 4'h0 : T8239;
  assign T8239 = T21 ? T8240 : hashCount1;
  assign T8240 = T10286 ? T9264 : T8241;
  assign T8241 = T9263 ? T8753 : T8242;
  assign T8242 = T8752 ? T8498 : T8243;
  assign T8243 = T8497 ? T8371 : T8244;
  assign T8244 = T8370 ? T8308 : T8245;
  assign T8245 = T8307 ? T8277 : T8246;
  assign T8246 = T8276 ? T8262 : T8247;
  assign T8247 = T8261 ? T8255 : T8248;
  assign T8248 = T8254 ? T8252 : T8249;
  assign T8249 = T8250 ? counts_1 : counts_0;
  assign T8250 = T8251[1'h0:1'h0];
  assign T8251 = curInfo_hash1;
  assign T8252 = T8253 ? counts_3 : counts_2;
  assign T8253 = T8251[1'h0:1'h0];
  assign T8254 = T8251[1'h1:1'h1];
  assign T8255 = T8260 ? T8258 : T8256;
  assign T8256 = T8257 ? counts_5 : counts_4;
  assign T8257 = T8251[1'h0:1'h0];
  assign T8258 = T8259 ? counts_7 : counts_6;
  assign T8259 = T8251[1'h0:1'h0];
  assign T8260 = T8251[1'h1:1'h1];
  assign T8261 = T8251[2'h2:2'h2];
  assign T8262 = T8275 ? T8269 : T8263;
  assign T8263 = T8268 ? T8266 : T8264;
  assign T8264 = T8265 ? counts_9 : counts_8;
  assign T8265 = T8251[1'h0:1'h0];
  assign T8266 = T8267 ? counts_11 : counts_10;
  assign T8267 = T8251[1'h0:1'h0];
  assign T8268 = T8251[1'h1:1'h1];
  assign T8269 = T8274 ? T8272 : T8270;
  assign T8270 = T8271 ? counts_13 : counts_12;
  assign T8271 = T8251[1'h0:1'h0];
  assign T8272 = T8273 ? counts_15 : counts_14;
  assign T8273 = T8251[1'h0:1'h0];
  assign T8274 = T8251[1'h1:1'h1];
  assign T8275 = T8251[2'h2:2'h2];
  assign T8276 = T8251[2'h3:2'h3];
  assign T8277 = T8306 ? T8292 : T8278;
  assign T8278 = T8291 ? T8285 : T8279;
  assign T8279 = T8284 ? T8282 : T8280;
  assign T8280 = T8281 ? counts_17 : counts_16;
  assign T8281 = T8251[1'h0:1'h0];
  assign T8282 = T8283 ? counts_19 : counts_18;
  assign T8283 = T8251[1'h0:1'h0];
  assign T8284 = T8251[1'h1:1'h1];
  assign T8285 = T8290 ? T8288 : T8286;
  assign T8286 = T8287 ? counts_21 : counts_20;
  assign T8287 = T8251[1'h0:1'h0];
  assign T8288 = T8289 ? counts_23 : counts_22;
  assign T8289 = T8251[1'h0:1'h0];
  assign T8290 = T8251[1'h1:1'h1];
  assign T8291 = T8251[2'h2:2'h2];
  assign T8292 = T8305 ? T8299 : T8293;
  assign T8293 = T8298 ? T8296 : T8294;
  assign T8294 = T8295 ? counts_25 : counts_24;
  assign T8295 = T8251[1'h0:1'h0];
  assign T8296 = T8297 ? counts_27 : counts_26;
  assign T8297 = T8251[1'h0:1'h0];
  assign T8298 = T8251[1'h1:1'h1];
  assign T8299 = T8304 ? T8302 : T8300;
  assign T8300 = T8301 ? counts_29 : counts_28;
  assign T8301 = T8251[1'h0:1'h0];
  assign T8302 = T8303 ? counts_31 : counts_30;
  assign T8303 = T8251[1'h0:1'h0];
  assign T8304 = T8251[1'h1:1'h1];
  assign T8305 = T8251[2'h2:2'h2];
  assign T8306 = T8251[2'h3:2'h3];
  assign T8307 = T8251[3'h4:3'h4];
  assign T8308 = T8369 ? T8339 : T8309;
  assign T8309 = T8338 ? T8324 : T8310;
  assign T8310 = T8323 ? T8317 : T8311;
  assign T8311 = T8316 ? T8314 : T8312;
  assign T8312 = T8313 ? counts_33 : counts_32;
  assign T8313 = T8251[1'h0:1'h0];
  assign T8314 = T8315 ? counts_35 : counts_34;
  assign T8315 = T8251[1'h0:1'h0];
  assign T8316 = T8251[1'h1:1'h1];
  assign T8317 = T8322 ? T8320 : T8318;
  assign T8318 = T8319 ? counts_37 : counts_36;
  assign T8319 = T8251[1'h0:1'h0];
  assign T8320 = T8321 ? counts_39 : counts_38;
  assign T8321 = T8251[1'h0:1'h0];
  assign T8322 = T8251[1'h1:1'h1];
  assign T8323 = T8251[2'h2:2'h2];
  assign T8324 = T8337 ? T8331 : T8325;
  assign T8325 = T8330 ? T8328 : T8326;
  assign T8326 = T8327 ? counts_41 : counts_40;
  assign T8327 = T8251[1'h0:1'h0];
  assign T8328 = T8329 ? counts_43 : counts_42;
  assign T8329 = T8251[1'h0:1'h0];
  assign T8330 = T8251[1'h1:1'h1];
  assign T8331 = T8336 ? T8334 : T8332;
  assign T8332 = T8333 ? counts_45 : counts_44;
  assign T8333 = T8251[1'h0:1'h0];
  assign T8334 = T8335 ? counts_47 : counts_46;
  assign T8335 = T8251[1'h0:1'h0];
  assign T8336 = T8251[1'h1:1'h1];
  assign T8337 = T8251[2'h2:2'h2];
  assign T8338 = T8251[2'h3:2'h3];
  assign T8339 = T8368 ? T8354 : T8340;
  assign T8340 = T8353 ? T8347 : T8341;
  assign T8341 = T8346 ? T8344 : T8342;
  assign T8342 = T8343 ? counts_49 : counts_48;
  assign T8343 = T8251[1'h0:1'h0];
  assign T8344 = T8345 ? counts_51 : counts_50;
  assign T8345 = T8251[1'h0:1'h0];
  assign T8346 = T8251[1'h1:1'h1];
  assign T8347 = T8352 ? T8350 : T8348;
  assign T8348 = T8349 ? counts_53 : counts_52;
  assign T8349 = T8251[1'h0:1'h0];
  assign T8350 = T8351 ? counts_55 : counts_54;
  assign T8351 = T8251[1'h0:1'h0];
  assign T8352 = T8251[1'h1:1'h1];
  assign T8353 = T8251[2'h2:2'h2];
  assign T8354 = T8367 ? T8361 : T8355;
  assign T8355 = T8360 ? T8358 : T8356;
  assign T8356 = T8357 ? counts_57 : counts_56;
  assign T8357 = T8251[1'h0:1'h0];
  assign T8358 = T8359 ? counts_59 : counts_58;
  assign T8359 = T8251[1'h0:1'h0];
  assign T8360 = T8251[1'h1:1'h1];
  assign T8361 = T8366 ? T8364 : T8362;
  assign T8362 = T8363 ? counts_61 : counts_60;
  assign T8363 = T8251[1'h0:1'h0];
  assign T8364 = T8365 ? counts_63 : counts_62;
  assign T8365 = T8251[1'h0:1'h0];
  assign T8366 = T8251[1'h1:1'h1];
  assign T8367 = T8251[2'h2:2'h2];
  assign T8368 = T8251[2'h3:2'h3];
  assign T8369 = T8251[3'h4:3'h4];
  assign T8370 = T8251[3'h5:3'h5];
  assign T8371 = T8496 ? T8434 : T8372;
  assign T8372 = T8433 ? T8403 : T8373;
  assign T8373 = T8402 ? T8388 : T8374;
  assign T8374 = T8387 ? T8381 : T8375;
  assign T8375 = T8380 ? T8378 : T8376;
  assign T8376 = T8377 ? counts_65 : counts_64;
  assign T8377 = T8251[1'h0:1'h0];
  assign T8378 = T8379 ? counts_67 : counts_66;
  assign T8379 = T8251[1'h0:1'h0];
  assign T8380 = T8251[1'h1:1'h1];
  assign T8381 = T8386 ? T8384 : T8382;
  assign T8382 = T8383 ? counts_69 : counts_68;
  assign T8383 = T8251[1'h0:1'h0];
  assign T8384 = T8385 ? counts_71 : counts_70;
  assign T8385 = T8251[1'h0:1'h0];
  assign T8386 = T8251[1'h1:1'h1];
  assign T8387 = T8251[2'h2:2'h2];
  assign T8388 = T8401 ? T8395 : T8389;
  assign T8389 = T8394 ? T8392 : T8390;
  assign T8390 = T8391 ? counts_73 : counts_72;
  assign T8391 = T8251[1'h0:1'h0];
  assign T8392 = T8393 ? counts_75 : counts_74;
  assign T8393 = T8251[1'h0:1'h0];
  assign T8394 = T8251[1'h1:1'h1];
  assign T8395 = T8400 ? T8398 : T8396;
  assign T8396 = T8397 ? counts_77 : counts_76;
  assign T8397 = T8251[1'h0:1'h0];
  assign T8398 = T8399 ? counts_79 : counts_78;
  assign T8399 = T8251[1'h0:1'h0];
  assign T8400 = T8251[1'h1:1'h1];
  assign T8401 = T8251[2'h2:2'h2];
  assign T8402 = T8251[2'h3:2'h3];
  assign T8403 = T8432 ? T8418 : T8404;
  assign T8404 = T8417 ? T8411 : T8405;
  assign T8405 = T8410 ? T8408 : T8406;
  assign T8406 = T8407 ? counts_81 : counts_80;
  assign T8407 = T8251[1'h0:1'h0];
  assign T8408 = T8409 ? counts_83 : counts_82;
  assign T8409 = T8251[1'h0:1'h0];
  assign T8410 = T8251[1'h1:1'h1];
  assign T8411 = T8416 ? T8414 : T8412;
  assign T8412 = T8413 ? counts_85 : counts_84;
  assign T8413 = T8251[1'h0:1'h0];
  assign T8414 = T8415 ? counts_87 : counts_86;
  assign T8415 = T8251[1'h0:1'h0];
  assign T8416 = T8251[1'h1:1'h1];
  assign T8417 = T8251[2'h2:2'h2];
  assign T8418 = T8431 ? T8425 : T8419;
  assign T8419 = T8424 ? T8422 : T8420;
  assign T8420 = T8421 ? counts_89 : counts_88;
  assign T8421 = T8251[1'h0:1'h0];
  assign T8422 = T8423 ? counts_91 : counts_90;
  assign T8423 = T8251[1'h0:1'h0];
  assign T8424 = T8251[1'h1:1'h1];
  assign T8425 = T8430 ? T8428 : T8426;
  assign T8426 = T8427 ? counts_93 : counts_92;
  assign T8427 = T8251[1'h0:1'h0];
  assign T8428 = T8429 ? counts_95 : counts_94;
  assign T8429 = T8251[1'h0:1'h0];
  assign T8430 = T8251[1'h1:1'h1];
  assign T8431 = T8251[2'h2:2'h2];
  assign T8432 = T8251[2'h3:2'h3];
  assign T8433 = T8251[3'h4:3'h4];
  assign T8434 = T8495 ? T8465 : T8435;
  assign T8435 = T8464 ? T8450 : T8436;
  assign T8436 = T8449 ? T8443 : T8437;
  assign T8437 = T8442 ? T8440 : T8438;
  assign T8438 = T8439 ? counts_97 : counts_96;
  assign T8439 = T8251[1'h0:1'h0];
  assign T8440 = T8441 ? counts_99 : counts_98;
  assign T8441 = T8251[1'h0:1'h0];
  assign T8442 = T8251[1'h1:1'h1];
  assign T8443 = T8448 ? T8446 : T8444;
  assign T8444 = T8445 ? counts_101 : counts_100;
  assign T8445 = T8251[1'h0:1'h0];
  assign T8446 = T8447 ? counts_103 : counts_102;
  assign T8447 = T8251[1'h0:1'h0];
  assign T8448 = T8251[1'h1:1'h1];
  assign T8449 = T8251[2'h2:2'h2];
  assign T8450 = T8463 ? T8457 : T8451;
  assign T8451 = T8456 ? T8454 : T8452;
  assign T8452 = T8453 ? counts_105 : counts_104;
  assign T8453 = T8251[1'h0:1'h0];
  assign T8454 = T8455 ? counts_107 : counts_106;
  assign T8455 = T8251[1'h0:1'h0];
  assign T8456 = T8251[1'h1:1'h1];
  assign T8457 = T8462 ? T8460 : T8458;
  assign T8458 = T8459 ? counts_109 : counts_108;
  assign T8459 = T8251[1'h0:1'h0];
  assign T8460 = T8461 ? counts_111 : counts_110;
  assign T8461 = T8251[1'h0:1'h0];
  assign T8462 = T8251[1'h1:1'h1];
  assign T8463 = T8251[2'h2:2'h2];
  assign T8464 = T8251[2'h3:2'h3];
  assign T8465 = T8494 ? T8480 : T8466;
  assign T8466 = T8479 ? T8473 : T8467;
  assign T8467 = T8472 ? T8470 : T8468;
  assign T8468 = T8469 ? counts_113 : counts_112;
  assign T8469 = T8251[1'h0:1'h0];
  assign T8470 = T8471 ? counts_115 : counts_114;
  assign T8471 = T8251[1'h0:1'h0];
  assign T8472 = T8251[1'h1:1'h1];
  assign T8473 = T8478 ? T8476 : T8474;
  assign T8474 = T8475 ? counts_117 : counts_116;
  assign T8475 = T8251[1'h0:1'h0];
  assign T8476 = T8477 ? counts_119 : counts_118;
  assign T8477 = T8251[1'h0:1'h0];
  assign T8478 = T8251[1'h1:1'h1];
  assign T8479 = T8251[2'h2:2'h2];
  assign T8480 = T8493 ? T8487 : T8481;
  assign T8481 = T8486 ? T8484 : T8482;
  assign T8482 = T8483 ? counts_121 : counts_120;
  assign T8483 = T8251[1'h0:1'h0];
  assign T8484 = T8485 ? counts_123 : counts_122;
  assign T8485 = T8251[1'h0:1'h0];
  assign T8486 = T8251[1'h1:1'h1];
  assign T8487 = T8492 ? T8490 : T8488;
  assign T8488 = T8489 ? counts_125 : counts_124;
  assign T8489 = T8251[1'h0:1'h0];
  assign T8490 = T8491 ? counts_127 : counts_126;
  assign T8491 = T8251[1'h0:1'h0];
  assign T8492 = T8251[1'h1:1'h1];
  assign T8493 = T8251[2'h2:2'h2];
  assign T8494 = T8251[2'h3:2'h3];
  assign T8495 = T8251[3'h4:3'h4];
  assign T8496 = T8251[3'h5:3'h5];
  assign T8497 = T8251[3'h6:3'h6];
  assign T8498 = T8751 ? T8625 : T8499;
  assign T8499 = T8624 ? T8562 : T8500;
  assign T8500 = T8561 ? T8531 : T8501;
  assign T8501 = T8530 ? T8516 : T8502;
  assign T8502 = T8515 ? T8509 : T8503;
  assign T8503 = T8508 ? T8506 : T8504;
  assign T8504 = T8505 ? counts_129 : counts_128;
  assign T8505 = T8251[1'h0:1'h0];
  assign T8506 = T8507 ? counts_131 : counts_130;
  assign T8507 = T8251[1'h0:1'h0];
  assign T8508 = T8251[1'h1:1'h1];
  assign T8509 = T8514 ? T8512 : T8510;
  assign T8510 = T8511 ? counts_133 : counts_132;
  assign T8511 = T8251[1'h0:1'h0];
  assign T8512 = T8513 ? counts_135 : counts_134;
  assign T8513 = T8251[1'h0:1'h0];
  assign T8514 = T8251[1'h1:1'h1];
  assign T8515 = T8251[2'h2:2'h2];
  assign T8516 = T8529 ? T8523 : T8517;
  assign T8517 = T8522 ? T8520 : T8518;
  assign T8518 = T8519 ? counts_137 : counts_136;
  assign T8519 = T8251[1'h0:1'h0];
  assign T8520 = T8521 ? counts_139 : counts_138;
  assign T8521 = T8251[1'h0:1'h0];
  assign T8522 = T8251[1'h1:1'h1];
  assign T8523 = T8528 ? T8526 : T8524;
  assign T8524 = T8525 ? counts_141 : counts_140;
  assign T8525 = T8251[1'h0:1'h0];
  assign T8526 = T8527 ? counts_143 : counts_142;
  assign T8527 = T8251[1'h0:1'h0];
  assign T8528 = T8251[1'h1:1'h1];
  assign T8529 = T8251[2'h2:2'h2];
  assign T8530 = T8251[2'h3:2'h3];
  assign T8531 = T8560 ? T8546 : T8532;
  assign T8532 = T8545 ? T8539 : T8533;
  assign T8533 = T8538 ? T8536 : T8534;
  assign T8534 = T8535 ? counts_145 : counts_144;
  assign T8535 = T8251[1'h0:1'h0];
  assign T8536 = T8537 ? counts_147 : counts_146;
  assign T8537 = T8251[1'h0:1'h0];
  assign T8538 = T8251[1'h1:1'h1];
  assign T8539 = T8544 ? T8542 : T8540;
  assign T8540 = T8541 ? counts_149 : counts_148;
  assign T8541 = T8251[1'h0:1'h0];
  assign T8542 = T8543 ? counts_151 : counts_150;
  assign T8543 = T8251[1'h0:1'h0];
  assign T8544 = T8251[1'h1:1'h1];
  assign T8545 = T8251[2'h2:2'h2];
  assign T8546 = T8559 ? T8553 : T8547;
  assign T8547 = T8552 ? T8550 : T8548;
  assign T8548 = T8549 ? counts_153 : counts_152;
  assign T8549 = T8251[1'h0:1'h0];
  assign T8550 = T8551 ? counts_155 : counts_154;
  assign T8551 = T8251[1'h0:1'h0];
  assign T8552 = T8251[1'h1:1'h1];
  assign T8553 = T8558 ? T8556 : T8554;
  assign T8554 = T8555 ? counts_157 : counts_156;
  assign T8555 = T8251[1'h0:1'h0];
  assign T8556 = T8557 ? counts_159 : counts_158;
  assign T8557 = T8251[1'h0:1'h0];
  assign T8558 = T8251[1'h1:1'h1];
  assign T8559 = T8251[2'h2:2'h2];
  assign T8560 = T8251[2'h3:2'h3];
  assign T8561 = T8251[3'h4:3'h4];
  assign T8562 = T8623 ? T8593 : T8563;
  assign T8563 = T8592 ? T8578 : T8564;
  assign T8564 = T8577 ? T8571 : T8565;
  assign T8565 = T8570 ? T8568 : T8566;
  assign T8566 = T8567 ? counts_161 : counts_160;
  assign T8567 = T8251[1'h0:1'h0];
  assign T8568 = T8569 ? counts_163 : counts_162;
  assign T8569 = T8251[1'h0:1'h0];
  assign T8570 = T8251[1'h1:1'h1];
  assign T8571 = T8576 ? T8574 : T8572;
  assign T8572 = T8573 ? counts_165 : counts_164;
  assign T8573 = T8251[1'h0:1'h0];
  assign T8574 = T8575 ? counts_167 : counts_166;
  assign T8575 = T8251[1'h0:1'h0];
  assign T8576 = T8251[1'h1:1'h1];
  assign T8577 = T8251[2'h2:2'h2];
  assign T8578 = T8591 ? T8585 : T8579;
  assign T8579 = T8584 ? T8582 : T8580;
  assign T8580 = T8581 ? counts_169 : counts_168;
  assign T8581 = T8251[1'h0:1'h0];
  assign T8582 = T8583 ? counts_171 : counts_170;
  assign T8583 = T8251[1'h0:1'h0];
  assign T8584 = T8251[1'h1:1'h1];
  assign T8585 = T8590 ? T8588 : T8586;
  assign T8586 = T8587 ? counts_173 : counts_172;
  assign T8587 = T8251[1'h0:1'h0];
  assign T8588 = T8589 ? counts_175 : counts_174;
  assign T8589 = T8251[1'h0:1'h0];
  assign T8590 = T8251[1'h1:1'h1];
  assign T8591 = T8251[2'h2:2'h2];
  assign T8592 = T8251[2'h3:2'h3];
  assign T8593 = T8622 ? T8608 : T8594;
  assign T8594 = T8607 ? T8601 : T8595;
  assign T8595 = T8600 ? T8598 : T8596;
  assign T8596 = T8597 ? counts_177 : counts_176;
  assign T8597 = T8251[1'h0:1'h0];
  assign T8598 = T8599 ? counts_179 : counts_178;
  assign T8599 = T8251[1'h0:1'h0];
  assign T8600 = T8251[1'h1:1'h1];
  assign T8601 = T8606 ? T8604 : T8602;
  assign T8602 = T8603 ? counts_181 : counts_180;
  assign T8603 = T8251[1'h0:1'h0];
  assign T8604 = T8605 ? counts_183 : counts_182;
  assign T8605 = T8251[1'h0:1'h0];
  assign T8606 = T8251[1'h1:1'h1];
  assign T8607 = T8251[2'h2:2'h2];
  assign T8608 = T8621 ? T8615 : T8609;
  assign T8609 = T8614 ? T8612 : T8610;
  assign T8610 = T8611 ? counts_185 : counts_184;
  assign T8611 = T8251[1'h0:1'h0];
  assign T8612 = T8613 ? counts_187 : counts_186;
  assign T8613 = T8251[1'h0:1'h0];
  assign T8614 = T8251[1'h1:1'h1];
  assign T8615 = T8620 ? T8618 : T8616;
  assign T8616 = T8617 ? counts_189 : counts_188;
  assign T8617 = T8251[1'h0:1'h0];
  assign T8618 = T8619 ? counts_191 : counts_190;
  assign T8619 = T8251[1'h0:1'h0];
  assign T8620 = T8251[1'h1:1'h1];
  assign T8621 = T8251[2'h2:2'h2];
  assign T8622 = T8251[2'h3:2'h3];
  assign T8623 = T8251[3'h4:3'h4];
  assign T8624 = T8251[3'h5:3'h5];
  assign T8625 = T8750 ? T8688 : T8626;
  assign T8626 = T8687 ? T8657 : T8627;
  assign T8627 = T8656 ? T8642 : T8628;
  assign T8628 = T8641 ? T8635 : T8629;
  assign T8629 = T8634 ? T8632 : T8630;
  assign T8630 = T8631 ? counts_193 : counts_192;
  assign T8631 = T8251[1'h0:1'h0];
  assign T8632 = T8633 ? counts_195 : counts_194;
  assign T8633 = T8251[1'h0:1'h0];
  assign T8634 = T8251[1'h1:1'h1];
  assign T8635 = T8640 ? T8638 : T8636;
  assign T8636 = T8637 ? counts_197 : counts_196;
  assign T8637 = T8251[1'h0:1'h0];
  assign T8638 = T8639 ? counts_199 : counts_198;
  assign T8639 = T8251[1'h0:1'h0];
  assign T8640 = T8251[1'h1:1'h1];
  assign T8641 = T8251[2'h2:2'h2];
  assign T8642 = T8655 ? T8649 : T8643;
  assign T8643 = T8648 ? T8646 : T8644;
  assign T8644 = T8645 ? counts_201 : counts_200;
  assign T8645 = T8251[1'h0:1'h0];
  assign T8646 = T8647 ? counts_203 : counts_202;
  assign T8647 = T8251[1'h0:1'h0];
  assign T8648 = T8251[1'h1:1'h1];
  assign T8649 = T8654 ? T8652 : T8650;
  assign T8650 = T8651 ? counts_205 : counts_204;
  assign T8651 = T8251[1'h0:1'h0];
  assign T8652 = T8653 ? counts_207 : counts_206;
  assign T8653 = T8251[1'h0:1'h0];
  assign T8654 = T8251[1'h1:1'h1];
  assign T8655 = T8251[2'h2:2'h2];
  assign T8656 = T8251[2'h3:2'h3];
  assign T8657 = T8686 ? T8672 : T8658;
  assign T8658 = T8671 ? T8665 : T8659;
  assign T8659 = T8664 ? T8662 : T8660;
  assign T8660 = T8661 ? counts_209 : counts_208;
  assign T8661 = T8251[1'h0:1'h0];
  assign T8662 = T8663 ? counts_211 : counts_210;
  assign T8663 = T8251[1'h0:1'h0];
  assign T8664 = T8251[1'h1:1'h1];
  assign T8665 = T8670 ? T8668 : T8666;
  assign T8666 = T8667 ? counts_213 : counts_212;
  assign T8667 = T8251[1'h0:1'h0];
  assign T8668 = T8669 ? counts_215 : counts_214;
  assign T8669 = T8251[1'h0:1'h0];
  assign T8670 = T8251[1'h1:1'h1];
  assign T8671 = T8251[2'h2:2'h2];
  assign T8672 = T8685 ? T8679 : T8673;
  assign T8673 = T8678 ? T8676 : T8674;
  assign T8674 = T8675 ? counts_217 : counts_216;
  assign T8675 = T8251[1'h0:1'h0];
  assign T8676 = T8677 ? counts_219 : counts_218;
  assign T8677 = T8251[1'h0:1'h0];
  assign T8678 = T8251[1'h1:1'h1];
  assign T8679 = T8684 ? T8682 : T8680;
  assign T8680 = T8681 ? counts_221 : counts_220;
  assign T8681 = T8251[1'h0:1'h0];
  assign T8682 = T8683 ? counts_223 : counts_222;
  assign T8683 = T8251[1'h0:1'h0];
  assign T8684 = T8251[1'h1:1'h1];
  assign T8685 = T8251[2'h2:2'h2];
  assign T8686 = T8251[2'h3:2'h3];
  assign T8687 = T8251[3'h4:3'h4];
  assign T8688 = T8749 ? T8719 : T8689;
  assign T8689 = T8718 ? T8704 : T8690;
  assign T8690 = T8703 ? T8697 : T8691;
  assign T8691 = T8696 ? T8694 : T8692;
  assign T8692 = T8693 ? counts_225 : counts_224;
  assign T8693 = T8251[1'h0:1'h0];
  assign T8694 = T8695 ? counts_227 : counts_226;
  assign T8695 = T8251[1'h0:1'h0];
  assign T8696 = T8251[1'h1:1'h1];
  assign T8697 = T8702 ? T8700 : T8698;
  assign T8698 = T8699 ? counts_229 : counts_228;
  assign T8699 = T8251[1'h0:1'h0];
  assign T8700 = T8701 ? counts_231 : counts_230;
  assign T8701 = T8251[1'h0:1'h0];
  assign T8702 = T8251[1'h1:1'h1];
  assign T8703 = T8251[2'h2:2'h2];
  assign T8704 = T8717 ? T8711 : T8705;
  assign T8705 = T8710 ? T8708 : T8706;
  assign T8706 = T8707 ? counts_233 : counts_232;
  assign T8707 = T8251[1'h0:1'h0];
  assign T8708 = T8709 ? counts_235 : counts_234;
  assign T8709 = T8251[1'h0:1'h0];
  assign T8710 = T8251[1'h1:1'h1];
  assign T8711 = T8716 ? T8714 : T8712;
  assign T8712 = T8713 ? counts_237 : counts_236;
  assign T8713 = T8251[1'h0:1'h0];
  assign T8714 = T8715 ? counts_239 : counts_238;
  assign T8715 = T8251[1'h0:1'h0];
  assign T8716 = T8251[1'h1:1'h1];
  assign T8717 = T8251[2'h2:2'h2];
  assign T8718 = T8251[2'h3:2'h3];
  assign T8719 = T8748 ? T8734 : T8720;
  assign T8720 = T8733 ? T8727 : T8721;
  assign T8721 = T8726 ? T8724 : T8722;
  assign T8722 = T8723 ? counts_241 : counts_240;
  assign T8723 = T8251[1'h0:1'h0];
  assign T8724 = T8725 ? counts_243 : counts_242;
  assign T8725 = T8251[1'h0:1'h0];
  assign T8726 = T8251[1'h1:1'h1];
  assign T8727 = T8732 ? T8730 : T8728;
  assign T8728 = T8729 ? counts_245 : counts_244;
  assign T8729 = T8251[1'h0:1'h0];
  assign T8730 = T8731 ? counts_247 : counts_246;
  assign T8731 = T8251[1'h0:1'h0];
  assign T8732 = T8251[1'h1:1'h1];
  assign T8733 = T8251[2'h2:2'h2];
  assign T8734 = T8747 ? T8741 : T8735;
  assign T8735 = T8740 ? T8738 : T8736;
  assign T8736 = T8737 ? counts_249 : counts_248;
  assign T8737 = T8251[1'h0:1'h0];
  assign T8738 = T8739 ? counts_251 : counts_250;
  assign T8739 = T8251[1'h0:1'h0];
  assign T8740 = T8251[1'h1:1'h1];
  assign T8741 = T8746 ? T8744 : T8742;
  assign T8742 = T8743 ? counts_253 : counts_252;
  assign T8743 = T8251[1'h0:1'h0];
  assign T8744 = T8745 ? counts_255 : counts_254;
  assign T8745 = T8251[1'h0:1'h0];
  assign T8746 = T8251[1'h1:1'h1];
  assign T8747 = T8251[2'h2:2'h2];
  assign T8748 = T8251[2'h3:2'h3];
  assign T8749 = T8251[3'h4:3'h4];
  assign T8750 = T8251[3'h5:3'h5];
  assign T8751 = T8251[3'h6:3'h6];
  assign T8752 = T8251[3'h7:3'h7];
  assign T8753 = T9262 ? T9008 : T8754;
  assign T8754 = T9007 ? T8881 : T8755;
  assign T8755 = T8880 ? T8818 : T8756;
  assign T8756 = T8817 ? T8787 : T8757;
  assign T8757 = T8786 ? T8772 : T8758;
  assign T8758 = T8771 ? T8765 : T8759;
  assign T8759 = T8764 ? T8762 : T8760;
  assign T8760 = T8761 ? counts_257 : counts_256;
  assign T8761 = T8251[1'h0:1'h0];
  assign T8762 = T8763 ? counts_259 : counts_258;
  assign T8763 = T8251[1'h0:1'h0];
  assign T8764 = T8251[1'h1:1'h1];
  assign T8765 = T8770 ? T8768 : T8766;
  assign T8766 = T8767 ? counts_261 : counts_260;
  assign T8767 = T8251[1'h0:1'h0];
  assign T8768 = T8769 ? counts_263 : counts_262;
  assign T8769 = T8251[1'h0:1'h0];
  assign T8770 = T8251[1'h1:1'h1];
  assign T8771 = T8251[2'h2:2'h2];
  assign T8772 = T8785 ? T8779 : T8773;
  assign T8773 = T8778 ? T8776 : T8774;
  assign T8774 = T8775 ? counts_265 : counts_264;
  assign T8775 = T8251[1'h0:1'h0];
  assign T8776 = T8777 ? counts_267 : counts_266;
  assign T8777 = T8251[1'h0:1'h0];
  assign T8778 = T8251[1'h1:1'h1];
  assign T8779 = T8784 ? T8782 : T8780;
  assign T8780 = T8781 ? counts_269 : counts_268;
  assign T8781 = T8251[1'h0:1'h0];
  assign T8782 = T8783 ? counts_271 : counts_270;
  assign T8783 = T8251[1'h0:1'h0];
  assign T8784 = T8251[1'h1:1'h1];
  assign T8785 = T8251[2'h2:2'h2];
  assign T8786 = T8251[2'h3:2'h3];
  assign T8787 = T8816 ? T8802 : T8788;
  assign T8788 = T8801 ? T8795 : T8789;
  assign T8789 = T8794 ? T8792 : T8790;
  assign T8790 = T8791 ? counts_273 : counts_272;
  assign T8791 = T8251[1'h0:1'h0];
  assign T8792 = T8793 ? counts_275 : counts_274;
  assign T8793 = T8251[1'h0:1'h0];
  assign T8794 = T8251[1'h1:1'h1];
  assign T8795 = T8800 ? T8798 : T8796;
  assign T8796 = T8797 ? counts_277 : counts_276;
  assign T8797 = T8251[1'h0:1'h0];
  assign T8798 = T8799 ? counts_279 : counts_278;
  assign T8799 = T8251[1'h0:1'h0];
  assign T8800 = T8251[1'h1:1'h1];
  assign T8801 = T8251[2'h2:2'h2];
  assign T8802 = T8815 ? T8809 : T8803;
  assign T8803 = T8808 ? T8806 : T8804;
  assign T8804 = T8805 ? counts_281 : counts_280;
  assign T8805 = T8251[1'h0:1'h0];
  assign T8806 = T8807 ? counts_283 : counts_282;
  assign T8807 = T8251[1'h0:1'h0];
  assign T8808 = T8251[1'h1:1'h1];
  assign T8809 = T8814 ? T8812 : T8810;
  assign T8810 = T8811 ? counts_285 : counts_284;
  assign T8811 = T8251[1'h0:1'h0];
  assign T8812 = T8813 ? counts_287 : counts_286;
  assign T8813 = T8251[1'h0:1'h0];
  assign T8814 = T8251[1'h1:1'h1];
  assign T8815 = T8251[2'h2:2'h2];
  assign T8816 = T8251[2'h3:2'h3];
  assign T8817 = T8251[3'h4:3'h4];
  assign T8818 = T8879 ? T8849 : T8819;
  assign T8819 = T8848 ? T8834 : T8820;
  assign T8820 = T8833 ? T8827 : T8821;
  assign T8821 = T8826 ? T8824 : T8822;
  assign T8822 = T8823 ? counts_289 : counts_288;
  assign T8823 = T8251[1'h0:1'h0];
  assign T8824 = T8825 ? counts_291 : counts_290;
  assign T8825 = T8251[1'h0:1'h0];
  assign T8826 = T8251[1'h1:1'h1];
  assign T8827 = T8832 ? T8830 : T8828;
  assign T8828 = T8829 ? counts_293 : counts_292;
  assign T8829 = T8251[1'h0:1'h0];
  assign T8830 = T8831 ? counts_295 : counts_294;
  assign T8831 = T8251[1'h0:1'h0];
  assign T8832 = T8251[1'h1:1'h1];
  assign T8833 = T8251[2'h2:2'h2];
  assign T8834 = T8847 ? T8841 : T8835;
  assign T8835 = T8840 ? T8838 : T8836;
  assign T8836 = T8837 ? counts_297 : counts_296;
  assign T8837 = T8251[1'h0:1'h0];
  assign T8838 = T8839 ? counts_299 : counts_298;
  assign T8839 = T8251[1'h0:1'h0];
  assign T8840 = T8251[1'h1:1'h1];
  assign T8841 = T8846 ? T8844 : T8842;
  assign T8842 = T8843 ? counts_301 : counts_300;
  assign T8843 = T8251[1'h0:1'h0];
  assign T8844 = T8845 ? counts_303 : counts_302;
  assign T8845 = T8251[1'h0:1'h0];
  assign T8846 = T8251[1'h1:1'h1];
  assign T8847 = T8251[2'h2:2'h2];
  assign T8848 = T8251[2'h3:2'h3];
  assign T8849 = T8878 ? T8864 : T8850;
  assign T8850 = T8863 ? T8857 : T8851;
  assign T8851 = T8856 ? T8854 : T8852;
  assign T8852 = T8853 ? counts_305 : counts_304;
  assign T8853 = T8251[1'h0:1'h0];
  assign T8854 = T8855 ? counts_307 : counts_306;
  assign T8855 = T8251[1'h0:1'h0];
  assign T8856 = T8251[1'h1:1'h1];
  assign T8857 = T8862 ? T8860 : T8858;
  assign T8858 = T8859 ? counts_309 : counts_308;
  assign T8859 = T8251[1'h0:1'h0];
  assign T8860 = T8861 ? counts_311 : counts_310;
  assign T8861 = T8251[1'h0:1'h0];
  assign T8862 = T8251[1'h1:1'h1];
  assign T8863 = T8251[2'h2:2'h2];
  assign T8864 = T8877 ? T8871 : T8865;
  assign T8865 = T8870 ? T8868 : T8866;
  assign T8866 = T8867 ? counts_313 : counts_312;
  assign T8867 = T8251[1'h0:1'h0];
  assign T8868 = T8869 ? counts_315 : counts_314;
  assign T8869 = T8251[1'h0:1'h0];
  assign T8870 = T8251[1'h1:1'h1];
  assign T8871 = T8876 ? T8874 : T8872;
  assign T8872 = T8873 ? counts_317 : counts_316;
  assign T8873 = T8251[1'h0:1'h0];
  assign T8874 = T8875 ? counts_319 : counts_318;
  assign T8875 = T8251[1'h0:1'h0];
  assign T8876 = T8251[1'h1:1'h1];
  assign T8877 = T8251[2'h2:2'h2];
  assign T8878 = T8251[2'h3:2'h3];
  assign T8879 = T8251[3'h4:3'h4];
  assign T8880 = T8251[3'h5:3'h5];
  assign T8881 = T9006 ? T8944 : T8882;
  assign T8882 = T8943 ? T8913 : T8883;
  assign T8883 = T8912 ? T8898 : T8884;
  assign T8884 = T8897 ? T8891 : T8885;
  assign T8885 = T8890 ? T8888 : T8886;
  assign T8886 = T8887 ? counts_321 : counts_320;
  assign T8887 = T8251[1'h0:1'h0];
  assign T8888 = T8889 ? counts_323 : counts_322;
  assign T8889 = T8251[1'h0:1'h0];
  assign T8890 = T8251[1'h1:1'h1];
  assign T8891 = T8896 ? T8894 : T8892;
  assign T8892 = T8893 ? counts_325 : counts_324;
  assign T8893 = T8251[1'h0:1'h0];
  assign T8894 = T8895 ? counts_327 : counts_326;
  assign T8895 = T8251[1'h0:1'h0];
  assign T8896 = T8251[1'h1:1'h1];
  assign T8897 = T8251[2'h2:2'h2];
  assign T8898 = T8911 ? T8905 : T8899;
  assign T8899 = T8904 ? T8902 : T8900;
  assign T8900 = T8901 ? counts_329 : counts_328;
  assign T8901 = T8251[1'h0:1'h0];
  assign T8902 = T8903 ? counts_331 : counts_330;
  assign T8903 = T8251[1'h0:1'h0];
  assign T8904 = T8251[1'h1:1'h1];
  assign T8905 = T8910 ? T8908 : T8906;
  assign T8906 = T8907 ? counts_333 : counts_332;
  assign T8907 = T8251[1'h0:1'h0];
  assign T8908 = T8909 ? counts_335 : counts_334;
  assign T8909 = T8251[1'h0:1'h0];
  assign T8910 = T8251[1'h1:1'h1];
  assign T8911 = T8251[2'h2:2'h2];
  assign T8912 = T8251[2'h3:2'h3];
  assign T8913 = T8942 ? T8928 : T8914;
  assign T8914 = T8927 ? T8921 : T8915;
  assign T8915 = T8920 ? T8918 : T8916;
  assign T8916 = T8917 ? counts_337 : counts_336;
  assign T8917 = T8251[1'h0:1'h0];
  assign T8918 = T8919 ? counts_339 : counts_338;
  assign T8919 = T8251[1'h0:1'h0];
  assign T8920 = T8251[1'h1:1'h1];
  assign T8921 = T8926 ? T8924 : T8922;
  assign T8922 = T8923 ? counts_341 : counts_340;
  assign T8923 = T8251[1'h0:1'h0];
  assign T8924 = T8925 ? counts_343 : counts_342;
  assign T8925 = T8251[1'h0:1'h0];
  assign T8926 = T8251[1'h1:1'h1];
  assign T8927 = T8251[2'h2:2'h2];
  assign T8928 = T8941 ? T8935 : T8929;
  assign T8929 = T8934 ? T8932 : T8930;
  assign T8930 = T8931 ? counts_345 : counts_344;
  assign T8931 = T8251[1'h0:1'h0];
  assign T8932 = T8933 ? counts_347 : counts_346;
  assign T8933 = T8251[1'h0:1'h0];
  assign T8934 = T8251[1'h1:1'h1];
  assign T8935 = T8940 ? T8938 : T8936;
  assign T8936 = T8937 ? counts_349 : counts_348;
  assign T8937 = T8251[1'h0:1'h0];
  assign T8938 = T8939 ? counts_351 : counts_350;
  assign T8939 = T8251[1'h0:1'h0];
  assign T8940 = T8251[1'h1:1'h1];
  assign T8941 = T8251[2'h2:2'h2];
  assign T8942 = T8251[2'h3:2'h3];
  assign T8943 = T8251[3'h4:3'h4];
  assign T8944 = T9005 ? T8975 : T8945;
  assign T8945 = T8974 ? T8960 : T8946;
  assign T8946 = T8959 ? T8953 : T8947;
  assign T8947 = T8952 ? T8950 : T8948;
  assign T8948 = T8949 ? counts_353 : counts_352;
  assign T8949 = T8251[1'h0:1'h0];
  assign T8950 = T8951 ? counts_355 : counts_354;
  assign T8951 = T8251[1'h0:1'h0];
  assign T8952 = T8251[1'h1:1'h1];
  assign T8953 = T8958 ? T8956 : T8954;
  assign T8954 = T8955 ? counts_357 : counts_356;
  assign T8955 = T8251[1'h0:1'h0];
  assign T8956 = T8957 ? counts_359 : counts_358;
  assign T8957 = T8251[1'h0:1'h0];
  assign T8958 = T8251[1'h1:1'h1];
  assign T8959 = T8251[2'h2:2'h2];
  assign T8960 = T8973 ? T8967 : T8961;
  assign T8961 = T8966 ? T8964 : T8962;
  assign T8962 = T8963 ? counts_361 : counts_360;
  assign T8963 = T8251[1'h0:1'h0];
  assign T8964 = T8965 ? counts_363 : counts_362;
  assign T8965 = T8251[1'h0:1'h0];
  assign T8966 = T8251[1'h1:1'h1];
  assign T8967 = T8972 ? T8970 : T8968;
  assign T8968 = T8969 ? counts_365 : counts_364;
  assign T8969 = T8251[1'h0:1'h0];
  assign T8970 = T8971 ? counts_367 : counts_366;
  assign T8971 = T8251[1'h0:1'h0];
  assign T8972 = T8251[1'h1:1'h1];
  assign T8973 = T8251[2'h2:2'h2];
  assign T8974 = T8251[2'h3:2'h3];
  assign T8975 = T9004 ? T8990 : T8976;
  assign T8976 = T8989 ? T8983 : T8977;
  assign T8977 = T8982 ? T8980 : T8978;
  assign T8978 = T8979 ? counts_369 : counts_368;
  assign T8979 = T8251[1'h0:1'h0];
  assign T8980 = T8981 ? counts_371 : counts_370;
  assign T8981 = T8251[1'h0:1'h0];
  assign T8982 = T8251[1'h1:1'h1];
  assign T8983 = T8988 ? T8986 : T8984;
  assign T8984 = T8985 ? counts_373 : counts_372;
  assign T8985 = T8251[1'h0:1'h0];
  assign T8986 = T8987 ? counts_375 : counts_374;
  assign T8987 = T8251[1'h0:1'h0];
  assign T8988 = T8251[1'h1:1'h1];
  assign T8989 = T8251[2'h2:2'h2];
  assign T8990 = T9003 ? T8997 : T8991;
  assign T8991 = T8996 ? T8994 : T8992;
  assign T8992 = T8993 ? counts_377 : counts_376;
  assign T8993 = T8251[1'h0:1'h0];
  assign T8994 = T8995 ? counts_379 : counts_378;
  assign T8995 = T8251[1'h0:1'h0];
  assign T8996 = T8251[1'h1:1'h1];
  assign T8997 = T9002 ? T9000 : T8998;
  assign T8998 = T8999 ? counts_381 : counts_380;
  assign T8999 = T8251[1'h0:1'h0];
  assign T9000 = T9001 ? counts_383 : counts_382;
  assign T9001 = T8251[1'h0:1'h0];
  assign T9002 = T8251[1'h1:1'h1];
  assign T9003 = T8251[2'h2:2'h2];
  assign T9004 = T8251[2'h3:2'h3];
  assign T9005 = T8251[3'h4:3'h4];
  assign T9006 = T8251[3'h5:3'h5];
  assign T9007 = T8251[3'h6:3'h6];
  assign T9008 = T9261 ? T9135 : T9009;
  assign T9009 = T9134 ? T9072 : T9010;
  assign T9010 = T9071 ? T9041 : T9011;
  assign T9011 = T9040 ? T9026 : T9012;
  assign T9012 = T9025 ? T9019 : T9013;
  assign T9013 = T9018 ? T9016 : T9014;
  assign T9014 = T9015 ? counts_385 : counts_384;
  assign T9015 = T8251[1'h0:1'h0];
  assign T9016 = T9017 ? counts_387 : counts_386;
  assign T9017 = T8251[1'h0:1'h0];
  assign T9018 = T8251[1'h1:1'h1];
  assign T9019 = T9024 ? T9022 : T9020;
  assign T9020 = T9021 ? counts_389 : counts_388;
  assign T9021 = T8251[1'h0:1'h0];
  assign T9022 = T9023 ? counts_391 : counts_390;
  assign T9023 = T8251[1'h0:1'h0];
  assign T9024 = T8251[1'h1:1'h1];
  assign T9025 = T8251[2'h2:2'h2];
  assign T9026 = T9039 ? T9033 : T9027;
  assign T9027 = T9032 ? T9030 : T9028;
  assign T9028 = T9029 ? counts_393 : counts_392;
  assign T9029 = T8251[1'h0:1'h0];
  assign T9030 = T9031 ? counts_395 : counts_394;
  assign T9031 = T8251[1'h0:1'h0];
  assign T9032 = T8251[1'h1:1'h1];
  assign T9033 = T9038 ? T9036 : T9034;
  assign T9034 = T9035 ? counts_397 : counts_396;
  assign T9035 = T8251[1'h0:1'h0];
  assign T9036 = T9037 ? counts_399 : counts_398;
  assign T9037 = T8251[1'h0:1'h0];
  assign T9038 = T8251[1'h1:1'h1];
  assign T9039 = T8251[2'h2:2'h2];
  assign T9040 = T8251[2'h3:2'h3];
  assign T9041 = T9070 ? T9056 : T9042;
  assign T9042 = T9055 ? T9049 : T9043;
  assign T9043 = T9048 ? T9046 : T9044;
  assign T9044 = T9045 ? counts_401 : counts_400;
  assign T9045 = T8251[1'h0:1'h0];
  assign T9046 = T9047 ? counts_403 : counts_402;
  assign T9047 = T8251[1'h0:1'h0];
  assign T9048 = T8251[1'h1:1'h1];
  assign T9049 = T9054 ? T9052 : T9050;
  assign T9050 = T9051 ? counts_405 : counts_404;
  assign T9051 = T8251[1'h0:1'h0];
  assign T9052 = T9053 ? counts_407 : counts_406;
  assign T9053 = T8251[1'h0:1'h0];
  assign T9054 = T8251[1'h1:1'h1];
  assign T9055 = T8251[2'h2:2'h2];
  assign T9056 = T9069 ? T9063 : T9057;
  assign T9057 = T9062 ? T9060 : T9058;
  assign T9058 = T9059 ? counts_409 : counts_408;
  assign T9059 = T8251[1'h0:1'h0];
  assign T9060 = T9061 ? counts_411 : counts_410;
  assign T9061 = T8251[1'h0:1'h0];
  assign T9062 = T8251[1'h1:1'h1];
  assign T9063 = T9068 ? T9066 : T9064;
  assign T9064 = T9065 ? counts_413 : counts_412;
  assign T9065 = T8251[1'h0:1'h0];
  assign T9066 = T9067 ? counts_415 : counts_414;
  assign T9067 = T8251[1'h0:1'h0];
  assign T9068 = T8251[1'h1:1'h1];
  assign T9069 = T8251[2'h2:2'h2];
  assign T9070 = T8251[2'h3:2'h3];
  assign T9071 = T8251[3'h4:3'h4];
  assign T9072 = T9133 ? T9103 : T9073;
  assign T9073 = T9102 ? T9088 : T9074;
  assign T9074 = T9087 ? T9081 : T9075;
  assign T9075 = T9080 ? T9078 : T9076;
  assign T9076 = T9077 ? counts_417 : counts_416;
  assign T9077 = T8251[1'h0:1'h0];
  assign T9078 = T9079 ? counts_419 : counts_418;
  assign T9079 = T8251[1'h0:1'h0];
  assign T9080 = T8251[1'h1:1'h1];
  assign T9081 = T9086 ? T9084 : T9082;
  assign T9082 = T9083 ? counts_421 : counts_420;
  assign T9083 = T8251[1'h0:1'h0];
  assign T9084 = T9085 ? counts_423 : counts_422;
  assign T9085 = T8251[1'h0:1'h0];
  assign T9086 = T8251[1'h1:1'h1];
  assign T9087 = T8251[2'h2:2'h2];
  assign T9088 = T9101 ? T9095 : T9089;
  assign T9089 = T9094 ? T9092 : T9090;
  assign T9090 = T9091 ? counts_425 : counts_424;
  assign T9091 = T8251[1'h0:1'h0];
  assign T9092 = T9093 ? counts_427 : counts_426;
  assign T9093 = T8251[1'h0:1'h0];
  assign T9094 = T8251[1'h1:1'h1];
  assign T9095 = T9100 ? T9098 : T9096;
  assign T9096 = T9097 ? counts_429 : counts_428;
  assign T9097 = T8251[1'h0:1'h0];
  assign T9098 = T9099 ? counts_431 : counts_430;
  assign T9099 = T8251[1'h0:1'h0];
  assign T9100 = T8251[1'h1:1'h1];
  assign T9101 = T8251[2'h2:2'h2];
  assign T9102 = T8251[2'h3:2'h3];
  assign T9103 = T9132 ? T9118 : T9104;
  assign T9104 = T9117 ? T9111 : T9105;
  assign T9105 = T9110 ? T9108 : T9106;
  assign T9106 = T9107 ? counts_433 : counts_432;
  assign T9107 = T8251[1'h0:1'h0];
  assign T9108 = T9109 ? counts_435 : counts_434;
  assign T9109 = T8251[1'h0:1'h0];
  assign T9110 = T8251[1'h1:1'h1];
  assign T9111 = T9116 ? T9114 : T9112;
  assign T9112 = T9113 ? counts_437 : counts_436;
  assign T9113 = T8251[1'h0:1'h0];
  assign T9114 = T9115 ? counts_439 : counts_438;
  assign T9115 = T8251[1'h0:1'h0];
  assign T9116 = T8251[1'h1:1'h1];
  assign T9117 = T8251[2'h2:2'h2];
  assign T9118 = T9131 ? T9125 : T9119;
  assign T9119 = T9124 ? T9122 : T9120;
  assign T9120 = T9121 ? counts_441 : counts_440;
  assign T9121 = T8251[1'h0:1'h0];
  assign T9122 = T9123 ? counts_443 : counts_442;
  assign T9123 = T8251[1'h0:1'h0];
  assign T9124 = T8251[1'h1:1'h1];
  assign T9125 = T9130 ? T9128 : T9126;
  assign T9126 = T9127 ? counts_445 : counts_444;
  assign T9127 = T8251[1'h0:1'h0];
  assign T9128 = T9129 ? counts_447 : counts_446;
  assign T9129 = T8251[1'h0:1'h0];
  assign T9130 = T8251[1'h1:1'h1];
  assign T9131 = T8251[2'h2:2'h2];
  assign T9132 = T8251[2'h3:2'h3];
  assign T9133 = T8251[3'h4:3'h4];
  assign T9134 = T8251[3'h5:3'h5];
  assign T9135 = T9260 ? T9198 : T9136;
  assign T9136 = T9197 ? T9167 : T9137;
  assign T9137 = T9166 ? T9152 : T9138;
  assign T9138 = T9151 ? T9145 : T9139;
  assign T9139 = T9144 ? T9142 : T9140;
  assign T9140 = T9141 ? counts_449 : counts_448;
  assign T9141 = T8251[1'h0:1'h0];
  assign T9142 = T9143 ? counts_451 : counts_450;
  assign T9143 = T8251[1'h0:1'h0];
  assign T9144 = T8251[1'h1:1'h1];
  assign T9145 = T9150 ? T9148 : T9146;
  assign T9146 = T9147 ? counts_453 : counts_452;
  assign T9147 = T8251[1'h0:1'h0];
  assign T9148 = T9149 ? counts_455 : counts_454;
  assign T9149 = T8251[1'h0:1'h0];
  assign T9150 = T8251[1'h1:1'h1];
  assign T9151 = T8251[2'h2:2'h2];
  assign T9152 = T9165 ? T9159 : T9153;
  assign T9153 = T9158 ? T9156 : T9154;
  assign T9154 = T9155 ? counts_457 : counts_456;
  assign T9155 = T8251[1'h0:1'h0];
  assign T9156 = T9157 ? counts_459 : counts_458;
  assign T9157 = T8251[1'h0:1'h0];
  assign T9158 = T8251[1'h1:1'h1];
  assign T9159 = T9164 ? T9162 : T9160;
  assign T9160 = T9161 ? counts_461 : counts_460;
  assign T9161 = T8251[1'h0:1'h0];
  assign T9162 = T9163 ? counts_463 : counts_462;
  assign T9163 = T8251[1'h0:1'h0];
  assign T9164 = T8251[1'h1:1'h1];
  assign T9165 = T8251[2'h2:2'h2];
  assign T9166 = T8251[2'h3:2'h3];
  assign T9167 = T9196 ? T9182 : T9168;
  assign T9168 = T9181 ? T9175 : T9169;
  assign T9169 = T9174 ? T9172 : T9170;
  assign T9170 = T9171 ? counts_465 : counts_464;
  assign T9171 = T8251[1'h0:1'h0];
  assign T9172 = T9173 ? counts_467 : counts_466;
  assign T9173 = T8251[1'h0:1'h0];
  assign T9174 = T8251[1'h1:1'h1];
  assign T9175 = T9180 ? T9178 : T9176;
  assign T9176 = T9177 ? counts_469 : counts_468;
  assign T9177 = T8251[1'h0:1'h0];
  assign T9178 = T9179 ? counts_471 : counts_470;
  assign T9179 = T8251[1'h0:1'h0];
  assign T9180 = T8251[1'h1:1'h1];
  assign T9181 = T8251[2'h2:2'h2];
  assign T9182 = T9195 ? T9189 : T9183;
  assign T9183 = T9188 ? T9186 : T9184;
  assign T9184 = T9185 ? counts_473 : counts_472;
  assign T9185 = T8251[1'h0:1'h0];
  assign T9186 = T9187 ? counts_475 : counts_474;
  assign T9187 = T8251[1'h0:1'h0];
  assign T9188 = T8251[1'h1:1'h1];
  assign T9189 = T9194 ? T9192 : T9190;
  assign T9190 = T9191 ? counts_477 : counts_476;
  assign T9191 = T8251[1'h0:1'h0];
  assign T9192 = T9193 ? counts_479 : counts_478;
  assign T9193 = T8251[1'h0:1'h0];
  assign T9194 = T8251[1'h1:1'h1];
  assign T9195 = T8251[2'h2:2'h2];
  assign T9196 = T8251[2'h3:2'h3];
  assign T9197 = T8251[3'h4:3'h4];
  assign T9198 = T9259 ? T9229 : T9199;
  assign T9199 = T9228 ? T9214 : T9200;
  assign T9200 = T9213 ? T9207 : T9201;
  assign T9201 = T9206 ? T9204 : T9202;
  assign T9202 = T9203 ? counts_481 : counts_480;
  assign T9203 = T8251[1'h0:1'h0];
  assign T9204 = T9205 ? counts_483 : counts_482;
  assign T9205 = T8251[1'h0:1'h0];
  assign T9206 = T8251[1'h1:1'h1];
  assign T9207 = T9212 ? T9210 : T9208;
  assign T9208 = T9209 ? counts_485 : counts_484;
  assign T9209 = T8251[1'h0:1'h0];
  assign T9210 = T9211 ? counts_487 : counts_486;
  assign T9211 = T8251[1'h0:1'h0];
  assign T9212 = T8251[1'h1:1'h1];
  assign T9213 = T8251[2'h2:2'h2];
  assign T9214 = T9227 ? T9221 : T9215;
  assign T9215 = T9220 ? T9218 : T9216;
  assign T9216 = T9217 ? counts_489 : counts_488;
  assign T9217 = T8251[1'h0:1'h0];
  assign T9218 = T9219 ? counts_491 : counts_490;
  assign T9219 = T8251[1'h0:1'h0];
  assign T9220 = T8251[1'h1:1'h1];
  assign T9221 = T9226 ? T9224 : T9222;
  assign T9222 = T9223 ? counts_493 : counts_492;
  assign T9223 = T8251[1'h0:1'h0];
  assign T9224 = T9225 ? counts_495 : counts_494;
  assign T9225 = T8251[1'h0:1'h0];
  assign T9226 = T8251[1'h1:1'h1];
  assign T9227 = T8251[2'h2:2'h2];
  assign T9228 = T8251[2'h3:2'h3];
  assign T9229 = T9258 ? T9244 : T9230;
  assign T9230 = T9243 ? T9237 : T9231;
  assign T9231 = T9236 ? T9234 : T9232;
  assign T9232 = T9233 ? counts_497 : counts_496;
  assign T9233 = T8251[1'h0:1'h0];
  assign T9234 = T9235 ? counts_499 : counts_498;
  assign T9235 = T8251[1'h0:1'h0];
  assign T9236 = T8251[1'h1:1'h1];
  assign T9237 = T9242 ? T9240 : T9238;
  assign T9238 = T9239 ? counts_501 : counts_500;
  assign T9239 = T8251[1'h0:1'h0];
  assign T9240 = T9241 ? counts_503 : counts_502;
  assign T9241 = T8251[1'h0:1'h0];
  assign T9242 = T8251[1'h1:1'h1];
  assign T9243 = T8251[2'h2:2'h2];
  assign T9244 = T9257 ? T9251 : T9245;
  assign T9245 = T9250 ? T9248 : T9246;
  assign T9246 = T9247 ? counts_505 : counts_504;
  assign T9247 = T8251[1'h0:1'h0];
  assign T9248 = T9249 ? counts_507 : counts_506;
  assign T9249 = T8251[1'h0:1'h0];
  assign T9250 = T8251[1'h1:1'h1];
  assign T9251 = T9256 ? T9254 : T9252;
  assign T9252 = T9253 ? counts_509 : counts_508;
  assign T9253 = T8251[1'h0:1'h0];
  assign T9254 = T9255 ? counts_511 : counts_510;
  assign T9255 = T8251[1'h0:1'h0];
  assign T9256 = T8251[1'h1:1'h1];
  assign T9257 = T8251[2'h2:2'h2];
  assign T9258 = T8251[2'h3:2'h3];
  assign T9259 = T8251[3'h4:3'h4];
  assign T9260 = T8251[3'h5:3'h5];
  assign T9261 = T8251[3'h6:3'h6];
  assign T9262 = T8251[3'h7:3'h7];
  assign T9263 = T8251[4'h8:4'h8];
  assign T9264 = T10285 ? T9775 : T9265;
  assign T9265 = T9774 ? T9520 : T9266;
  assign T9266 = T9519 ? T9393 : T9267;
  assign T9267 = T9392 ? T9330 : T9268;
  assign T9268 = T9329 ? T9299 : T9269;
  assign T9269 = T9298 ? T9284 : T9270;
  assign T9270 = T9283 ? T9277 : T9271;
  assign T9271 = T9276 ? T9274 : T9272;
  assign T9272 = T9273 ? counts_513 : counts_512;
  assign T9273 = T8251[1'h0:1'h0];
  assign T9274 = T9275 ? counts_515 : counts_514;
  assign T9275 = T8251[1'h0:1'h0];
  assign T9276 = T8251[1'h1:1'h1];
  assign T9277 = T9282 ? T9280 : T9278;
  assign T9278 = T9279 ? counts_517 : counts_516;
  assign T9279 = T8251[1'h0:1'h0];
  assign T9280 = T9281 ? counts_519 : counts_518;
  assign T9281 = T8251[1'h0:1'h0];
  assign T9282 = T8251[1'h1:1'h1];
  assign T9283 = T8251[2'h2:2'h2];
  assign T9284 = T9297 ? T9291 : T9285;
  assign T9285 = T9290 ? T9288 : T9286;
  assign T9286 = T9287 ? counts_521 : counts_520;
  assign T9287 = T8251[1'h0:1'h0];
  assign T9288 = T9289 ? counts_523 : counts_522;
  assign T9289 = T8251[1'h0:1'h0];
  assign T9290 = T8251[1'h1:1'h1];
  assign T9291 = T9296 ? T9294 : T9292;
  assign T9292 = T9293 ? counts_525 : counts_524;
  assign T9293 = T8251[1'h0:1'h0];
  assign T9294 = T9295 ? counts_527 : counts_526;
  assign T9295 = T8251[1'h0:1'h0];
  assign T9296 = T8251[1'h1:1'h1];
  assign T9297 = T8251[2'h2:2'h2];
  assign T9298 = T8251[2'h3:2'h3];
  assign T9299 = T9328 ? T9314 : T9300;
  assign T9300 = T9313 ? T9307 : T9301;
  assign T9301 = T9306 ? T9304 : T9302;
  assign T9302 = T9303 ? counts_529 : counts_528;
  assign T9303 = T8251[1'h0:1'h0];
  assign T9304 = T9305 ? counts_531 : counts_530;
  assign T9305 = T8251[1'h0:1'h0];
  assign T9306 = T8251[1'h1:1'h1];
  assign T9307 = T9312 ? T9310 : T9308;
  assign T9308 = T9309 ? counts_533 : counts_532;
  assign T9309 = T8251[1'h0:1'h0];
  assign T9310 = T9311 ? counts_535 : counts_534;
  assign T9311 = T8251[1'h0:1'h0];
  assign T9312 = T8251[1'h1:1'h1];
  assign T9313 = T8251[2'h2:2'h2];
  assign T9314 = T9327 ? T9321 : T9315;
  assign T9315 = T9320 ? T9318 : T9316;
  assign T9316 = T9317 ? counts_537 : counts_536;
  assign T9317 = T8251[1'h0:1'h0];
  assign T9318 = T9319 ? counts_539 : counts_538;
  assign T9319 = T8251[1'h0:1'h0];
  assign T9320 = T8251[1'h1:1'h1];
  assign T9321 = T9326 ? T9324 : T9322;
  assign T9322 = T9323 ? counts_541 : counts_540;
  assign T9323 = T8251[1'h0:1'h0];
  assign T9324 = T9325 ? counts_543 : counts_542;
  assign T9325 = T8251[1'h0:1'h0];
  assign T9326 = T8251[1'h1:1'h1];
  assign T9327 = T8251[2'h2:2'h2];
  assign T9328 = T8251[2'h3:2'h3];
  assign T9329 = T8251[3'h4:3'h4];
  assign T9330 = T9391 ? T9361 : T9331;
  assign T9331 = T9360 ? T9346 : T9332;
  assign T9332 = T9345 ? T9339 : T9333;
  assign T9333 = T9338 ? T9336 : T9334;
  assign T9334 = T9335 ? counts_545 : counts_544;
  assign T9335 = T8251[1'h0:1'h0];
  assign T9336 = T9337 ? counts_547 : counts_546;
  assign T9337 = T8251[1'h0:1'h0];
  assign T9338 = T8251[1'h1:1'h1];
  assign T9339 = T9344 ? T9342 : T9340;
  assign T9340 = T9341 ? counts_549 : counts_548;
  assign T9341 = T8251[1'h0:1'h0];
  assign T9342 = T9343 ? counts_551 : counts_550;
  assign T9343 = T8251[1'h0:1'h0];
  assign T9344 = T8251[1'h1:1'h1];
  assign T9345 = T8251[2'h2:2'h2];
  assign T9346 = T9359 ? T9353 : T9347;
  assign T9347 = T9352 ? T9350 : T9348;
  assign T9348 = T9349 ? counts_553 : counts_552;
  assign T9349 = T8251[1'h0:1'h0];
  assign T9350 = T9351 ? counts_555 : counts_554;
  assign T9351 = T8251[1'h0:1'h0];
  assign T9352 = T8251[1'h1:1'h1];
  assign T9353 = T9358 ? T9356 : T9354;
  assign T9354 = T9355 ? counts_557 : counts_556;
  assign T9355 = T8251[1'h0:1'h0];
  assign T9356 = T9357 ? counts_559 : counts_558;
  assign T9357 = T8251[1'h0:1'h0];
  assign T9358 = T8251[1'h1:1'h1];
  assign T9359 = T8251[2'h2:2'h2];
  assign T9360 = T8251[2'h3:2'h3];
  assign T9361 = T9390 ? T9376 : T9362;
  assign T9362 = T9375 ? T9369 : T9363;
  assign T9363 = T9368 ? T9366 : T9364;
  assign T9364 = T9365 ? counts_561 : counts_560;
  assign T9365 = T8251[1'h0:1'h0];
  assign T9366 = T9367 ? counts_563 : counts_562;
  assign T9367 = T8251[1'h0:1'h0];
  assign T9368 = T8251[1'h1:1'h1];
  assign T9369 = T9374 ? T9372 : T9370;
  assign T9370 = T9371 ? counts_565 : counts_564;
  assign T9371 = T8251[1'h0:1'h0];
  assign T9372 = T9373 ? counts_567 : counts_566;
  assign T9373 = T8251[1'h0:1'h0];
  assign T9374 = T8251[1'h1:1'h1];
  assign T9375 = T8251[2'h2:2'h2];
  assign T9376 = T9389 ? T9383 : T9377;
  assign T9377 = T9382 ? T9380 : T9378;
  assign T9378 = T9379 ? counts_569 : counts_568;
  assign T9379 = T8251[1'h0:1'h0];
  assign T9380 = T9381 ? counts_571 : counts_570;
  assign T9381 = T8251[1'h0:1'h0];
  assign T9382 = T8251[1'h1:1'h1];
  assign T9383 = T9388 ? T9386 : T9384;
  assign T9384 = T9385 ? counts_573 : counts_572;
  assign T9385 = T8251[1'h0:1'h0];
  assign T9386 = T9387 ? counts_575 : counts_574;
  assign T9387 = T8251[1'h0:1'h0];
  assign T9388 = T8251[1'h1:1'h1];
  assign T9389 = T8251[2'h2:2'h2];
  assign T9390 = T8251[2'h3:2'h3];
  assign T9391 = T8251[3'h4:3'h4];
  assign T9392 = T8251[3'h5:3'h5];
  assign T9393 = T9518 ? T9456 : T9394;
  assign T9394 = T9455 ? T9425 : T9395;
  assign T9395 = T9424 ? T9410 : T9396;
  assign T9396 = T9409 ? T9403 : T9397;
  assign T9397 = T9402 ? T9400 : T9398;
  assign T9398 = T9399 ? counts_577 : counts_576;
  assign T9399 = T8251[1'h0:1'h0];
  assign T9400 = T9401 ? counts_579 : counts_578;
  assign T9401 = T8251[1'h0:1'h0];
  assign T9402 = T8251[1'h1:1'h1];
  assign T9403 = T9408 ? T9406 : T9404;
  assign T9404 = T9405 ? counts_581 : counts_580;
  assign T9405 = T8251[1'h0:1'h0];
  assign T9406 = T9407 ? counts_583 : counts_582;
  assign T9407 = T8251[1'h0:1'h0];
  assign T9408 = T8251[1'h1:1'h1];
  assign T9409 = T8251[2'h2:2'h2];
  assign T9410 = T9423 ? T9417 : T9411;
  assign T9411 = T9416 ? T9414 : T9412;
  assign T9412 = T9413 ? counts_585 : counts_584;
  assign T9413 = T8251[1'h0:1'h0];
  assign T9414 = T9415 ? counts_587 : counts_586;
  assign T9415 = T8251[1'h0:1'h0];
  assign T9416 = T8251[1'h1:1'h1];
  assign T9417 = T9422 ? T9420 : T9418;
  assign T9418 = T9419 ? counts_589 : counts_588;
  assign T9419 = T8251[1'h0:1'h0];
  assign T9420 = T9421 ? counts_591 : counts_590;
  assign T9421 = T8251[1'h0:1'h0];
  assign T9422 = T8251[1'h1:1'h1];
  assign T9423 = T8251[2'h2:2'h2];
  assign T9424 = T8251[2'h3:2'h3];
  assign T9425 = T9454 ? T9440 : T9426;
  assign T9426 = T9439 ? T9433 : T9427;
  assign T9427 = T9432 ? T9430 : T9428;
  assign T9428 = T9429 ? counts_593 : counts_592;
  assign T9429 = T8251[1'h0:1'h0];
  assign T9430 = T9431 ? counts_595 : counts_594;
  assign T9431 = T8251[1'h0:1'h0];
  assign T9432 = T8251[1'h1:1'h1];
  assign T9433 = T9438 ? T9436 : T9434;
  assign T9434 = T9435 ? counts_597 : counts_596;
  assign T9435 = T8251[1'h0:1'h0];
  assign T9436 = T9437 ? counts_599 : counts_598;
  assign T9437 = T8251[1'h0:1'h0];
  assign T9438 = T8251[1'h1:1'h1];
  assign T9439 = T8251[2'h2:2'h2];
  assign T9440 = T9453 ? T9447 : T9441;
  assign T9441 = T9446 ? T9444 : T9442;
  assign T9442 = T9443 ? counts_601 : counts_600;
  assign T9443 = T8251[1'h0:1'h0];
  assign T9444 = T9445 ? counts_603 : counts_602;
  assign T9445 = T8251[1'h0:1'h0];
  assign T9446 = T8251[1'h1:1'h1];
  assign T9447 = T9452 ? T9450 : T9448;
  assign T9448 = T9449 ? counts_605 : counts_604;
  assign T9449 = T8251[1'h0:1'h0];
  assign T9450 = T9451 ? counts_607 : counts_606;
  assign T9451 = T8251[1'h0:1'h0];
  assign T9452 = T8251[1'h1:1'h1];
  assign T9453 = T8251[2'h2:2'h2];
  assign T9454 = T8251[2'h3:2'h3];
  assign T9455 = T8251[3'h4:3'h4];
  assign T9456 = T9517 ? T9487 : T9457;
  assign T9457 = T9486 ? T9472 : T9458;
  assign T9458 = T9471 ? T9465 : T9459;
  assign T9459 = T9464 ? T9462 : T9460;
  assign T9460 = T9461 ? counts_609 : counts_608;
  assign T9461 = T8251[1'h0:1'h0];
  assign T9462 = T9463 ? counts_611 : counts_610;
  assign T9463 = T8251[1'h0:1'h0];
  assign T9464 = T8251[1'h1:1'h1];
  assign T9465 = T9470 ? T9468 : T9466;
  assign T9466 = T9467 ? counts_613 : counts_612;
  assign T9467 = T8251[1'h0:1'h0];
  assign T9468 = T9469 ? counts_615 : counts_614;
  assign T9469 = T8251[1'h0:1'h0];
  assign T9470 = T8251[1'h1:1'h1];
  assign T9471 = T8251[2'h2:2'h2];
  assign T9472 = T9485 ? T9479 : T9473;
  assign T9473 = T9478 ? T9476 : T9474;
  assign T9474 = T9475 ? counts_617 : counts_616;
  assign T9475 = T8251[1'h0:1'h0];
  assign T9476 = T9477 ? counts_619 : counts_618;
  assign T9477 = T8251[1'h0:1'h0];
  assign T9478 = T8251[1'h1:1'h1];
  assign T9479 = T9484 ? T9482 : T9480;
  assign T9480 = T9481 ? counts_621 : counts_620;
  assign T9481 = T8251[1'h0:1'h0];
  assign T9482 = T9483 ? counts_623 : counts_622;
  assign T9483 = T8251[1'h0:1'h0];
  assign T9484 = T8251[1'h1:1'h1];
  assign T9485 = T8251[2'h2:2'h2];
  assign T9486 = T8251[2'h3:2'h3];
  assign T9487 = T9516 ? T9502 : T9488;
  assign T9488 = T9501 ? T9495 : T9489;
  assign T9489 = T9494 ? T9492 : T9490;
  assign T9490 = T9491 ? counts_625 : counts_624;
  assign T9491 = T8251[1'h0:1'h0];
  assign T9492 = T9493 ? counts_627 : counts_626;
  assign T9493 = T8251[1'h0:1'h0];
  assign T9494 = T8251[1'h1:1'h1];
  assign T9495 = T9500 ? T9498 : T9496;
  assign T9496 = T9497 ? counts_629 : counts_628;
  assign T9497 = T8251[1'h0:1'h0];
  assign T9498 = T9499 ? counts_631 : counts_630;
  assign T9499 = T8251[1'h0:1'h0];
  assign T9500 = T8251[1'h1:1'h1];
  assign T9501 = T8251[2'h2:2'h2];
  assign T9502 = T9515 ? T9509 : T9503;
  assign T9503 = T9508 ? T9506 : T9504;
  assign T9504 = T9505 ? counts_633 : counts_632;
  assign T9505 = T8251[1'h0:1'h0];
  assign T9506 = T9507 ? counts_635 : counts_634;
  assign T9507 = T8251[1'h0:1'h0];
  assign T9508 = T8251[1'h1:1'h1];
  assign T9509 = T9514 ? T9512 : T9510;
  assign T9510 = T9511 ? counts_637 : counts_636;
  assign T9511 = T8251[1'h0:1'h0];
  assign T9512 = T9513 ? counts_639 : counts_638;
  assign T9513 = T8251[1'h0:1'h0];
  assign T9514 = T8251[1'h1:1'h1];
  assign T9515 = T8251[2'h2:2'h2];
  assign T9516 = T8251[2'h3:2'h3];
  assign T9517 = T8251[3'h4:3'h4];
  assign T9518 = T8251[3'h5:3'h5];
  assign T9519 = T8251[3'h6:3'h6];
  assign T9520 = T9773 ? T9647 : T9521;
  assign T9521 = T9646 ? T9584 : T9522;
  assign T9522 = T9583 ? T9553 : T9523;
  assign T9523 = T9552 ? T9538 : T9524;
  assign T9524 = T9537 ? T9531 : T9525;
  assign T9525 = T9530 ? T9528 : T9526;
  assign T9526 = T9527 ? counts_641 : counts_640;
  assign T9527 = T8251[1'h0:1'h0];
  assign T9528 = T9529 ? counts_643 : counts_642;
  assign T9529 = T8251[1'h0:1'h0];
  assign T9530 = T8251[1'h1:1'h1];
  assign T9531 = T9536 ? T9534 : T9532;
  assign T9532 = T9533 ? counts_645 : counts_644;
  assign T9533 = T8251[1'h0:1'h0];
  assign T9534 = T9535 ? counts_647 : counts_646;
  assign T9535 = T8251[1'h0:1'h0];
  assign T9536 = T8251[1'h1:1'h1];
  assign T9537 = T8251[2'h2:2'h2];
  assign T9538 = T9551 ? T9545 : T9539;
  assign T9539 = T9544 ? T9542 : T9540;
  assign T9540 = T9541 ? counts_649 : counts_648;
  assign T9541 = T8251[1'h0:1'h0];
  assign T9542 = T9543 ? counts_651 : counts_650;
  assign T9543 = T8251[1'h0:1'h0];
  assign T9544 = T8251[1'h1:1'h1];
  assign T9545 = T9550 ? T9548 : T9546;
  assign T9546 = T9547 ? counts_653 : counts_652;
  assign T9547 = T8251[1'h0:1'h0];
  assign T9548 = T9549 ? counts_655 : counts_654;
  assign T9549 = T8251[1'h0:1'h0];
  assign T9550 = T8251[1'h1:1'h1];
  assign T9551 = T8251[2'h2:2'h2];
  assign T9552 = T8251[2'h3:2'h3];
  assign T9553 = T9582 ? T9568 : T9554;
  assign T9554 = T9567 ? T9561 : T9555;
  assign T9555 = T9560 ? T9558 : T9556;
  assign T9556 = T9557 ? counts_657 : counts_656;
  assign T9557 = T8251[1'h0:1'h0];
  assign T9558 = T9559 ? counts_659 : counts_658;
  assign T9559 = T8251[1'h0:1'h0];
  assign T9560 = T8251[1'h1:1'h1];
  assign T9561 = T9566 ? T9564 : T9562;
  assign T9562 = T9563 ? counts_661 : counts_660;
  assign T9563 = T8251[1'h0:1'h0];
  assign T9564 = T9565 ? counts_663 : counts_662;
  assign T9565 = T8251[1'h0:1'h0];
  assign T9566 = T8251[1'h1:1'h1];
  assign T9567 = T8251[2'h2:2'h2];
  assign T9568 = T9581 ? T9575 : T9569;
  assign T9569 = T9574 ? T9572 : T9570;
  assign T9570 = T9571 ? counts_665 : counts_664;
  assign T9571 = T8251[1'h0:1'h0];
  assign T9572 = T9573 ? counts_667 : counts_666;
  assign T9573 = T8251[1'h0:1'h0];
  assign T9574 = T8251[1'h1:1'h1];
  assign T9575 = T9580 ? T9578 : T9576;
  assign T9576 = T9577 ? counts_669 : counts_668;
  assign T9577 = T8251[1'h0:1'h0];
  assign T9578 = T9579 ? counts_671 : counts_670;
  assign T9579 = T8251[1'h0:1'h0];
  assign T9580 = T8251[1'h1:1'h1];
  assign T9581 = T8251[2'h2:2'h2];
  assign T9582 = T8251[2'h3:2'h3];
  assign T9583 = T8251[3'h4:3'h4];
  assign T9584 = T9645 ? T9615 : T9585;
  assign T9585 = T9614 ? T9600 : T9586;
  assign T9586 = T9599 ? T9593 : T9587;
  assign T9587 = T9592 ? T9590 : T9588;
  assign T9588 = T9589 ? counts_673 : counts_672;
  assign T9589 = T8251[1'h0:1'h0];
  assign T9590 = T9591 ? counts_675 : counts_674;
  assign T9591 = T8251[1'h0:1'h0];
  assign T9592 = T8251[1'h1:1'h1];
  assign T9593 = T9598 ? T9596 : T9594;
  assign T9594 = T9595 ? counts_677 : counts_676;
  assign T9595 = T8251[1'h0:1'h0];
  assign T9596 = T9597 ? counts_679 : counts_678;
  assign T9597 = T8251[1'h0:1'h0];
  assign T9598 = T8251[1'h1:1'h1];
  assign T9599 = T8251[2'h2:2'h2];
  assign T9600 = T9613 ? T9607 : T9601;
  assign T9601 = T9606 ? T9604 : T9602;
  assign T9602 = T9603 ? counts_681 : counts_680;
  assign T9603 = T8251[1'h0:1'h0];
  assign T9604 = T9605 ? counts_683 : counts_682;
  assign T9605 = T8251[1'h0:1'h0];
  assign T9606 = T8251[1'h1:1'h1];
  assign T9607 = T9612 ? T9610 : T9608;
  assign T9608 = T9609 ? counts_685 : counts_684;
  assign T9609 = T8251[1'h0:1'h0];
  assign T9610 = T9611 ? counts_687 : counts_686;
  assign T9611 = T8251[1'h0:1'h0];
  assign T9612 = T8251[1'h1:1'h1];
  assign T9613 = T8251[2'h2:2'h2];
  assign T9614 = T8251[2'h3:2'h3];
  assign T9615 = T9644 ? T9630 : T9616;
  assign T9616 = T9629 ? T9623 : T9617;
  assign T9617 = T9622 ? T9620 : T9618;
  assign T9618 = T9619 ? counts_689 : counts_688;
  assign T9619 = T8251[1'h0:1'h0];
  assign T9620 = T9621 ? counts_691 : counts_690;
  assign T9621 = T8251[1'h0:1'h0];
  assign T9622 = T8251[1'h1:1'h1];
  assign T9623 = T9628 ? T9626 : T9624;
  assign T9624 = T9625 ? counts_693 : counts_692;
  assign T9625 = T8251[1'h0:1'h0];
  assign T9626 = T9627 ? counts_695 : counts_694;
  assign T9627 = T8251[1'h0:1'h0];
  assign T9628 = T8251[1'h1:1'h1];
  assign T9629 = T8251[2'h2:2'h2];
  assign T9630 = T9643 ? T9637 : T9631;
  assign T9631 = T9636 ? T9634 : T9632;
  assign T9632 = T9633 ? counts_697 : counts_696;
  assign T9633 = T8251[1'h0:1'h0];
  assign T9634 = T9635 ? counts_699 : counts_698;
  assign T9635 = T8251[1'h0:1'h0];
  assign T9636 = T8251[1'h1:1'h1];
  assign T9637 = T9642 ? T9640 : T9638;
  assign T9638 = T9639 ? counts_701 : counts_700;
  assign T9639 = T8251[1'h0:1'h0];
  assign T9640 = T9641 ? counts_703 : counts_702;
  assign T9641 = T8251[1'h0:1'h0];
  assign T9642 = T8251[1'h1:1'h1];
  assign T9643 = T8251[2'h2:2'h2];
  assign T9644 = T8251[2'h3:2'h3];
  assign T9645 = T8251[3'h4:3'h4];
  assign T9646 = T8251[3'h5:3'h5];
  assign T9647 = T9772 ? T9710 : T9648;
  assign T9648 = T9709 ? T9679 : T9649;
  assign T9649 = T9678 ? T9664 : T9650;
  assign T9650 = T9663 ? T9657 : T9651;
  assign T9651 = T9656 ? T9654 : T9652;
  assign T9652 = T9653 ? counts_705 : counts_704;
  assign T9653 = T8251[1'h0:1'h0];
  assign T9654 = T9655 ? counts_707 : counts_706;
  assign T9655 = T8251[1'h0:1'h0];
  assign T9656 = T8251[1'h1:1'h1];
  assign T9657 = T9662 ? T9660 : T9658;
  assign T9658 = T9659 ? counts_709 : counts_708;
  assign T9659 = T8251[1'h0:1'h0];
  assign T9660 = T9661 ? counts_711 : counts_710;
  assign T9661 = T8251[1'h0:1'h0];
  assign T9662 = T8251[1'h1:1'h1];
  assign T9663 = T8251[2'h2:2'h2];
  assign T9664 = T9677 ? T9671 : T9665;
  assign T9665 = T9670 ? T9668 : T9666;
  assign T9666 = T9667 ? counts_713 : counts_712;
  assign T9667 = T8251[1'h0:1'h0];
  assign T9668 = T9669 ? counts_715 : counts_714;
  assign T9669 = T8251[1'h0:1'h0];
  assign T9670 = T8251[1'h1:1'h1];
  assign T9671 = T9676 ? T9674 : T9672;
  assign T9672 = T9673 ? counts_717 : counts_716;
  assign T9673 = T8251[1'h0:1'h0];
  assign T9674 = T9675 ? counts_719 : counts_718;
  assign T9675 = T8251[1'h0:1'h0];
  assign T9676 = T8251[1'h1:1'h1];
  assign T9677 = T8251[2'h2:2'h2];
  assign T9678 = T8251[2'h3:2'h3];
  assign T9679 = T9708 ? T9694 : T9680;
  assign T9680 = T9693 ? T9687 : T9681;
  assign T9681 = T9686 ? T9684 : T9682;
  assign T9682 = T9683 ? counts_721 : counts_720;
  assign T9683 = T8251[1'h0:1'h0];
  assign T9684 = T9685 ? counts_723 : counts_722;
  assign T9685 = T8251[1'h0:1'h0];
  assign T9686 = T8251[1'h1:1'h1];
  assign T9687 = T9692 ? T9690 : T9688;
  assign T9688 = T9689 ? counts_725 : counts_724;
  assign T9689 = T8251[1'h0:1'h0];
  assign T9690 = T9691 ? counts_727 : counts_726;
  assign T9691 = T8251[1'h0:1'h0];
  assign T9692 = T8251[1'h1:1'h1];
  assign T9693 = T8251[2'h2:2'h2];
  assign T9694 = T9707 ? T9701 : T9695;
  assign T9695 = T9700 ? T9698 : T9696;
  assign T9696 = T9697 ? counts_729 : counts_728;
  assign T9697 = T8251[1'h0:1'h0];
  assign T9698 = T9699 ? counts_731 : counts_730;
  assign T9699 = T8251[1'h0:1'h0];
  assign T9700 = T8251[1'h1:1'h1];
  assign T9701 = T9706 ? T9704 : T9702;
  assign T9702 = T9703 ? counts_733 : counts_732;
  assign T9703 = T8251[1'h0:1'h0];
  assign T9704 = T9705 ? counts_735 : counts_734;
  assign T9705 = T8251[1'h0:1'h0];
  assign T9706 = T8251[1'h1:1'h1];
  assign T9707 = T8251[2'h2:2'h2];
  assign T9708 = T8251[2'h3:2'h3];
  assign T9709 = T8251[3'h4:3'h4];
  assign T9710 = T9771 ? T9741 : T9711;
  assign T9711 = T9740 ? T9726 : T9712;
  assign T9712 = T9725 ? T9719 : T9713;
  assign T9713 = T9718 ? T9716 : T9714;
  assign T9714 = T9715 ? counts_737 : counts_736;
  assign T9715 = T8251[1'h0:1'h0];
  assign T9716 = T9717 ? counts_739 : counts_738;
  assign T9717 = T8251[1'h0:1'h0];
  assign T9718 = T8251[1'h1:1'h1];
  assign T9719 = T9724 ? T9722 : T9720;
  assign T9720 = T9721 ? counts_741 : counts_740;
  assign T9721 = T8251[1'h0:1'h0];
  assign T9722 = T9723 ? counts_743 : counts_742;
  assign T9723 = T8251[1'h0:1'h0];
  assign T9724 = T8251[1'h1:1'h1];
  assign T9725 = T8251[2'h2:2'h2];
  assign T9726 = T9739 ? T9733 : T9727;
  assign T9727 = T9732 ? T9730 : T9728;
  assign T9728 = T9729 ? counts_745 : counts_744;
  assign T9729 = T8251[1'h0:1'h0];
  assign T9730 = T9731 ? counts_747 : counts_746;
  assign T9731 = T8251[1'h0:1'h0];
  assign T9732 = T8251[1'h1:1'h1];
  assign T9733 = T9738 ? T9736 : T9734;
  assign T9734 = T9735 ? counts_749 : counts_748;
  assign T9735 = T8251[1'h0:1'h0];
  assign T9736 = T9737 ? counts_751 : counts_750;
  assign T9737 = T8251[1'h0:1'h0];
  assign T9738 = T8251[1'h1:1'h1];
  assign T9739 = T8251[2'h2:2'h2];
  assign T9740 = T8251[2'h3:2'h3];
  assign T9741 = T9770 ? T9756 : T9742;
  assign T9742 = T9755 ? T9749 : T9743;
  assign T9743 = T9748 ? T9746 : T9744;
  assign T9744 = T9745 ? counts_753 : counts_752;
  assign T9745 = T8251[1'h0:1'h0];
  assign T9746 = T9747 ? counts_755 : counts_754;
  assign T9747 = T8251[1'h0:1'h0];
  assign T9748 = T8251[1'h1:1'h1];
  assign T9749 = T9754 ? T9752 : T9750;
  assign T9750 = T9751 ? counts_757 : counts_756;
  assign T9751 = T8251[1'h0:1'h0];
  assign T9752 = T9753 ? counts_759 : counts_758;
  assign T9753 = T8251[1'h0:1'h0];
  assign T9754 = T8251[1'h1:1'h1];
  assign T9755 = T8251[2'h2:2'h2];
  assign T9756 = T9769 ? T9763 : T9757;
  assign T9757 = T9762 ? T9760 : T9758;
  assign T9758 = T9759 ? counts_761 : counts_760;
  assign T9759 = T8251[1'h0:1'h0];
  assign T9760 = T9761 ? counts_763 : counts_762;
  assign T9761 = T8251[1'h0:1'h0];
  assign T9762 = T8251[1'h1:1'h1];
  assign T9763 = T9768 ? T9766 : T9764;
  assign T9764 = T9765 ? counts_765 : counts_764;
  assign T9765 = T8251[1'h0:1'h0];
  assign T9766 = T9767 ? counts_767 : counts_766;
  assign T9767 = T8251[1'h0:1'h0];
  assign T9768 = T8251[1'h1:1'h1];
  assign T9769 = T8251[2'h2:2'h2];
  assign T9770 = T8251[2'h3:2'h3];
  assign T9771 = T8251[3'h4:3'h4];
  assign T9772 = T8251[3'h5:3'h5];
  assign T9773 = T8251[3'h6:3'h6];
  assign T9774 = T8251[3'h7:3'h7];
  assign T9775 = T10284 ? T10030 : T9776;
  assign T9776 = T10029 ? T9903 : T9777;
  assign T9777 = T9902 ? T9840 : T9778;
  assign T9778 = T9839 ? T9809 : T9779;
  assign T9779 = T9808 ? T9794 : T9780;
  assign T9780 = T9793 ? T9787 : T9781;
  assign T9781 = T9786 ? T9784 : T9782;
  assign T9782 = T9783 ? counts_769 : counts_768;
  assign T9783 = T8251[1'h0:1'h0];
  assign T9784 = T9785 ? counts_771 : counts_770;
  assign T9785 = T8251[1'h0:1'h0];
  assign T9786 = T8251[1'h1:1'h1];
  assign T9787 = T9792 ? T9790 : T9788;
  assign T9788 = T9789 ? counts_773 : counts_772;
  assign T9789 = T8251[1'h0:1'h0];
  assign T9790 = T9791 ? counts_775 : counts_774;
  assign T9791 = T8251[1'h0:1'h0];
  assign T9792 = T8251[1'h1:1'h1];
  assign T9793 = T8251[2'h2:2'h2];
  assign T9794 = T9807 ? T9801 : T9795;
  assign T9795 = T9800 ? T9798 : T9796;
  assign T9796 = T9797 ? counts_777 : counts_776;
  assign T9797 = T8251[1'h0:1'h0];
  assign T9798 = T9799 ? counts_779 : counts_778;
  assign T9799 = T8251[1'h0:1'h0];
  assign T9800 = T8251[1'h1:1'h1];
  assign T9801 = T9806 ? T9804 : T9802;
  assign T9802 = T9803 ? counts_781 : counts_780;
  assign T9803 = T8251[1'h0:1'h0];
  assign T9804 = T9805 ? counts_783 : counts_782;
  assign T9805 = T8251[1'h0:1'h0];
  assign T9806 = T8251[1'h1:1'h1];
  assign T9807 = T8251[2'h2:2'h2];
  assign T9808 = T8251[2'h3:2'h3];
  assign T9809 = T9838 ? T9824 : T9810;
  assign T9810 = T9823 ? T9817 : T9811;
  assign T9811 = T9816 ? T9814 : T9812;
  assign T9812 = T9813 ? counts_785 : counts_784;
  assign T9813 = T8251[1'h0:1'h0];
  assign T9814 = T9815 ? counts_787 : counts_786;
  assign T9815 = T8251[1'h0:1'h0];
  assign T9816 = T8251[1'h1:1'h1];
  assign T9817 = T9822 ? T9820 : T9818;
  assign T9818 = T9819 ? counts_789 : counts_788;
  assign T9819 = T8251[1'h0:1'h0];
  assign T9820 = T9821 ? counts_791 : counts_790;
  assign T9821 = T8251[1'h0:1'h0];
  assign T9822 = T8251[1'h1:1'h1];
  assign T9823 = T8251[2'h2:2'h2];
  assign T9824 = T9837 ? T9831 : T9825;
  assign T9825 = T9830 ? T9828 : T9826;
  assign T9826 = T9827 ? counts_793 : counts_792;
  assign T9827 = T8251[1'h0:1'h0];
  assign T9828 = T9829 ? counts_795 : counts_794;
  assign T9829 = T8251[1'h0:1'h0];
  assign T9830 = T8251[1'h1:1'h1];
  assign T9831 = T9836 ? T9834 : T9832;
  assign T9832 = T9833 ? counts_797 : counts_796;
  assign T9833 = T8251[1'h0:1'h0];
  assign T9834 = T9835 ? counts_799 : counts_798;
  assign T9835 = T8251[1'h0:1'h0];
  assign T9836 = T8251[1'h1:1'h1];
  assign T9837 = T8251[2'h2:2'h2];
  assign T9838 = T8251[2'h3:2'h3];
  assign T9839 = T8251[3'h4:3'h4];
  assign T9840 = T9901 ? T9871 : T9841;
  assign T9841 = T9870 ? T9856 : T9842;
  assign T9842 = T9855 ? T9849 : T9843;
  assign T9843 = T9848 ? T9846 : T9844;
  assign T9844 = T9845 ? counts_801 : counts_800;
  assign T9845 = T8251[1'h0:1'h0];
  assign T9846 = T9847 ? counts_803 : counts_802;
  assign T9847 = T8251[1'h0:1'h0];
  assign T9848 = T8251[1'h1:1'h1];
  assign T9849 = T9854 ? T9852 : T9850;
  assign T9850 = T9851 ? counts_805 : counts_804;
  assign T9851 = T8251[1'h0:1'h0];
  assign T9852 = T9853 ? counts_807 : counts_806;
  assign T9853 = T8251[1'h0:1'h0];
  assign T9854 = T8251[1'h1:1'h1];
  assign T9855 = T8251[2'h2:2'h2];
  assign T9856 = T9869 ? T9863 : T9857;
  assign T9857 = T9862 ? T9860 : T9858;
  assign T9858 = T9859 ? counts_809 : counts_808;
  assign T9859 = T8251[1'h0:1'h0];
  assign T9860 = T9861 ? counts_811 : counts_810;
  assign T9861 = T8251[1'h0:1'h0];
  assign T9862 = T8251[1'h1:1'h1];
  assign T9863 = T9868 ? T9866 : T9864;
  assign T9864 = T9865 ? counts_813 : counts_812;
  assign T9865 = T8251[1'h0:1'h0];
  assign T9866 = T9867 ? counts_815 : counts_814;
  assign T9867 = T8251[1'h0:1'h0];
  assign T9868 = T8251[1'h1:1'h1];
  assign T9869 = T8251[2'h2:2'h2];
  assign T9870 = T8251[2'h3:2'h3];
  assign T9871 = T9900 ? T9886 : T9872;
  assign T9872 = T9885 ? T9879 : T9873;
  assign T9873 = T9878 ? T9876 : T9874;
  assign T9874 = T9875 ? counts_817 : counts_816;
  assign T9875 = T8251[1'h0:1'h0];
  assign T9876 = T9877 ? counts_819 : counts_818;
  assign T9877 = T8251[1'h0:1'h0];
  assign T9878 = T8251[1'h1:1'h1];
  assign T9879 = T9884 ? T9882 : T9880;
  assign T9880 = T9881 ? counts_821 : counts_820;
  assign T9881 = T8251[1'h0:1'h0];
  assign T9882 = T9883 ? counts_823 : counts_822;
  assign T9883 = T8251[1'h0:1'h0];
  assign T9884 = T8251[1'h1:1'h1];
  assign T9885 = T8251[2'h2:2'h2];
  assign T9886 = T9899 ? T9893 : T9887;
  assign T9887 = T9892 ? T9890 : T9888;
  assign T9888 = T9889 ? counts_825 : counts_824;
  assign T9889 = T8251[1'h0:1'h0];
  assign T9890 = T9891 ? counts_827 : counts_826;
  assign T9891 = T8251[1'h0:1'h0];
  assign T9892 = T8251[1'h1:1'h1];
  assign T9893 = T9898 ? T9896 : T9894;
  assign T9894 = T9895 ? counts_829 : counts_828;
  assign T9895 = T8251[1'h0:1'h0];
  assign T9896 = T9897 ? counts_831 : counts_830;
  assign T9897 = T8251[1'h0:1'h0];
  assign T9898 = T8251[1'h1:1'h1];
  assign T9899 = T8251[2'h2:2'h2];
  assign T9900 = T8251[2'h3:2'h3];
  assign T9901 = T8251[3'h4:3'h4];
  assign T9902 = T8251[3'h5:3'h5];
  assign T9903 = T10028 ? T9966 : T9904;
  assign T9904 = T9965 ? T9935 : T9905;
  assign T9905 = T9934 ? T9920 : T9906;
  assign T9906 = T9919 ? T9913 : T9907;
  assign T9907 = T9912 ? T9910 : T9908;
  assign T9908 = T9909 ? counts_833 : counts_832;
  assign T9909 = T8251[1'h0:1'h0];
  assign T9910 = T9911 ? counts_835 : counts_834;
  assign T9911 = T8251[1'h0:1'h0];
  assign T9912 = T8251[1'h1:1'h1];
  assign T9913 = T9918 ? T9916 : T9914;
  assign T9914 = T9915 ? counts_837 : counts_836;
  assign T9915 = T8251[1'h0:1'h0];
  assign T9916 = T9917 ? counts_839 : counts_838;
  assign T9917 = T8251[1'h0:1'h0];
  assign T9918 = T8251[1'h1:1'h1];
  assign T9919 = T8251[2'h2:2'h2];
  assign T9920 = T9933 ? T9927 : T9921;
  assign T9921 = T9926 ? T9924 : T9922;
  assign T9922 = T9923 ? counts_841 : counts_840;
  assign T9923 = T8251[1'h0:1'h0];
  assign T9924 = T9925 ? counts_843 : counts_842;
  assign T9925 = T8251[1'h0:1'h0];
  assign T9926 = T8251[1'h1:1'h1];
  assign T9927 = T9932 ? T9930 : T9928;
  assign T9928 = T9929 ? counts_845 : counts_844;
  assign T9929 = T8251[1'h0:1'h0];
  assign T9930 = T9931 ? counts_847 : counts_846;
  assign T9931 = T8251[1'h0:1'h0];
  assign T9932 = T8251[1'h1:1'h1];
  assign T9933 = T8251[2'h2:2'h2];
  assign T9934 = T8251[2'h3:2'h3];
  assign T9935 = T9964 ? T9950 : T9936;
  assign T9936 = T9949 ? T9943 : T9937;
  assign T9937 = T9942 ? T9940 : T9938;
  assign T9938 = T9939 ? counts_849 : counts_848;
  assign T9939 = T8251[1'h0:1'h0];
  assign T9940 = T9941 ? counts_851 : counts_850;
  assign T9941 = T8251[1'h0:1'h0];
  assign T9942 = T8251[1'h1:1'h1];
  assign T9943 = T9948 ? T9946 : T9944;
  assign T9944 = T9945 ? counts_853 : counts_852;
  assign T9945 = T8251[1'h0:1'h0];
  assign T9946 = T9947 ? counts_855 : counts_854;
  assign T9947 = T8251[1'h0:1'h0];
  assign T9948 = T8251[1'h1:1'h1];
  assign T9949 = T8251[2'h2:2'h2];
  assign T9950 = T9963 ? T9957 : T9951;
  assign T9951 = T9956 ? T9954 : T9952;
  assign T9952 = T9953 ? counts_857 : counts_856;
  assign T9953 = T8251[1'h0:1'h0];
  assign T9954 = T9955 ? counts_859 : counts_858;
  assign T9955 = T8251[1'h0:1'h0];
  assign T9956 = T8251[1'h1:1'h1];
  assign T9957 = T9962 ? T9960 : T9958;
  assign T9958 = T9959 ? counts_861 : counts_860;
  assign T9959 = T8251[1'h0:1'h0];
  assign T9960 = T9961 ? counts_863 : counts_862;
  assign T9961 = T8251[1'h0:1'h0];
  assign T9962 = T8251[1'h1:1'h1];
  assign T9963 = T8251[2'h2:2'h2];
  assign T9964 = T8251[2'h3:2'h3];
  assign T9965 = T8251[3'h4:3'h4];
  assign T9966 = T10027 ? T9997 : T9967;
  assign T9967 = T9996 ? T9982 : T9968;
  assign T9968 = T9981 ? T9975 : T9969;
  assign T9969 = T9974 ? T9972 : T9970;
  assign T9970 = T9971 ? counts_865 : counts_864;
  assign T9971 = T8251[1'h0:1'h0];
  assign T9972 = T9973 ? counts_867 : counts_866;
  assign T9973 = T8251[1'h0:1'h0];
  assign T9974 = T8251[1'h1:1'h1];
  assign T9975 = T9980 ? T9978 : T9976;
  assign T9976 = T9977 ? counts_869 : counts_868;
  assign T9977 = T8251[1'h0:1'h0];
  assign T9978 = T9979 ? counts_871 : counts_870;
  assign T9979 = T8251[1'h0:1'h0];
  assign T9980 = T8251[1'h1:1'h1];
  assign T9981 = T8251[2'h2:2'h2];
  assign T9982 = T9995 ? T9989 : T9983;
  assign T9983 = T9988 ? T9986 : T9984;
  assign T9984 = T9985 ? counts_873 : counts_872;
  assign T9985 = T8251[1'h0:1'h0];
  assign T9986 = T9987 ? counts_875 : counts_874;
  assign T9987 = T8251[1'h0:1'h0];
  assign T9988 = T8251[1'h1:1'h1];
  assign T9989 = T9994 ? T9992 : T9990;
  assign T9990 = T9991 ? counts_877 : counts_876;
  assign T9991 = T8251[1'h0:1'h0];
  assign T9992 = T9993 ? counts_879 : counts_878;
  assign T9993 = T8251[1'h0:1'h0];
  assign T9994 = T8251[1'h1:1'h1];
  assign T9995 = T8251[2'h2:2'h2];
  assign T9996 = T8251[2'h3:2'h3];
  assign T9997 = T10026 ? T10012 : T9998;
  assign T9998 = T10011 ? T10005 : T9999;
  assign T9999 = T10004 ? T10002 : T10000;
  assign T10000 = T10001 ? counts_881 : counts_880;
  assign T10001 = T8251[1'h0:1'h0];
  assign T10002 = T10003 ? counts_883 : counts_882;
  assign T10003 = T8251[1'h0:1'h0];
  assign T10004 = T8251[1'h1:1'h1];
  assign T10005 = T10010 ? T10008 : T10006;
  assign T10006 = T10007 ? counts_885 : counts_884;
  assign T10007 = T8251[1'h0:1'h0];
  assign T10008 = T10009 ? counts_887 : counts_886;
  assign T10009 = T8251[1'h0:1'h0];
  assign T10010 = T8251[1'h1:1'h1];
  assign T10011 = T8251[2'h2:2'h2];
  assign T10012 = T10025 ? T10019 : T10013;
  assign T10013 = T10018 ? T10016 : T10014;
  assign T10014 = T10015 ? counts_889 : counts_888;
  assign T10015 = T8251[1'h0:1'h0];
  assign T10016 = T10017 ? counts_891 : counts_890;
  assign T10017 = T8251[1'h0:1'h0];
  assign T10018 = T8251[1'h1:1'h1];
  assign T10019 = T10024 ? T10022 : T10020;
  assign T10020 = T10021 ? counts_893 : counts_892;
  assign T10021 = T8251[1'h0:1'h0];
  assign T10022 = T10023 ? counts_895 : counts_894;
  assign T10023 = T8251[1'h0:1'h0];
  assign T10024 = T8251[1'h1:1'h1];
  assign T10025 = T8251[2'h2:2'h2];
  assign T10026 = T8251[2'h3:2'h3];
  assign T10027 = T8251[3'h4:3'h4];
  assign T10028 = T8251[3'h5:3'h5];
  assign T10029 = T8251[3'h6:3'h6];
  assign T10030 = T10283 ? T10157 : T10031;
  assign T10031 = T10156 ? T10094 : T10032;
  assign T10032 = T10093 ? T10063 : T10033;
  assign T10033 = T10062 ? T10048 : T10034;
  assign T10034 = T10047 ? T10041 : T10035;
  assign T10035 = T10040 ? T10038 : T10036;
  assign T10036 = T10037 ? counts_897 : counts_896;
  assign T10037 = T8251[1'h0:1'h0];
  assign T10038 = T10039 ? counts_899 : counts_898;
  assign T10039 = T8251[1'h0:1'h0];
  assign T10040 = T8251[1'h1:1'h1];
  assign T10041 = T10046 ? T10044 : T10042;
  assign T10042 = T10043 ? counts_901 : counts_900;
  assign T10043 = T8251[1'h0:1'h0];
  assign T10044 = T10045 ? counts_903 : counts_902;
  assign T10045 = T8251[1'h0:1'h0];
  assign T10046 = T8251[1'h1:1'h1];
  assign T10047 = T8251[2'h2:2'h2];
  assign T10048 = T10061 ? T10055 : T10049;
  assign T10049 = T10054 ? T10052 : T10050;
  assign T10050 = T10051 ? counts_905 : counts_904;
  assign T10051 = T8251[1'h0:1'h0];
  assign T10052 = T10053 ? counts_907 : counts_906;
  assign T10053 = T8251[1'h0:1'h0];
  assign T10054 = T8251[1'h1:1'h1];
  assign T10055 = T10060 ? T10058 : T10056;
  assign T10056 = T10057 ? counts_909 : counts_908;
  assign T10057 = T8251[1'h0:1'h0];
  assign T10058 = T10059 ? counts_911 : counts_910;
  assign T10059 = T8251[1'h0:1'h0];
  assign T10060 = T8251[1'h1:1'h1];
  assign T10061 = T8251[2'h2:2'h2];
  assign T10062 = T8251[2'h3:2'h3];
  assign T10063 = T10092 ? T10078 : T10064;
  assign T10064 = T10077 ? T10071 : T10065;
  assign T10065 = T10070 ? T10068 : T10066;
  assign T10066 = T10067 ? counts_913 : counts_912;
  assign T10067 = T8251[1'h0:1'h0];
  assign T10068 = T10069 ? counts_915 : counts_914;
  assign T10069 = T8251[1'h0:1'h0];
  assign T10070 = T8251[1'h1:1'h1];
  assign T10071 = T10076 ? T10074 : T10072;
  assign T10072 = T10073 ? counts_917 : counts_916;
  assign T10073 = T8251[1'h0:1'h0];
  assign T10074 = T10075 ? counts_919 : counts_918;
  assign T10075 = T8251[1'h0:1'h0];
  assign T10076 = T8251[1'h1:1'h1];
  assign T10077 = T8251[2'h2:2'h2];
  assign T10078 = T10091 ? T10085 : T10079;
  assign T10079 = T10084 ? T10082 : T10080;
  assign T10080 = T10081 ? counts_921 : counts_920;
  assign T10081 = T8251[1'h0:1'h0];
  assign T10082 = T10083 ? counts_923 : counts_922;
  assign T10083 = T8251[1'h0:1'h0];
  assign T10084 = T8251[1'h1:1'h1];
  assign T10085 = T10090 ? T10088 : T10086;
  assign T10086 = T10087 ? counts_925 : counts_924;
  assign T10087 = T8251[1'h0:1'h0];
  assign T10088 = T10089 ? counts_927 : counts_926;
  assign T10089 = T8251[1'h0:1'h0];
  assign T10090 = T8251[1'h1:1'h1];
  assign T10091 = T8251[2'h2:2'h2];
  assign T10092 = T8251[2'h3:2'h3];
  assign T10093 = T8251[3'h4:3'h4];
  assign T10094 = T10155 ? T10125 : T10095;
  assign T10095 = T10124 ? T10110 : T10096;
  assign T10096 = T10109 ? T10103 : T10097;
  assign T10097 = T10102 ? T10100 : T10098;
  assign T10098 = T10099 ? counts_929 : counts_928;
  assign T10099 = T8251[1'h0:1'h0];
  assign T10100 = T10101 ? counts_931 : counts_930;
  assign T10101 = T8251[1'h0:1'h0];
  assign T10102 = T8251[1'h1:1'h1];
  assign T10103 = T10108 ? T10106 : T10104;
  assign T10104 = T10105 ? counts_933 : counts_932;
  assign T10105 = T8251[1'h0:1'h0];
  assign T10106 = T10107 ? counts_935 : counts_934;
  assign T10107 = T8251[1'h0:1'h0];
  assign T10108 = T8251[1'h1:1'h1];
  assign T10109 = T8251[2'h2:2'h2];
  assign T10110 = T10123 ? T10117 : T10111;
  assign T10111 = T10116 ? T10114 : T10112;
  assign T10112 = T10113 ? counts_937 : counts_936;
  assign T10113 = T8251[1'h0:1'h0];
  assign T10114 = T10115 ? counts_939 : counts_938;
  assign T10115 = T8251[1'h0:1'h0];
  assign T10116 = T8251[1'h1:1'h1];
  assign T10117 = T10122 ? T10120 : T10118;
  assign T10118 = T10119 ? counts_941 : counts_940;
  assign T10119 = T8251[1'h0:1'h0];
  assign T10120 = T10121 ? counts_943 : counts_942;
  assign T10121 = T8251[1'h0:1'h0];
  assign T10122 = T8251[1'h1:1'h1];
  assign T10123 = T8251[2'h2:2'h2];
  assign T10124 = T8251[2'h3:2'h3];
  assign T10125 = T10154 ? T10140 : T10126;
  assign T10126 = T10139 ? T10133 : T10127;
  assign T10127 = T10132 ? T10130 : T10128;
  assign T10128 = T10129 ? counts_945 : counts_944;
  assign T10129 = T8251[1'h0:1'h0];
  assign T10130 = T10131 ? counts_947 : counts_946;
  assign T10131 = T8251[1'h0:1'h0];
  assign T10132 = T8251[1'h1:1'h1];
  assign T10133 = T10138 ? T10136 : T10134;
  assign T10134 = T10135 ? counts_949 : counts_948;
  assign T10135 = T8251[1'h0:1'h0];
  assign T10136 = T10137 ? counts_951 : counts_950;
  assign T10137 = T8251[1'h0:1'h0];
  assign T10138 = T8251[1'h1:1'h1];
  assign T10139 = T8251[2'h2:2'h2];
  assign T10140 = T10153 ? T10147 : T10141;
  assign T10141 = T10146 ? T10144 : T10142;
  assign T10142 = T10143 ? counts_953 : counts_952;
  assign T10143 = T8251[1'h0:1'h0];
  assign T10144 = T10145 ? counts_955 : counts_954;
  assign T10145 = T8251[1'h0:1'h0];
  assign T10146 = T8251[1'h1:1'h1];
  assign T10147 = T10152 ? T10150 : T10148;
  assign T10148 = T10149 ? counts_957 : counts_956;
  assign T10149 = T8251[1'h0:1'h0];
  assign T10150 = T10151 ? counts_959 : counts_958;
  assign T10151 = T8251[1'h0:1'h0];
  assign T10152 = T8251[1'h1:1'h1];
  assign T10153 = T8251[2'h2:2'h2];
  assign T10154 = T8251[2'h3:2'h3];
  assign T10155 = T8251[3'h4:3'h4];
  assign T10156 = T8251[3'h5:3'h5];
  assign T10157 = T10282 ? T10220 : T10158;
  assign T10158 = T10219 ? T10189 : T10159;
  assign T10159 = T10188 ? T10174 : T10160;
  assign T10160 = T10173 ? T10167 : T10161;
  assign T10161 = T10166 ? T10164 : T10162;
  assign T10162 = T10163 ? counts_961 : counts_960;
  assign T10163 = T8251[1'h0:1'h0];
  assign T10164 = T10165 ? counts_963 : counts_962;
  assign T10165 = T8251[1'h0:1'h0];
  assign T10166 = T8251[1'h1:1'h1];
  assign T10167 = T10172 ? T10170 : T10168;
  assign T10168 = T10169 ? counts_965 : counts_964;
  assign T10169 = T8251[1'h0:1'h0];
  assign T10170 = T10171 ? counts_967 : counts_966;
  assign T10171 = T8251[1'h0:1'h0];
  assign T10172 = T8251[1'h1:1'h1];
  assign T10173 = T8251[2'h2:2'h2];
  assign T10174 = T10187 ? T10181 : T10175;
  assign T10175 = T10180 ? T10178 : T10176;
  assign T10176 = T10177 ? counts_969 : counts_968;
  assign T10177 = T8251[1'h0:1'h0];
  assign T10178 = T10179 ? counts_971 : counts_970;
  assign T10179 = T8251[1'h0:1'h0];
  assign T10180 = T8251[1'h1:1'h1];
  assign T10181 = T10186 ? T10184 : T10182;
  assign T10182 = T10183 ? counts_973 : counts_972;
  assign T10183 = T8251[1'h0:1'h0];
  assign T10184 = T10185 ? counts_975 : counts_974;
  assign T10185 = T8251[1'h0:1'h0];
  assign T10186 = T8251[1'h1:1'h1];
  assign T10187 = T8251[2'h2:2'h2];
  assign T10188 = T8251[2'h3:2'h3];
  assign T10189 = T10218 ? T10204 : T10190;
  assign T10190 = T10203 ? T10197 : T10191;
  assign T10191 = T10196 ? T10194 : T10192;
  assign T10192 = T10193 ? counts_977 : counts_976;
  assign T10193 = T8251[1'h0:1'h0];
  assign T10194 = T10195 ? counts_979 : counts_978;
  assign T10195 = T8251[1'h0:1'h0];
  assign T10196 = T8251[1'h1:1'h1];
  assign T10197 = T10202 ? T10200 : T10198;
  assign T10198 = T10199 ? counts_981 : counts_980;
  assign T10199 = T8251[1'h0:1'h0];
  assign T10200 = T10201 ? counts_983 : counts_982;
  assign T10201 = T8251[1'h0:1'h0];
  assign T10202 = T8251[1'h1:1'h1];
  assign T10203 = T8251[2'h2:2'h2];
  assign T10204 = T10217 ? T10211 : T10205;
  assign T10205 = T10210 ? T10208 : T10206;
  assign T10206 = T10207 ? counts_985 : counts_984;
  assign T10207 = T8251[1'h0:1'h0];
  assign T10208 = T10209 ? counts_987 : counts_986;
  assign T10209 = T8251[1'h0:1'h0];
  assign T10210 = T8251[1'h1:1'h1];
  assign T10211 = T10216 ? T10214 : T10212;
  assign T10212 = T10213 ? counts_989 : counts_988;
  assign T10213 = T8251[1'h0:1'h0];
  assign T10214 = T10215 ? counts_991 : counts_990;
  assign T10215 = T8251[1'h0:1'h0];
  assign T10216 = T8251[1'h1:1'h1];
  assign T10217 = T8251[2'h2:2'h2];
  assign T10218 = T8251[2'h3:2'h3];
  assign T10219 = T8251[3'h4:3'h4];
  assign T10220 = T10281 ? T10251 : T10221;
  assign T10221 = T10250 ? T10236 : T10222;
  assign T10222 = T10235 ? T10229 : T10223;
  assign T10223 = T10228 ? T10226 : T10224;
  assign T10224 = T10225 ? counts_993 : counts_992;
  assign T10225 = T8251[1'h0:1'h0];
  assign T10226 = T10227 ? counts_995 : counts_994;
  assign T10227 = T8251[1'h0:1'h0];
  assign T10228 = T8251[1'h1:1'h1];
  assign T10229 = T10234 ? T10232 : T10230;
  assign T10230 = T10231 ? counts_997 : counts_996;
  assign T10231 = T8251[1'h0:1'h0];
  assign T10232 = T10233 ? counts_999 : counts_998;
  assign T10233 = T8251[1'h0:1'h0];
  assign T10234 = T8251[1'h1:1'h1];
  assign T10235 = T8251[2'h2:2'h2];
  assign T10236 = T10249 ? T10243 : T10237;
  assign T10237 = T10242 ? T10240 : T10238;
  assign T10238 = T10239 ? counts_1001 : counts_1000;
  assign T10239 = T8251[1'h0:1'h0];
  assign T10240 = T10241 ? counts_1003 : counts_1002;
  assign T10241 = T8251[1'h0:1'h0];
  assign T10242 = T8251[1'h1:1'h1];
  assign T10243 = T10248 ? T10246 : T10244;
  assign T10244 = T10245 ? counts_1005 : counts_1004;
  assign T10245 = T8251[1'h0:1'h0];
  assign T10246 = T10247 ? counts_1007 : counts_1006;
  assign T10247 = T8251[1'h0:1'h0];
  assign T10248 = T8251[1'h1:1'h1];
  assign T10249 = T8251[2'h2:2'h2];
  assign T10250 = T8251[2'h3:2'h3];
  assign T10251 = T10280 ? T10266 : T10252;
  assign T10252 = T10265 ? T10259 : T10253;
  assign T10253 = T10258 ? T10256 : T10254;
  assign T10254 = T10255 ? counts_1009 : counts_1008;
  assign T10255 = T8251[1'h0:1'h0];
  assign T10256 = T10257 ? counts_1011 : counts_1010;
  assign T10257 = T8251[1'h0:1'h0];
  assign T10258 = T8251[1'h1:1'h1];
  assign T10259 = T10264 ? T10262 : T10260;
  assign T10260 = T10261 ? counts_1013 : counts_1012;
  assign T10261 = T8251[1'h0:1'h0];
  assign T10262 = T10263 ? counts_1015 : counts_1014;
  assign T10263 = T8251[1'h0:1'h0];
  assign T10264 = T8251[1'h1:1'h1];
  assign T10265 = T8251[2'h2:2'h2];
  assign T10266 = T10279 ? T10273 : T10267;
  assign T10267 = T10272 ? T10270 : T10268;
  assign T10268 = T10269 ? counts_1017 : counts_1016;
  assign T10269 = T8251[1'h0:1'h0];
  assign T10270 = T10271 ? counts_1019 : counts_1018;
  assign T10271 = T8251[1'h0:1'h0];
  assign T10272 = T8251[1'h1:1'h1];
  assign T10273 = T10278 ? T10276 : T10274;
  assign T10274 = T10275 ? counts_1021 : counts_1020;
  assign T10275 = T8251[1'h0:1'h0];
  assign T10276 = T10277 ? counts_1023 : counts_1022;
  assign T10277 = T8251[1'h0:1'h0];
  assign T10278 = T8251[1'h1:1'h1];
  assign T10279 = T8251[2'h2:2'h2];
  assign T10280 = T8251[2'h3:2'h3];
  assign T10281 = T8251[3'h4:3'h4];
  assign T10282 = T8251[3'h5:3'h5];
  assign T10283 = T8251[3'h6:3'h6];
  assign T10284 = T8251[3'h7:3'h7];
  assign T10285 = T8251[4'h8:4'h8];
  assign T10286 = T8251[4'h9:4'h9];
  assign T10287 = T10316 & T10288;
  assign T10288 = T38 ^ 1'h1;
  assign T10289 = T10290 ^ 1'h1;
  assign T10290 = T27 | T24;
  assign T10291 = T29 & T10292;
  assign T10292 = T10293 & io_findAvailable;
  assign T10293 = T10294 ^ 1'h1;
  assign T10294 = T10290 | checkFirst;
  assign T10295 = T29 & T10296;
  assign T10296 = T10297 ^ 1'h1;
  assign T10297 = T10294 | io_findAvailable;
  assign T10298 = T10305 & T10299;
  assign T10299 = delayCount == 1'h0;
  assign T10300 = T10303 ? T10302 : T10301;
  assign T10301 = T22 ? 1'h1 : delayCount;
  assign T10302 = delayCount - 1'h1;
  assign T10303 = T10305 & T10304;
  assign T10304 = T10299 ^ 1'h1;
  assign T10305 = 3'h3 == state;
  assign T10306 = T10307 & checkFirst;
  assign T10307 = T10309 & T10308;
  assign T10308 = io_curKeyData != io_allKeyData;
  assign T10309 = 3'h4 == state;
  assign T10310 = T10307 & T10311;
  assign T10311 = T10312 & io_findAvailable;
  assign T10312 = checkFirst ^ 1'h1;
  assign T10313 = T10307 & T10314;
  assign T10314 = T10315 ^ 1'h1;
  assign T10315 = checkFirst | io_findAvailable;
  assign T10316 = 3'h5 == state;
  assign T10317 = T10318 & io_hashOut_ready;
  assign T10318 = 3'h7 == state;
  assign T10319 = T29 & T27;
  assign T10320 = T10309 & T10321;
  assign T10321 = T10336 & reachedEnd;
  assign reachedEnd = T10334 ? T10332 : T10322;
  assign T10322 = delayedIndex == wordLen;
  assign wordLen = curInfo_len[3'h7:2'h2];
  assign T10324 = T10329 ? T10328 : T10325;
  assign T10325 = T10303 ? T10327 : T10326;
  assign T10326 = T22 ? 6'h0 : index;
  assign T10327 = index + 6'h1;
  assign T10328 = index + 6'h1;
  assign T10329 = T10309 & T10330;
  assign T10330 = T10331 ^ 1'h1;
  assign T10331 = T10308 | reachedEnd;
  assign T10332 = delayedIndex == T10333;
  assign T10333 = wordLen - 6'h1;
  assign T10334 = T10335 == 2'h0;
  assign T10335 = curInfo_len[1'h1:1'h0];
  assign T10336 = T10308 ^ 1'h1;
  assign T10337 = curCount < curInfo_tag;
  assign T10338 = T20 ? io_hashIn_bits_tag : curInfo_tag;
  assign curCount = checkFirst ? hashCount1 : hashCount2;
  assign T10339 = 3'h6 == state;
  assign io_hashOut_bits_hash = curHash;
  assign io_hashOut_bits_tag = curInfo_tag;
  assign io_hashOut_valid = T10340;
  assign T10340 = state == 3'h7;
  assign io_hashIn_ready = T10341;
  assign T10341 = state == 3'h0;
  assign io_lenAddr = curHash;
  assign io_allKeyAddr = T10342;
  assign T10342 = {curHash, index};
  assign io_curKeyAddr = index;

  always @(posedge clk) begin
    if(T10339) begin
      hashFound <= T10337;
    end else if(T10320) begin
      hashFound <= 1'h1;
    end else if(T10319) begin
      hashFound <= 1'h1;
    end else if(T4) begin
      hashFound <= 1'h0;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T10317) begin
      state <= 3'h0;
    end else if(T10339) begin
      state <= 3'h7;
    end else if(T10316) begin
      state <= 3'h6;
    end else if(T10320) begin
      state <= 3'h7;
    end else if(T10313) begin
      state <= 3'h7;
    end else if(T10310) begin
      state <= 3'h5;
    end else if(T10306) begin
      state <= 3'h1;
    end else if(T10298) begin
      state <= 3'h4;
    end else if(T10295) begin
      state <= 3'h7;
    end else if(T10291) begin
      state <= 3'h5;
    end else if(T30) begin
      state <= 3'h1;
    end else if(T22) begin
      state <= 3'h3;
    end else if(T10319) begin
      state <= 3'h7;
    end else if(T21) begin
      state <= 3'h2;
    end else if(T20) begin
      state <= 3'h1;
    end
    if(T20) begin
      curInfo_len <= io_hashIn_bits_len;
    end
    if(T10287) begin
      checkFirst <= 1'h0;
    end else if(T37) begin
      checkFirst <= 1'h1;
    end else if(T10306) begin
      checkFirst <= 1'h0;
    end else if(T30) begin
      checkFirst <= 1'h0;
    end else if(T4) begin
      checkFirst <= 1'h1;
    end
    if(reset) begin
      hashCount2 <= 4'h0;
    end else if(T21) begin
      hashCount2 <= T40;
    end
    if(reset) begin
      counts_0 <= 4'h0;
    end else if(T6196) begin
      counts_0 <= T52;
    end else if(io_resetCounts) begin
      counts_0 <= 4'h0;
    end
    if(T20) begin
      curInfo_hash2 <= io_hashIn_bits_hash2;
    end
    if(T20) begin
      curInfo_hash1 <= io_hashIn_bits_hash1;
    end
    if(reset) begin
      counts_2 <= 4'h0;
    end else if(T74) begin
      counts_2 <= T52;
    end else if(io_resetCounts) begin
      counts_2 <= 4'h0;
    end
    if(reset) begin
      counts_3 <= 4'h0;
    end else if(T79) begin
      counts_3 <= T52;
    end else if(io_resetCounts) begin
      counts_3 <= 4'h0;
    end
    if(reset) begin
      counts_4 <= 4'h0;
    end else if(T87) begin
      counts_4 <= T52;
    end else if(io_resetCounts) begin
      counts_4 <= 4'h0;
    end
    if(reset) begin
      counts_5 <= 4'h0;
    end else if(T91) begin
      counts_5 <= T52;
    end else if(io_resetCounts) begin
      counts_5 <= 4'h0;
    end
    if(reset) begin
      counts_6 <= 4'h0;
    end else if(T97) begin
      counts_6 <= T52;
    end else if(io_resetCounts) begin
      counts_6 <= 4'h0;
    end
    if(reset) begin
      counts_7 <= 4'h0;
    end else if(T101) begin
      counts_7 <= T52;
    end else if(io_resetCounts) begin
      counts_7 <= 4'h0;
    end
    if(reset) begin
      counts_8 <= 4'h0;
    end else if(T111) begin
      counts_8 <= T52;
    end else if(io_resetCounts) begin
      counts_8 <= 4'h0;
    end
    if(reset) begin
      counts_9 <= 4'h0;
    end else if(T115) begin
      counts_9 <= T52;
    end else if(io_resetCounts) begin
      counts_9 <= 4'h0;
    end
    if(reset) begin
      counts_10 <= 4'h0;
    end else if(T121) begin
      counts_10 <= T52;
    end else if(io_resetCounts) begin
      counts_10 <= 4'h0;
    end
    if(reset) begin
      counts_11 <= 4'h0;
    end else if(T125) begin
      counts_11 <= T52;
    end else if(io_resetCounts) begin
      counts_11 <= 4'h0;
    end
    if(reset) begin
      counts_12 <= 4'h0;
    end else if(T133) begin
      counts_12 <= T52;
    end else if(io_resetCounts) begin
      counts_12 <= 4'h0;
    end
    if(reset) begin
      counts_13 <= 4'h0;
    end else if(T137) begin
      counts_13 <= T52;
    end else if(io_resetCounts) begin
      counts_13 <= 4'h0;
    end
    if(reset) begin
      counts_14 <= 4'h0;
    end else if(T143) begin
      counts_14 <= T52;
    end else if(io_resetCounts) begin
      counts_14 <= 4'h0;
    end
    if(reset) begin
      counts_15 <= 4'h0;
    end else if(T147) begin
      counts_15 <= T52;
    end else if(io_resetCounts) begin
      counts_15 <= 4'h0;
    end
    if(reset) begin
      counts_16 <= 4'h0;
    end else if(T159) begin
      counts_16 <= T52;
    end else if(io_resetCounts) begin
      counts_16 <= 4'h0;
    end
    if(reset) begin
      counts_17 <= 4'h0;
    end else if(T163) begin
      counts_17 <= T52;
    end else if(io_resetCounts) begin
      counts_17 <= 4'h0;
    end
    if(reset) begin
      counts_18 <= 4'h0;
    end else if(T169) begin
      counts_18 <= T52;
    end else if(io_resetCounts) begin
      counts_18 <= 4'h0;
    end
    if(reset) begin
      counts_19 <= 4'h0;
    end else if(T173) begin
      counts_19 <= T52;
    end else if(io_resetCounts) begin
      counts_19 <= 4'h0;
    end
    if(reset) begin
      counts_20 <= 4'h0;
    end else if(T181) begin
      counts_20 <= T52;
    end else if(io_resetCounts) begin
      counts_20 <= 4'h0;
    end
    if(reset) begin
      counts_21 <= 4'h0;
    end else if(T185) begin
      counts_21 <= T52;
    end else if(io_resetCounts) begin
      counts_21 <= 4'h0;
    end
    if(reset) begin
      counts_22 <= 4'h0;
    end else if(T191) begin
      counts_22 <= T52;
    end else if(io_resetCounts) begin
      counts_22 <= 4'h0;
    end
    if(reset) begin
      counts_23 <= 4'h0;
    end else if(T195) begin
      counts_23 <= T52;
    end else if(io_resetCounts) begin
      counts_23 <= 4'h0;
    end
    if(reset) begin
      counts_24 <= 4'h0;
    end else if(T205) begin
      counts_24 <= T52;
    end else if(io_resetCounts) begin
      counts_24 <= 4'h0;
    end
    if(reset) begin
      counts_25 <= 4'h0;
    end else if(T209) begin
      counts_25 <= T52;
    end else if(io_resetCounts) begin
      counts_25 <= 4'h0;
    end
    if(reset) begin
      counts_26 <= 4'h0;
    end else if(T215) begin
      counts_26 <= T52;
    end else if(io_resetCounts) begin
      counts_26 <= 4'h0;
    end
    if(reset) begin
      counts_27 <= 4'h0;
    end else if(T219) begin
      counts_27 <= T52;
    end else if(io_resetCounts) begin
      counts_27 <= 4'h0;
    end
    if(reset) begin
      counts_28 <= 4'h0;
    end else if(T227) begin
      counts_28 <= T52;
    end else if(io_resetCounts) begin
      counts_28 <= 4'h0;
    end
    if(reset) begin
      counts_29 <= 4'h0;
    end else if(T231) begin
      counts_29 <= T52;
    end else if(io_resetCounts) begin
      counts_29 <= 4'h0;
    end
    if(reset) begin
      counts_30 <= 4'h0;
    end else if(T237) begin
      counts_30 <= T52;
    end else if(io_resetCounts) begin
      counts_30 <= 4'h0;
    end
    if(reset) begin
      counts_31 <= 4'h0;
    end else if(T241) begin
      counts_31 <= T52;
    end else if(io_resetCounts) begin
      counts_31 <= 4'h0;
    end
    if(reset) begin
      counts_32 <= 4'h0;
    end else if(T255) begin
      counts_32 <= T52;
    end else if(io_resetCounts) begin
      counts_32 <= 4'h0;
    end
    if(reset) begin
      counts_33 <= 4'h0;
    end else if(T259) begin
      counts_33 <= T52;
    end else if(io_resetCounts) begin
      counts_33 <= 4'h0;
    end
    if(reset) begin
      counts_34 <= 4'h0;
    end else if(T265) begin
      counts_34 <= T52;
    end else if(io_resetCounts) begin
      counts_34 <= 4'h0;
    end
    if(reset) begin
      counts_35 <= 4'h0;
    end else if(T269) begin
      counts_35 <= T52;
    end else if(io_resetCounts) begin
      counts_35 <= 4'h0;
    end
    if(reset) begin
      counts_36 <= 4'h0;
    end else if(T277) begin
      counts_36 <= T52;
    end else if(io_resetCounts) begin
      counts_36 <= 4'h0;
    end
    if(reset) begin
      counts_37 <= 4'h0;
    end else if(T281) begin
      counts_37 <= T52;
    end else if(io_resetCounts) begin
      counts_37 <= 4'h0;
    end
    if(reset) begin
      counts_38 <= 4'h0;
    end else if(T287) begin
      counts_38 <= T52;
    end else if(io_resetCounts) begin
      counts_38 <= 4'h0;
    end
    if(reset) begin
      counts_39 <= 4'h0;
    end else if(T291) begin
      counts_39 <= T52;
    end else if(io_resetCounts) begin
      counts_39 <= 4'h0;
    end
    if(reset) begin
      counts_40 <= 4'h0;
    end else if(T301) begin
      counts_40 <= T52;
    end else if(io_resetCounts) begin
      counts_40 <= 4'h0;
    end
    if(reset) begin
      counts_41 <= 4'h0;
    end else if(T305) begin
      counts_41 <= T52;
    end else if(io_resetCounts) begin
      counts_41 <= 4'h0;
    end
    if(reset) begin
      counts_42 <= 4'h0;
    end else if(T311) begin
      counts_42 <= T52;
    end else if(io_resetCounts) begin
      counts_42 <= 4'h0;
    end
    if(reset) begin
      counts_43 <= 4'h0;
    end else if(T315) begin
      counts_43 <= T52;
    end else if(io_resetCounts) begin
      counts_43 <= 4'h0;
    end
    if(reset) begin
      counts_44 <= 4'h0;
    end else if(T323) begin
      counts_44 <= T52;
    end else if(io_resetCounts) begin
      counts_44 <= 4'h0;
    end
    if(reset) begin
      counts_45 <= 4'h0;
    end else if(T327) begin
      counts_45 <= T52;
    end else if(io_resetCounts) begin
      counts_45 <= 4'h0;
    end
    if(reset) begin
      counts_46 <= 4'h0;
    end else if(T333) begin
      counts_46 <= T52;
    end else if(io_resetCounts) begin
      counts_46 <= 4'h0;
    end
    if(reset) begin
      counts_47 <= 4'h0;
    end else if(T337) begin
      counts_47 <= T52;
    end else if(io_resetCounts) begin
      counts_47 <= 4'h0;
    end
    if(reset) begin
      counts_48 <= 4'h0;
    end else if(T349) begin
      counts_48 <= T52;
    end else if(io_resetCounts) begin
      counts_48 <= 4'h0;
    end
    if(reset) begin
      counts_49 <= 4'h0;
    end else if(T353) begin
      counts_49 <= T52;
    end else if(io_resetCounts) begin
      counts_49 <= 4'h0;
    end
    if(reset) begin
      counts_50 <= 4'h0;
    end else if(T359) begin
      counts_50 <= T52;
    end else if(io_resetCounts) begin
      counts_50 <= 4'h0;
    end
    if(reset) begin
      counts_51 <= 4'h0;
    end else if(T363) begin
      counts_51 <= T52;
    end else if(io_resetCounts) begin
      counts_51 <= 4'h0;
    end
    if(reset) begin
      counts_52 <= 4'h0;
    end else if(T371) begin
      counts_52 <= T52;
    end else if(io_resetCounts) begin
      counts_52 <= 4'h0;
    end
    if(reset) begin
      counts_53 <= 4'h0;
    end else if(T375) begin
      counts_53 <= T52;
    end else if(io_resetCounts) begin
      counts_53 <= 4'h0;
    end
    if(reset) begin
      counts_54 <= 4'h0;
    end else if(T381) begin
      counts_54 <= T52;
    end else if(io_resetCounts) begin
      counts_54 <= 4'h0;
    end
    if(reset) begin
      counts_55 <= 4'h0;
    end else if(T385) begin
      counts_55 <= T52;
    end else if(io_resetCounts) begin
      counts_55 <= 4'h0;
    end
    if(reset) begin
      counts_56 <= 4'h0;
    end else if(T395) begin
      counts_56 <= T52;
    end else if(io_resetCounts) begin
      counts_56 <= 4'h0;
    end
    if(reset) begin
      counts_57 <= 4'h0;
    end else if(T399) begin
      counts_57 <= T52;
    end else if(io_resetCounts) begin
      counts_57 <= 4'h0;
    end
    if(reset) begin
      counts_58 <= 4'h0;
    end else if(T405) begin
      counts_58 <= T52;
    end else if(io_resetCounts) begin
      counts_58 <= 4'h0;
    end
    if(reset) begin
      counts_59 <= 4'h0;
    end else if(T409) begin
      counts_59 <= T52;
    end else if(io_resetCounts) begin
      counts_59 <= 4'h0;
    end
    if(reset) begin
      counts_60 <= 4'h0;
    end else if(T417) begin
      counts_60 <= T52;
    end else if(io_resetCounts) begin
      counts_60 <= 4'h0;
    end
    if(reset) begin
      counts_61 <= 4'h0;
    end else if(T421) begin
      counts_61 <= T52;
    end else if(io_resetCounts) begin
      counts_61 <= 4'h0;
    end
    if(reset) begin
      counts_62 <= 4'h0;
    end else if(T427) begin
      counts_62 <= T52;
    end else if(io_resetCounts) begin
      counts_62 <= 4'h0;
    end
    if(reset) begin
      counts_63 <= 4'h0;
    end else if(T431) begin
      counts_63 <= T52;
    end else if(io_resetCounts) begin
      counts_63 <= 4'h0;
    end
    if(reset) begin
      counts_64 <= 4'h0;
    end else if(T447) begin
      counts_64 <= T52;
    end else if(io_resetCounts) begin
      counts_64 <= 4'h0;
    end
    if(reset) begin
      counts_65 <= 4'h0;
    end else if(T451) begin
      counts_65 <= T52;
    end else if(io_resetCounts) begin
      counts_65 <= 4'h0;
    end
    if(reset) begin
      counts_66 <= 4'h0;
    end else if(T457) begin
      counts_66 <= T52;
    end else if(io_resetCounts) begin
      counts_66 <= 4'h0;
    end
    if(reset) begin
      counts_67 <= 4'h0;
    end else if(T461) begin
      counts_67 <= T52;
    end else if(io_resetCounts) begin
      counts_67 <= 4'h0;
    end
    if(reset) begin
      counts_68 <= 4'h0;
    end else if(T469) begin
      counts_68 <= T52;
    end else if(io_resetCounts) begin
      counts_68 <= 4'h0;
    end
    if(reset) begin
      counts_69 <= 4'h0;
    end else if(T473) begin
      counts_69 <= T52;
    end else if(io_resetCounts) begin
      counts_69 <= 4'h0;
    end
    if(reset) begin
      counts_70 <= 4'h0;
    end else if(T479) begin
      counts_70 <= T52;
    end else if(io_resetCounts) begin
      counts_70 <= 4'h0;
    end
    if(reset) begin
      counts_71 <= 4'h0;
    end else if(T483) begin
      counts_71 <= T52;
    end else if(io_resetCounts) begin
      counts_71 <= 4'h0;
    end
    if(reset) begin
      counts_72 <= 4'h0;
    end else if(T493) begin
      counts_72 <= T52;
    end else if(io_resetCounts) begin
      counts_72 <= 4'h0;
    end
    if(reset) begin
      counts_73 <= 4'h0;
    end else if(T497) begin
      counts_73 <= T52;
    end else if(io_resetCounts) begin
      counts_73 <= 4'h0;
    end
    if(reset) begin
      counts_74 <= 4'h0;
    end else if(T503) begin
      counts_74 <= T52;
    end else if(io_resetCounts) begin
      counts_74 <= 4'h0;
    end
    if(reset) begin
      counts_75 <= 4'h0;
    end else if(T507) begin
      counts_75 <= T52;
    end else if(io_resetCounts) begin
      counts_75 <= 4'h0;
    end
    if(reset) begin
      counts_76 <= 4'h0;
    end else if(T515) begin
      counts_76 <= T52;
    end else if(io_resetCounts) begin
      counts_76 <= 4'h0;
    end
    if(reset) begin
      counts_77 <= 4'h0;
    end else if(T519) begin
      counts_77 <= T52;
    end else if(io_resetCounts) begin
      counts_77 <= 4'h0;
    end
    if(reset) begin
      counts_78 <= 4'h0;
    end else if(T525) begin
      counts_78 <= T52;
    end else if(io_resetCounts) begin
      counts_78 <= 4'h0;
    end
    if(reset) begin
      counts_79 <= 4'h0;
    end else if(T529) begin
      counts_79 <= T52;
    end else if(io_resetCounts) begin
      counts_79 <= 4'h0;
    end
    if(reset) begin
      counts_80 <= 4'h0;
    end else if(T541) begin
      counts_80 <= T52;
    end else if(io_resetCounts) begin
      counts_80 <= 4'h0;
    end
    if(reset) begin
      counts_81 <= 4'h0;
    end else if(T545) begin
      counts_81 <= T52;
    end else if(io_resetCounts) begin
      counts_81 <= 4'h0;
    end
    if(reset) begin
      counts_82 <= 4'h0;
    end else if(T551) begin
      counts_82 <= T52;
    end else if(io_resetCounts) begin
      counts_82 <= 4'h0;
    end
    if(reset) begin
      counts_83 <= 4'h0;
    end else if(T555) begin
      counts_83 <= T52;
    end else if(io_resetCounts) begin
      counts_83 <= 4'h0;
    end
    if(reset) begin
      counts_84 <= 4'h0;
    end else if(T563) begin
      counts_84 <= T52;
    end else if(io_resetCounts) begin
      counts_84 <= 4'h0;
    end
    if(reset) begin
      counts_85 <= 4'h0;
    end else if(T567) begin
      counts_85 <= T52;
    end else if(io_resetCounts) begin
      counts_85 <= 4'h0;
    end
    if(reset) begin
      counts_86 <= 4'h0;
    end else if(T573) begin
      counts_86 <= T52;
    end else if(io_resetCounts) begin
      counts_86 <= 4'h0;
    end
    if(reset) begin
      counts_87 <= 4'h0;
    end else if(T577) begin
      counts_87 <= T52;
    end else if(io_resetCounts) begin
      counts_87 <= 4'h0;
    end
    if(reset) begin
      counts_88 <= 4'h0;
    end else if(T587) begin
      counts_88 <= T52;
    end else if(io_resetCounts) begin
      counts_88 <= 4'h0;
    end
    if(reset) begin
      counts_89 <= 4'h0;
    end else if(T591) begin
      counts_89 <= T52;
    end else if(io_resetCounts) begin
      counts_89 <= 4'h0;
    end
    if(reset) begin
      counts_90 <= 4'h0;
    end else if(T597) begin
      counts_90 <= T52;
    end else if(io_resetCounts) begin
      counts_90 <= 4'h0;
    end
    if(reset) begin
      counts_91 <= 4'h0;
    end else if(T601) begin
      counts_91 <= T52;
    end else if(io_resetCounts) begin
      counts_91 <= 4'h0;
    end
    if(reset) begin
      counts_92 <= 4'h0;
    end else if(T609) begin
      counts_92 <= T52;
    end else if(io_resetCounts) begin
      counts_92 <= 4'h0;
    end
    if(reset) begin
      counts_93 <= 4'h0;
    end else if(T613) begin
      counts_93 <= T52;
    end else if(io_resetCounts) begin
      counts_93 <= 4'h0;
    end
    if(reset) begin
      counts_94 <= 4'h0;
    end else if(T619) begin
      counts_94 <= T52;
    end else if(io_resetCounts) begin
      counts_94 <= 4'h0;
    end
    if(reset) begin
      counts_95 <= 4'h0;
    end else if(T623) begin
      counts_95 <= T52;
    end else if(io_resetCounts) begin
      counts_95 <= 4'h0;
    end
    if(reset) begin
      counts_96 <= 4'h0;
    end else if(T637) begin
      counts_96 <= T52;
    end else if(io_resetCounts) begin
      counts_96 <= 4'h0;
    end
    if(reset) begin
      counts_97 <= 4'h0;
    end else if(T641) begin
      counts_97 <= T52;
    end else if(io_resetCounts) begin
      counts_97 <= 4'h0;
    end
    if(reset) begin
      counts_98 <= 4'h0;
    end else if(T647) begin
      counts_98 <= T52;
    end else if(io_resetCounts) begin
      counts_98 <= 4'h0;
    end
    if(reset) begin
      counts_99 <= 4'h0;
    end else if(T651) begin
      counts_99 <= T52;
    end else if(io_resetCounts) begin
      counts_99 <= 4'h0;
    end
    if(reset) begin
      counts_100 <= 4'h0;
    end else if(T659) begin
      counts_100 <= T52;
    end else if(io_resetCounts) begin
      counts_100 <= 4'h0;
    end
    if(reset) begin
      counts_101 <= 4'h0;
    end else if(T663) begin
      counts_101 <= T52;
    end else if(io_resetCounts) begin
      counts_101 <= 4'h0;
    end
    if(reset) begin
      counts_102 <= 4'h0;
    end else if(T669) begin
      counts_102 <= T52;
    end else if(io_resetCounts) begin
      counts_102 <= 4'h0;
    end
    if(reset) begin
      counts_103 <= 4'h0;
    end else if(T673) begin
      counts_103 <= T52;
    end else if(io_resetCounts) begin
      counts_103 <= 4'h0;
    end
    if(reset) begin
      counts_104 <= 4'h0;
    end else if(T683) begin
      counts_104 <= T52;
    end else if(io_resetCounts) begin
      counts_104 <= 4'h0;
    end
    if(reset) begin
      counts_105 <= 4'h0;
    end else if(T687) begin
      counts_105 <= T52;
    end else if(io_resetCounts) begin
      counts_105 <= 4'h0;
    end
    if(reset) begin
      counts_106 <= 4'h0;
    end else if(T693) begin
      counts_106 <= T52;
    end else if(io_resetCounts) begin
      counts_106 <= 4'h0;
    end
    if(reset) begin
      counts_107 <= 4'h0;
    end else if(T697) begin
      counts_107 <= T52;
    end else if(io_resetCounts) begin
      counts_107 <= 4'h0;
    end
    if(reset) begin
      counts_108 <= 4'h0;
    end else if(T705) begin
      counts_108 <= T52;
    end else if(io_resetCounts) begin
      counts_108 <= 4'h0;
    end
    if(reset) begin
      counts_109 <= 4'h0;
    end else if(T709) begin
      counts_109 <= T52;
    end else if(io_resetCounts) begin
      counts_109 <= 4'h0;
    end
    if(reset) begin
      counts_110 <= 4'h0;
    end else if(T715) begin
      counts_110 <= T52;
    end else if(io_resetCounts) begin
      counts_110 <= 4'h0;
    end
    if(reset) begin
      counts_111 <= 4'h0;
    end else if(T719) begin
      counts_111 <= T52;
    end else if(io_resetCounts) begin
      counts_111 <= 4'h0;
    end
    if(reset) begin
      counts_112 <= 4'h0;
    end else if(T731) begin
      counts_112 <= T52;
    end else if(io_resetCounts) begin
      counts_112 <= 4'h0;
    end
    if(reset) begin
      counts_113 <= 4'h0;
    end else if(T735) begin
      counts_113 <= T52;
    end else if(io_resetCounts) begin
      counts_113 <= 4'h0;
    end
    if(reset) begin
      counts_114 <= 4'h0;
    end else if(T741) begin
      counts_114 <= T52;
    end else if(io_resetCounts) begin
      counts_114 <= 4'h0;
    end
    if(reset) begin
      counts_115 <= 4'h0;
    end else if(T745) begin
      counts_115 <= T52;
    end else if(io_resetCounts) begin
      counts_115 <= 4'h0;
    end
    if(reset) begin
      counts_116 <= 4'h0;
    end else if(T753) begin
      counts_116 <= T52;
    end else if(io_resetCounts) begin
      counts_116 <= 4'h0;
    end
    if(reset) begin
      counts_117 <= 4'h0;
    end else if(T757) begin
      counts_117 <= T52;
    end else if(io_resetCounts) begin
      counts_117 <= 4'h0;
    end
    if(reset) begin
      counts_118 <= 4'h0;
    end else if(T763) begin
      counts_118 <= T52;
    end else if(io_resetCounts) begin
      counts_118 <= 4'h0;
    end
    if(reset) begin
      counts_119 <= 4'h0;
    end else if(T767) begin
      counts_119 <= T52;
    end else if(io_resetCounts) begin
      counts_119 <= 4'h0;
    end
    if(reset) begin
      counts_120 <= 4'h0;
    end else if(T777) begin
      counts_120 <= T52;
    end else if(io_resetCounts) begin
      counts_120 <= 4'h0;
    end
    if(reset) begin
      counts_121 <= 4'h0;
    end else if(T781) begin
      counts_121 <= T52;
    end else if(io_resetCounts) begin
      counts_121 <= 4'h0;
    end
    if(reset) begin
      counts_122 <= 4'h0;
    end else if(T787) begin
      counts_122 <= T52;
    end else if(io_resetCounts) begin
      counts_122 <= 4'h0;
    end
    if(reset) begin
      counts_123 <= 4'h0;
    end else if(T791) begin
      counts_123 <= T52;
    end else if(io_resetCounts) begin
      counts_123 <= 4'h0;
    end
    if(reset) begin
      counts_124 <= 4'h0;
    end else if(T799) begin
      counts_124 <= T52;
    end else if(io_resetCounts) begin
      counts_124 <= 4'h0;
    end
    if(reset) begin
      counts_125 <= 4'h0;
    end else if(T803) begin
      counts_125 <= T52;
    end else if(io_resetCounts) begin
      counts_125 <= 4'h0;
    end
    if(reset) begin
      counts_126 <= 4'h0;
    end else if(T809) begin
      counts_126 <= T52;
    end else if(io_resetCounts) begin
      counts_126 <= 4'h0;
    end
    if(reset) begin
      counts_127 <= 4'h0;
    end else if(T813) begin
      counts_127 <= T52;
    end else if(io_resetCounts) begin
      counts_127 <= 4'h0;
    end
    if(reset) begin
      counts_128 <= 4'h0;
    end else if(T831) begin
      counts_128 <= T52;
    end else if(io_resetCounts) begin
      counts_128 <= 4'h0;
    end
    if(reset) begin
      counts_129 <= 4'h0;
    end else if(T835) begin
      counts_129 <= T52;
    end else if(io_resetCounts) begin
      counts_129 <= 4'h0;
    end
    if(reset) begin
      counts_130 <= 4'h0;
    end else if(T841) begin
      counts_130 <= T52;
    end else if(io_resetCounts) begin
      counts_130 <= 4'h0;
    end
    if(reset) begin
      counts_131 <= 4'h0;
    end else if(T845) begin
      counts_131 <= T52;
    end else if(io_resetCounts) begin
      counts_131 <= 4'h0;
    end
    if(reset) begin
      counts_132 <= 4'h0;
    end else if(T853) begin
      counts_132 <= T52;
    end else if(io_resetCounts) begin
      counts_132 <= 4'h0;
    end
    if(reset) begin
      counts_133 <= 4'h0;
    end else if(T857) begin
      counts_133 <= T52;
    end else if(io_resetCounts) begin
      counts_133 <= 4'h0;
    end
    if(reset) begin
      counts_134 <= 4'h0;
    end else if(T863) begin
      counts_134 <= T52;
    end else if(io_resetCounts) begin
      counts_134 <= 4'h0;
    end
    if(reset) begin
      counts_135 <= 4'h0;
    end else if(T867) begin
      counts_135 <= T52;
    end else if(io_resetCounts) begin
      counts_135 <= 4'h0;
    end
    if(reset) begin
      counts_136 <= 4'h0;
    end else if(T877) begin
      counts_136 <= T52;
    end else if(io_resetCounts) begin
      counts_136 <= 4'h0;
    end
    if(reset) begin
      counts_137 <= 4'h0;
    end else if(T881) begin
      counts_137 <= T52;
    end else if(io_resetCounts) begin
      counts_137 <= 4'h0;
    end
    if(reset) begin
      counts_138 <= 4'h0;
    end else if(T887) begin
      counts_138 <= T52;
    end else if(io_resetCounts) begin
      counts_138 <= 4'h0;
    end
    if(reset) begin
      counts_139 <= 4'h0;
    end else if(T891) begin
      counts_139 <= T52;
    end else if(io_resetCounts) begin
      counts_139 <= 4'h0;
    end
    if(reset) begin
      counts_140 <= 4'h0;
    end else if(T899) begin
      counts_140 <= T52;
    end else if(io_resetCounts) begin
      counts_140 <= 4'h0;
    end
    if(reset) begin
      counts_141 <= 4'h0;
    end else if(T903) begin
      counts_141 <= T52;
    end else if(io_resetCounts) begin
      counts_141 <= 4'h0;
    end
    if(reset) begin
      counts_142 <= 4'h0;
    end else if(T909) begin
      counts_142 <= T52;
    end else if(io_resetCounts) begin
      counts_142 <= 4'h0;
    end
    if(reset) begin
      counts_143 <= 4'h0;
    end else if(T913) begin
      counts_143 <= T52;
    end else if(io_resetCounts) begin
      counts_143 <= 4'h0;
    end
    if(reset) begin
      counts_144 <= 4'h0;
    end else if(T925) begin
      counts_144 <= T52;
    end else if(io_resetCounts) begin
      counts_144 <= 4'h0;
    end
    if(reset) begin
      counts_145 <= 4'h0;
    end else if(T929) begin
      counts_145 <= T52;
    end else if(io_resetCounts) begin
      counts_145 <= 4'h0;
    end
    if(reset) begin
      counts_146 <= 4'h0;
    end else if(T935) begin
      counts_146 <= T52;
    end else if(io_resetCounts) begin
      counts_146 <= 4'h0;
    end
    if(reset) begin
      counts_147 <= 4'h0;
    end else if(T939) begin
      counts_147 <= T52;
    end else if(io_resetCounts) begin
      counts_147 <= 4'h0;
    end
    if(reset) begin
      counts_148 <= 4'h0;
    end else if(T947) begin
      counts_148 <= T52;
    end else if(io_resetCounts) begin
      counts_148 <= 4'h0;
    end
    if(reset) begin
      counts_149 <= 4'h0;
    end else if(T951) begin
      counts_149 <= T52;
    end else if(io_resetCounts) begin
      counts_149 <= 4'h0;
    end
    if(reset) begin
      counts_150 <= 4'h0;
    end else if(T957) begin
      counts_150 <= T52;
    end else if(io_resetCounts) begin
      counts_150 <= 4'h0;
    end
    if(reset) begin
      counts_151 <= 4'h0;
    end else if(T961) begin
      counts_151 <= T52;
    end else if(io_resetCounts) begin
      counts_151 <= 4'h0;
    end
    if(reset) begin
      counts_152 <= 4'h0;
    end else if(T971) begin
      counts_152 <= T52;
    end else if(io_resetCounts) begin
      counts_152 <= 4'h0;
    end
    if(reset) begin
      counts_153 <= 4'h0;
    end else if(T975) begin
      counts_153 <= T52;
    end else if(io_resetCounts) begin
      counts_153 <= 4'h0;
    end
    if(reset) begin
      counts_154 <= 4'h0;
    end else if(T981) begin
      counts_154 <= T52;
    end else if(io_resetCounts) begin
      counts_154 <= 4'h0;
    end
    if(reset) begin
      counts_155 <= 4'h0;
    end else if(T985) begin
      counts_155 <= T52;
    end else if(io_resetCounts) begin
      counts_155 <= 4'h0;
    end
    if(reset) begin
      counts_156 <= 4'h0;
    end else if(T993) begin
      counts_156 <= T52;
    end else if(io_resetCounts) begin
      counts_156 <= 4'h0;
    end
    if(reset) begin
      counts_157 <= 4'h0;
    end else if(T997) begin
      counts_157 <= T52;
    end else if(io_resetCounts) begin
      counts_157 <= 4'h0;
    end
    if(reset) begin
      counts_158 <= 4'h0;
    end else if(T1003) begin
      counts_158 <= T52;
    end else if(io_resetCounts) begin
      counts_158 <= 4'h0;
    end
    if(reset) begin
      counts_159 <= 4'h0;
    end else if(T1007) begin
      counts_159 <= T52;
    end else if(io_resetCounts) begin
      counts_159 <= 4'h0;
    end
    if(reset) begin
      counts_160 <= 4'h0;
    end else if(T1021) begin
      counts_160 <= T52;
    end else if(io_resetCounts) begin
      counts_160 <= 4'h0;
    end
    if(reset) begin
      counts_161 <= 4'h0;
    end else if(T1025) begin
      counts_161 <= T52;
    end else if(io_resetCounts) begin
      counts_161 <= 4'h0;
    end
    if(reset) begin
      counts_162 <= 4'h0;
    end else if(T1031) begin
      counts_162 <= T52;
    end else if(io_resetCounts) begin
      counts_162 <= 4'h0;
    end
    if(reset) begin
      counts_163 <= 4'h0;
    end else if(T1035) begin
      counts_163 <= T52;
    end else if(io_resetCounts) begin
      counts_163 <= 4'h0;
    end
    if(reset) begin
      counts_164 <= 4'h0;
    end else if(T1043) begin
      counts_164 <= T52;
    end else if(io_resetCounts) begin
      counts_164 <= 4'h0;
    end
    if(reset) begin
      counts_165 <= 4'h0;
    end else if(T1047) begin
      counts_165 <= T52;
    end else if(io_resetCounts) begin
      counts_165 <= 4'h0;
    end
    if(reset) begin
      counts_166 <= 4'h0;
    end else if(T1053) begin
      counts_166 <= T52;
    end else if(io_resetCounts) begin
      counts_166 <= 4'h0;
    end
    if(reset) begin
      counts_167 <= 4'h0;
    end else if(T1057) begin
      counts_167 <= T52;
    end else if(io_resetCounts) begin
      counts_167 <= 4'h0;
    end
    if(reset) begin
      counts_168 <= 4'h0;
    end else if(T1067) begin
      counts_168 <= T52;
    end else if(io_resetCounts) begin
      counts_168 <= 4'h0;
    end
    if(reset) begin
      counts_169 <= 4'h0;
    end else if(T1071) begin
      counts_169 <= T52;
    end else if(io_resetCounts) begin
      counts_169 <= 4'h0;
    end
    if(reset) begin
      counts_170 <= 4'h0;
    end else if(T1077) begin
      counts_170 <= T52;
    end else if(io_resetCounts) begin
      counts_170 <= 4'h0;
    end
    if(reset) begin
      counts_171 <= 4'h0;
    end else if(T1081) begin
      counts_171 <= T52;
    end else if(io_resetCounts) begin
      counts_171 <= 4'h0;
    end
    if(reset) begin
      counts_172 <= 4'h0;
    end else if(T1089) begin
      counts_172 <= T52;
    end else if(io_resetCounts) begin
      counts_172 <= 4'h0;
    end
    if(reset) begin
      counts_173 <= 4'h0;
    end else if(T1093) begin
      counts_173 <= T52;
    end else if(io_resetCounts) begin
      counts_173 <= 4'h0;
    end
    if(reset) begin
      counts_174 <= 4'h0;
    end else if(T1099) begin
      counts_174 <= T52;
    end else if(io_resetCounts) begin
      counts_174 <= 4'h0;
    end
    if(reset) begin
      counts_175 <= 4'h0;
    end else if(T1103) begin
      counts_175 <= T52;
    end else if(io_resetCounts) begin
      counts_175 <= 4'h0;
    end
    if(reset) begin
      counts_176 <= 4'h0;
    end else if(T1115) begin
      counts_176 <= T52;
    end else if(io_resetCounts) begin
      counts_176 <= 4'h0;
    end
    if(reset) begin
      counts_177 <= 4'h0;
    end else if(T1119) begin
      counts_177 <= T52;
    end else if(io_resetCounts) begin
      counts_177 <= 4'h0;
    end
    if(reset) begin
      counts_178 <= 4'h0;
    end else if(T1125) begin
      counts_178 <= T52;
    end else if(io_resetCounts) begin
      counts_178 <= 4'h0;
    end
    if(reset) begin
      counts_179 <= 4'h0;
    end else if(T1129) begin
      counts_179 <= T52;
    end else if(io_resetCounts) begin
      counts_179 <= 4'h0;
    end
    if(reset) begin
      counts_180 <= 4'h0;
    end else if(T1137) begin
      counts_180 <= T52;
    end else if(io_resetCounts) begin
      counts_180 <= 4'h0;
    end
    if(reset) begin
      counts_181 <= 4'h0;
    end else if(T1141) begin
      counts_181 <= T52;
    end else if(io_resetCounts) begin
      counts_181 <= 4'h0;
    end
    if(reset) begin
      counts_182 <= 4'h0;
    end else if(T1147) begin
      counts_182 <= T52;
    end else if(io_resetCounts) begin
      counts_182 <= 4'h0;
    end
    if(reset) begin
      counts_183 <= 4'h0;
    end else if(T1151) begin
      counts_183 <= T52;
    end else if(io_resetCounts) begin
      counts_183 <= 4'h0;
    end
    if(reset) begin
      counts_184 <= 4'h0;
    end else if(T1161) begin
      counts_184 <= T52;
    end else if(io_resetCounts) begin
      counts_184 <= 4'h0;
    end
    if(reset) begin
      counts_185 <= 4'h0;
    end else if(T1165) begin
      counts_185 <= T52;
    end else if(io_resetCounts) begin
      counts_185 <= 4'h0;
    end
    if(reset) begin
      counts_186 <= 4'h0;
    end else if(T1171) begin
      counts_186 <= T52;
    end else if(io_resetCounts) begin
      counts_186 <= 4'h0;
    end
    if(reset) begin
      counts_187 <= 4'h0;
    end else if(T1175) begin
      counts_187 <= T52;
    end else if(io_resetCounts) begin
      counts_187 <= 4'h0;
    end
    if(reset) begin
      counts_188 <= 4'h0;
    end else if(T1183) begin
      counts_188 <= T52;
    end else if(io_resetCounts) begin
      counts_188 <= 4'h0;
    end
    if(reset) begin
      counts_189 <= 4'h0;
    end else if(T1187) begin
      counts_189 <= T52;
    end else if(io_resetCounts) begin
      counts_189 <= 4'h0;
    end
    if(reset) begin
      counts_190 <= 4'h0;
    end else if(T1193) begin
      counts_190 <= T52;
    end else if(io_resetCounts) begin
      counts_190 <= 4'h0;
    end
    if(reset) begin
      counts_191 <= 4'h0;
    end else if(T1197) begin
      counts_191 <= T52;
    end else if(io_resetCounts) begin
      counts_191 <= 4'h0;
    end
    if(reset) begin
      counts_192 <= 4'h0;
    end else if(T1213) begin
      counts_192 <= T52;
    end else if(io_resetCounts) begin
      counts_192 <= 4'h0;
    end
    if(reset) begin
      counts_193 <= 4'h0;
    end else if(T1217) begin
      counts_193 <= T52;
    end else if(io_resetCounts) begin
      counts_193 <= 4'h0;
    end
    if(reset) begin
      counts_194 <= 4'h0;
    end else if(T1223) begin
      counts_194 <= T52;
    end else if(io_resetCounts) begin
      counts_194 <= 4'h0;
    end
    if(reset) begin
      counts_195 <= 4'h0;
    end else if(T1227) begin
      counts_195 <= T52;
    end else if(io_resetCounts) begin
      counts_195 <= 4'h0;
    end
    if(reset) begin
      counts_196 <= 4'h0;
    end else if(T1235) begin
      counts_196 <= T52;
    end else if(io_resetCounts) begin
      counts_196 <= 4'h0;
    end
    if(reset) begin
      counts_197 <= 4'h0;
    end else if(T1239) begin
      counts_197 <= T52;
    end else if(io_resetCounts) begin
      counts_197 <= 4'h0;
    end
    if(reset) begin
      counts_198 <= 4'h0;
    end else if(T1245) begin
      counts_198 <= T52;
    end else if(io_resetCounts) begin
      counts_198 <= 4'h0;
    end
    if(reset) begin
      counts_199 <= 4'h0;
    end else if(T1249) begin
      counts_199 <= T52;
    end else if(io_resetCounts) begin
      counts_199 <= 4'h0;
    end
    if(reset) begin
      counts_200 <= 4'h0;
    end else if(T1259) begin
      counts_200 <= T52;
    end else if(io_resetCounts) begin
      counts_200 <= 4'h0;
    end
    if(reset) begin
      counts_201 <= 4'h0;
    end else if(T1263) begin
      counts_201 <= T52;
    end else if(io_resetCounts) begin
      counts_201 <= 4'h0;
    end
    if(reset) begin
      counts_202 <= 4'h0;
    end else if(T1269) begin
      counts_202 <= T52;
    end else if(io_resetCounts) begin
      counts_202 <= 4'h0;
    end
    if(reset) begin
      counts_203 <= 4'h0;
    end else if(T1273) begin
      counts_203 <= T52;
    end else if(io_resetCounts) begin
      counts_203 <= 4'h0;
    end
    if(reset) begin
      counts_204 <= 4'h0;
    end else if(T1281) begin
      counts_204 <= T52;
    end else if(io_resetCounts) begin
      counts_204 <= 4'h0;
    end
    if(reset) begin
      counts_205 <= 4'h0;
    end else if(T1285) begin
      counts_205 <= T52;
    end else if(io_resetCounts) begin
      counts_205 <= 4'h0;
    end
    if(reset) begin
      counts_206 <= 4'h0;
    end else if(T1291) begin
      counts_206 <= T52;
    end else if(io_resetCounts) begin
      counts_206 <= 4'h0;
    end
    if(reset) begin
      counts_207 <= 4'h0;
    end else if(T1295) begin
      counts_207 <= T52;
    end else if(io_resetCounts) begin
      counts_207 <= 4'h0;
    end
    if(reset) begin
      counts_208 <= 4'h0;
    end else if(T1307) begin
      counts_208 <= T52;
    end else if(io_resetCounts) begin
      counts_208 <= 4'h0;
    end
    if(reset) begin
      counts_209 <= 4'h0;
    end else if(T1311) begin
      counts_209 <= T52;
    end else if(io_resetCounts) begin
      counts_209 <= 4'h0;
    end
    if(reset) begin
      counts_210 <= 4'h0;
    end else if(T1317) begin
      counts_210 <= T52;
    end else if(io_resetCounts) begin
      counts_210 <= 4'h0;
    end
    if(reset) begin
      counts_211 <= 4'h0;
    end else if(T1321) begin
      counts_211 <= T52;
    end else if(io_resetCounts) begin
      counts_211 <= 4'h0;
    end
    if(reset) begin
      counts_212 <= 4'h0;
    end else if(T1329) begin
      counts_212 <= T52;
    end else if(io_resetCounts) begin
      counts_212 <= 4'h0;
    end
    if(reset) begin
      counts_213 <= 4'h0;
    end else if(T1333) begin
      counts_213 <= T52;
    end else if(io_resetCounts) begin
      counts_213 <= 4'h0;
    end
    if(reset) begin
      counts_214 <= 4'h0;
    end else if(T1339) begin
      counts_214 <= T52;
    end else if(io_resetCounts) begin
      counts_214 <= 4'h0;
    end
    if(reset) begin
      counts_215 <= 4'h0;
    end else if(T1343) begin
      counts_215 <= T52;
    end else if(io_resetCounts) begin
      counts_215 <= 4'h0;
    end
    if(reset) begin
      counts_216 <= 4'h0;
    end else if(T1353) begin
      counts_216 <= T52;
    end else if(io_resetCounts) begin
      counts_216 <= 4'h0;
    end
    if(reset) begin
      counts_217 <= 4'h0;
    end else if(T1357) begin
      counts_217 <= T52;
    end else if(io_resetCounts) begin
      counts_217 <= 4'h0;
    end
    if(reset) begin
      counts_218 <= 4'h0;
    end else if(T1363) begin
      counts_218 <= T52;
    end else if(io_resetCounts) begin
      counts_218 <= 4'h0;
    end
    if(reset) begin
      counts_219 <= 4'h0;
    end else if(T1367) begin
      counts_219 <= T52;
    end else if(io_resetCounts) begin
      counts_219 <= 4'h0;
    end
    if(reset) begin
      counts_220 <= 4'h0;
    end else if(T1375) begin
      counts_220 <= T52;
    end else if(io_resetCounts) begin
      counts_220 <= 4'h0;
    end
    if(reset) begin
      counts_221 <= 4'h0;
    end else if(T1379) begin
      counts_221 <= T52;
    end else if(io_resetCounts) begin
      counts_221 <= 4'h0;
    end
    if(reset) begin
      counts_222 <= 4'h0;
    end else if(T1385) begin
      counts_222 <= T52;
    end else if(io_resetCounts) begin
      counts_222 <= 4'h0;
    end
    if(reset) begin
      counts_223 <= 4'h0;
    end else if(T1389) begin
      counts_223 <= T52;
    end else if(io_resetCounts) begin
      counts_223 <= 4'h0;
    end
    if(reset) begin
      counts_224 <= 4'h0;
    end else if(T1403) begin
      counts_224 <= T52;
    end else if(io_resetCounts) begin
      counts_224 <= 4'h0;
    end
    if(reset) begin
      counts_225 <= 4'h0;
    end else if(T1407) begin
      counts_225 <= T52;
    end else if(io_resetCounts) begin
      counts_225 <= 4'h0;
    end
    if(reset) begin
      counts_226 <= 4'h0;
    end else if(T1413) begin
      counts_226 <= T52;
    end else if(io_resetCounts) begin
      counts_226 <= 4'h0;
    end
    if(reset) begin
      counts_227 <= 4'h0;
    end else if(T1417) begin
      counts_227 <= T52;
    end else if(io_resetCounts) begin
      counts_227 <= 4'h0;
    end
    if(reset) begin
      counts_228 <= 4'h0;
    end else if(T1425) begin
      counts_228 <= T52;
    end else if(io_resetCounts) begin
      counts_228 <= 4'h0;
    end
    if(reset) begin
      counts_229 <= 4'h0;
    end else if(T1429) begin
      counts_229 <= T52;
    end else if(io_resetCounts) begin
      counts_229 <= 4'h0;
    end
    if(reset) begin
      counts_230 <= 4'h0;
    end else if(T1435) begin
      counts_230 <= T52;
    end else if(io_resetCounts) begin
      counts_230 <= 4'h0;
    end
    if(reset) begin
      counts_231 <= 4'h0;
    end else if(T1439) begin
      counts_231 <= T52;
    end else if(io_resetCounts) begin
      counts_231 <= 4'h0;
    end
    if(reset) begin
      counts_232 <= 4'h0;
    end else if(T1449) begin
      counts_232 <= T52;
    end else if(io_resetCounts) begin
      counts_232 <= 4'h0;
    end
    if(reset) begin
      counts_233 <= 4'h0;
    end else if(T1453) begin
      counts_233 <= T52;
    end else if(io_resetCounts) begin
      counts_233 <= 4'h0;
    end
    if(reset) begin
      counts_234 <= 4'h0;
    end else if(T1459) begin
      counts_234 <= T52;
    end else if(io_resetCounts) begin
      counts_234 <= 4'h0;
    end
    if(reset) begin
      counts_235 <= 4'h0;
    end else if(T1463) begin
      counts_235 <= T52;
    end else if(io_resetCounts) begin
      counts_235 <= 4'h0;
    end
    if(reset) begin
      counts_236 <= 4'h0;
    end else if(T1471) begin
      counts_236 <= T52;
    end else if(io_resetCounts) begin
      counts_236 <= 4'h0;
    end
    if(reset) begin
      counts_237 <= 4'h0;
    end else if(T1475) begin
      counts_237 <= T52;
    end else if(io_resetCounts) begin
      counts_237 <= 4'h0;
    end
    if(reset) begin
      counts_238 <= 4'h0;
    end else if(T1481) begin
      counts_238 <= T52;
    end else if(io_resetCounts) begin
      counts_238 <= 4'h0;
    end
    if(reset) begin
      counts_239 <= 4'h0;
    end else if(T1485) begin
      counts_239 <= T52;
    end else if(io_resetCounts) begin
      counts_239 <= 4'h0;
    end
    if(reset) begin
      counts_240 <= 4'h0;
    end else if(T1497) begin
      counts_240 <= T52;
    end else if(io_resetCounts) begin
      counts_240 <= 4'h0;
    end
    if(reset) begin
      counts_241 <= 4'h0;
    end else if(T1501) begin
      counts_241 <= T52;
    end else if(io_resetCounts) begin
      counts_241 <= 4'h0;
    end
    if(reset) begin
      counts_242 <= 4'h0;
    end else if(T1507) begin
      counts_242 <= T52;
    end else if(io_resetCounts) begin
      counts_242 <= 4'h0;
    end
    if(reset) begin
      counts_243 <= 4'h0;
    end else if(T1511) begin
      counts_243 <= T52;
    end else if(io_resetCounts) begin
      counts_243 <= 4'h0;
    end
    if(reset) begin
      counts_244 <= 4'h0;
    end else if(T1519) begin
      counts_244 <= T52;
    end else if(io_resetCounts) begin
      counts_244 <= 4'h0;
    end
    if(reset) begin
      counts_245 <= 4'h0;
    end else if(T1523) begin
      counts_245 <= T52;
    end else if(io_resetCounts) begin
      counts_245 <= 4'h0;
    end
    if(reset) begin
      counts_246 <= 4'h0;
    end else if(T1529) begin
      counts_246 <= T52;
    end else if(io_resetCounts) begin
      counts_246 <= 4'h0;
    end
    if(reset) begin
      counts_247 <= 4'h0;
    end else if(T1533) begin
      counts_247 <= T52;
    end else if(io_resetCounts) begin
      counts_247 <= 4'h0;
    end
    if(reset) begin
      counts_248 <= 4'h0;
    end else if(T1543) begin
      counts_248 <= T52;
    end else if(io_resetCounts) begin
      counts_248 <= 4'h0;
    end
    if(reset) begin
      counts_249 <= 4'h0;
    end else if(T1547) begin
      counts_249 <= T52;
    end else if(io_resetCounts) begin
      counts_249 <= 4'h0;
    end
    if(reset) begin
      counts_250 <= 4'h0;
    end else if(T1553) begin
      counts_250 <= T52;
    end else if(io_resetCounts) begin
      counts_250 <= 4'h0;
    end
    if(reset) begin
      counts_251 <= 4'h0;
    end else if(T1557) begin
      counts_251 <= T52;
    end else if(io_resetCounts) begin
      counts_251 <= 4'h0;
    end
    if(reset) begin
      counts_252 <= 4'h0;
    end else if(T1565) begin
      counts_252 <= T52;
    end else if(io_resetCounts) begin
      counts_252 <= 4'h0;
    end
    if(reset) begin
      counts_253 <= 4'h0;
    end else if(T1569) begin
      counts_253 <= T52;
    end else if(io_resetCounts) begin
      counts_253 <= 4'h0;
    end
    if(reset) begin
      counts_254 <= 4'h0;
    end else if(T1575) begin
      counts_254 <= T52;
    end else if(io_resetCounts) begin
      counts_254 <= 4'h0;
    end
    if(reset) begin
      counts_255 <= 4'h0;
    end else if(T1579) begin
      counts_255 <= T52;
    end else if(io_resetCounts) begin
      counts_255 <= 4'h0;
    end
    if(reset) begin
      counts_256 <= 4'h0;
    end else if(T1599) begin
      counts_256 <= T52;
    end else if(io_resetCounts) begin
      counts_256 <= 4'h0;
    end
    if(reset) begin
      counts_257 <= 4'h0;
    end else if(T1603) begin
      counts_257 <= T52;
    end else if(io_resetCounts) begin
      counts_257 <= 4'h0;
    end
    if(reset) begin
      counts_258 <= 4'h0;
    end else if(T1609) begin
      counts_258 <= T52;
    end else if(io_resetCounts) begin
      counts_258 <= 4'h0;
    end
    if(reset) begin
      counts_259 <= 4'h0;
    end else if(T1613) begin
      counts_259 <= T52;
    end else if(io_resetCounts) begin
      counts_259 <= 4'h0;
    end
    if(reset) begin
      counts_260 <= 4'h0;
    end else if(T1621) begin
      counts_260 <= T52;
    end else if(io_resetCounts) begin
      counts_260 <= 4'h0;
    end
    if(reset) begin
      counts_261 <= 4'h0;
    end else if(T1625) begin
      counts_261 <= T52;
    end else if(io_resetCounts) begin
      counts_261 <= 4'h0;
    end
    if(reset) begin
      counts_262 <= 4'h0;
    end else if(T1631) begin
      counts_262 <= T52;
    end else if(io_resetCounts) begin
      counts_262 <= 4'h0;
    end
    if(reset) begin
      counts_263 <= 4'h0;
    end else if(T1635) begin
      counts_263 <= T52;
    end else if(io_resetCounts) begin
      counts_263 <= 4'h0;
    end
    if(reset) begin
      counts_264 <= 4'h0;
    end else if(T1645) begin
      counts_264 <= T52;
    end else if(io_resetCounts) begin
      counts_264 <= 4'h0;
    end
    if(reset) begin
      counts_265 <= 4'h0;
    end else if(T1649) begin
      counts_265 <= T52;
    end else if(io_resetCounts) begin
      counts_265 <= 4'h0;
    end
    if(reset) begin
      counts_266 <= 4'h0;
    end else if(T1655) begin
      counts_266 <= T52;
    end else if(io_resetCounts) begin
      counts_266 <= 4'h0;
    end
    if(reset) begin
      counts_267 <= 4'h0;
    end else if(T1659) begin
      counts_267 <= T52;
    end else if(io_resetCounts) begin
      counts_267 <= 4'h0;
    end
    if(reset) begin
      counts_268 <= 4'h0;
    end else if(T1667) begin
      counts_268 <= T52;
    end else if(io_resetCounts) begin
      counts_268 <= 4'h0;
    end
    if(reset) begin
      counts_269 <= 4'h0;
    end else if(T1671) begin
      counts_269 <= T52;
    end else if(io_resetCounts) begin
      counts_269 <= 4'h0;
    end
    if(reset) begin
      counts_270 <= 4'h0;
    end else if(T1677) begin
      counts_270 <= T52;
    end else if(io_resetCounts) begin
      counts_270 <= 4'h0;
    end
    if(reset) begin
      counts_271 <= 4'h0;
    end else if(T1681) begin
      counts_271 <= T52;
    end else if(io_resetCounts) begin
      counts_271 <= 4'h0;
    end
    if(reset) begin
      counts_272 <= 4'h0;
    end else if(T1693) begin
      counts_272 <= T52;
    end else if(io_resetCounts) begin
      counts_272 <= 4'h0;
    end
    if(reset) begin
      counts_273 <= 4'h0;
    end else if(T1697) begin
      counts_273 <= T52;
    end else if(io_resetCounts) begin
      counts_273 <= 4'h0;
    end
    if(reset) begin
      counts_274 <= 4'h0;
    end else if(T1703) begin
      counts_274 <= T52;
    end else if(io_resetCounts) begin
      counts_274 <= 4'h0;
    end
    if(reset) begin
      counts_275 <= 4'h0;
    end else if(T1707) begin
      counts_275 <= T52;
    end else if(io_resetCounts) begin
      counts_275 <= 4'h0;
    end
    if(reset) begin
      counts_276 <= 4'h0;
    end else if(T1715) begin
      counts_276 <= T52;
    end else if(io_resetCounts) begin
      counts_276 <= 4'h0;
    end
    if(reset) begin
      counts_277 <= 4'h0;
    end else if(T1719) begin
      counts_277 <= T52;
    end else if(io_resetCounts) begin
      counts_277 <= 4'h0;
    end
    if(reset) begin
      counts_278 <= 4'h0;
    end else if(T1725) begin
      counts_278 <= T52;
    end else if(io_resetCounts) begin
      counts_278 <= 4'h0;
    end
    if(reset) begin
      counts_279 <= 4'h0;
    end else if(T1729) begin
      counts_279 <= T52;
    end else if(io_resetCounts) begin
      counts_279 <= 4'h0;
    end
    if(reset) begin
      counts_280 <= 4'h0;
    end else if(T1739) begin
      counts_280 <= T52;
    end else if(io_resetCounts) begin
      counts_280 <= 4'h0;
    end
    if(reset) begin
      counts_281 <= 4'h0;
    end else if(T1743) begin
      counts_281 <= T52;
    end else if(io_resetCounts) begin
      counts_281 <= 4'h0;
    end
    if(reset) begin
      counts_282 <= 4'h0;
    end else if(T1749) begin
      counts_282 <= T52;
    end else if(io_resetCounts) begin
      counts_282 <= 4'h0;
    end
    if(reset) begin
      counts_283 <= 4'h0;
    end else if(T1753) begin
      counts_283 <= T52;
    end else if(io_resetCounts) begin
      counts_283 <= 4'h0;
    end
    if(reset) begin
      counts_284 <= 4'h0;
    end else if(T1761) begin
      counts_284 <= T52;
    end else if(io_resetCounts) begin
      counts_284 <= 4'h0;
    end
    if(reset) begin
      counts_285 <= 4'h0;
    end else if(T1765) begin
      counts_285 <= T52;
    end else if(io_resetCounts) begin
      counts_285 <= 4'h0;
    end
    if(reset) begin
      counts_286 <= 4'h0;
    end else if(T1771) begin
      counts_286 <= T52;
    end else if(io_resetCounts) begin
      counts_286 <= 4'h0;
    end
    if(reset) begin
      counts_287 <= 4'h0;
    end else if(T1775) begin
      counts_287 <= T52;
    end else if(io_resetCounts) begin
      counts_287 <= 4'h0;
    end
    if(reset) begin
      counts_288 <= 4'h0;
    end else if(T1789) begin
      counts_288 <= T52;
    end else if(io_resetCounts) begin
      counts_288 <= 4'h0;
    end
    if(reset) begin
      counts_289 <= 4'h0;
    end else if(T1793) begin
      counts_289 <= T52;
    end else if(io_resetCounts) begin
      counts_289 <= 4'h0;
    end
    if(reset) begin
      counts_290 <= 4'h0;
    end else if(T1799) begin
      counts_290 <= T52;
    end else if(io_resetCounts) begin
      counts_290 <= 4'h0;
    end
    if(reset) begin
      counts_291 <= 4'h0;
    end else if(T1803) begin
      counts_291 <= T52;
    end else if(io_resetCounts) begin
      counts_291 <= 4'h0;
    end
    if(reset) begin
      counts_292 <= 4'h0;
    end else if(T1811) begin
      counts_292 <= T52;
    end else if(io_resetCounts) begin
      counts_292 <= 4'h0;
    end
    if(reset) begin
      counts_293 <= 4'h0;
    end else if(T1815) begin
      counts_293 <= T52;
    end else if(io_resetCounts) begin
      counts_293 <= 4'h0;
    end
    if(reset) begin
      counts_294 <= 4'h0;
    end else if(T1821) begin
      counts_294 <= T52;
    end else if(io_resetCounts) begin
      counts_294 <= 4'h0;
    end
    if(reset) begin
      counts_295 <= 4'h0;
    end else if(T1825) begin
      counts_295 <= T52;
    end else if(io_resetCounts) begin
      counts_295 <= 4'h0;
    end
    if(reset) begin
      counts_296 <= 4'h0;
    end else if(T1835) begin
      counts_296 <= T52;
    end else if(io_resetCounts) begin
      counts_296 <= 4'h0;
    end
    if(reset) begin
      counts_297 <= 4'h0;
    end else if(T1839) begin
      counts_297 <= T52;
    end else if(io_resetCounts) begin
      counts_297 <= 4'h0;
    end
    if(reset) begin
      counts_298 <= 4'h0;
    end else if(T1845) begin
      counts_298 <= T52;
    end else if(io_resetCounts) begin
      counts_298 <= 4'h0;
    end
    if(reset) begin
      counts_299 <= 4'h0;
    end else if(T1849) begin
      counts_299 <= T52;
    end else if(io_resetCounts) begin
      counts_299 <= 4'h0;
    end
    if(reset) begin
      counts_300 <= 4'h0;
    end else if(T1857) begin
      counts_300 <= T52;
    end else if(io_resetCounts) begin
      counts_300 <= 4'h0;
    end
    if(reset) begin
      counts_301 <= 4'h0;
    end else if(T1861) begin
      counts_301 <= T52;
    end else if(io_resetCounts) begin
      counts_301 <= 4'h0;
    end
    if(reset) begin
      counts_302 <= 4'h0;
    end else if(T1867) begin
      counts_302 <= T52;
    end else if(io_resetCounts) begin
      counts_302 <= 4'h0;
    end
    if(reset) begin
      counts_303 <= 4'h0;
    end else if(T1871) begin
      counts_303 <= T52;
    end else if(io_resetCounts) begin
      counts_303 <= 4'h0;
    end
    if(reset) begin
      counts_304 <= 4'h0;
    end else if(T1883) begin
      counts_304 <= T52;
    end else if(io_resetCounts) begin
      counts_304 <= 4'h0;
    end
    if(reset) begin
      counts_305 <= 4'h0;
    end else if(T1887) begin
      counts_305 <= T52;
    end else if(io_resetCounts) begin
      counts_305 <= 4'h0;
    end
    if(reset) begin
      counts_306 <= 4'h0;
    end else if(T1893) begin
      counts_306 <= T52;
    end else if(io_resetCounts) begin
      counts_306 <= 4'h0;
    end
    if(reset) begin
      counts_307 <= 4'h0;
    end else if(T1897) begin
      counts_307 <= T52;
    end else if(io_resetCounts) begin
      counts_307 <= 4'h0;
    end
    if(reset) begin
      counts_308 <= 4'h0;
    end else if(T1905) begin
      counts_308 <= T52;
    end else if(io_resetCounts) begin
      counts_308 <= 4'h0;
    end
    if(reset) begin
      counts_309 <= 4'h0;
    end else if(T1909) begin
      counts_309 <= T52;
    end else if(io_resetCounts) begin
      counts_309 <= 4'h0;
    end
    if(reset) begin
      counts_310 <= 4'h0;
    end else if(T1915) begin
      counts_310 <= T52;
    end else if(io_resetCounts) begin
      counts_310 <= 4'h0;
    end
    if(reset) begin
      counts_311 <= 4'h0;
    end else if(T1919) begin
      counts_311 <= T52;
    end else if(io_resetCounts) begin
      counts_311 <= 4'h0;
    end
    if(reset) begin
      counts_312 <= 4'h0;
    end else if(T1929) begin
      counts_312 <= T52;
    end else if(io_resetCounts) begin
      counts_312 <= 4'h0;
    end
    if(reset) begin
      counts_313 <= 4'h0;
    end else if(T1933) begin
      counts_313 <= T52;
    end else if(io_resetCounts) begin
      counts_313 <= 4'h0;
    end
    if(reset) begin
      counts_314 <= 4'h0;
    end else if(T1939) begin
      counts_314 <= T52;
    end else if(io_resetCounts) begin
      counts_314 <= 4'h0;
    end
    if(reset) begin
      counts_315 <= 4'h0;
    end else if(T1943) begin
      counts_315 <= T52;
    end else if(io_resetCounts) begin
      counts_315 <= 4'h0;
    end
    if(reset) begin
      counts_316 <= 4'h0;
    end else if(T1951) begin
      counts_316 <= T52;
    end else if(io_resetCounts) begin
      counts_316 <= 4'h0;
    end
    if(reset) begin
      counts_317 <= 4'h0;
    end else if(T1955) begin
      counts_317 <= T52;
    end else if(io_resetCounts) begin
      counts_317 <= 4'h0;
    end
    if(reset) begin
      counts_318 <= 4'h0;
    end else if(T1961) begin
      counts_318 <= T52;
    end else if(io_resetCounts) begin
      counts_318 <= 4'h0;
    end
    if(reset) begin
      counts_319 <= 4'h0;
    end else if(T1965) begin
      counts_319 <= T52;
    end else if(io_resetCounts) begin
      counts_319 <= 4'h0;
    end
    if(reset) begin
      counts_320 <= 4'h0;
    end else if(T1981) begin
      counts_320 <= T52;
    end else if(io_resetCounts) begin
      counts_320 <= 4'h0;
    end
    if(reset) begin
      counts_321 <= 4'h0;
    end else if(T1985) begin
      counts_321 <= T52;
    end else if(io_resetCounts) begin
      counts_321 <= 4'h0;
    end
    if(reset) begin
      counts_322 <= 4'h0;
    end else if(T1991) begin
      counts_322 <= T52;
    end else if(io_resetCounts) begin
      counts_322 <= 4'h0;
    end
    if(reset) begin
      counts_323 <= 4'h0;
    end else if(T1995) begin
      counts_323 <= T52;
    end else if(io_resetCounts) begin
      counts_323 <= 4'h0;
    end
    if(reset) begin
      counts_324 <= 4'h0;
    end else if(T2003) begin
      counts_324 <= T52;
    end else if(io_resetCounts) begin
      counts_324 <= 4'h0;
    end
    if(reset) begin
      counts_325 <= 4'h0;
    end else if(T2007) begin
      counts_325 <= T52;
    end else if(io_resetCounts) begin
      counts_325 <= 4'h0;
    end
    if(reset) begin
      counts_326 <= 4'h0;
    end else if(T2013) begin
      counts_326 <= T52;
    end else if(io_resetCounts) begin
      counts_326 <= 4'h0;
    end
    if(reset) begin
      counts_327 <= 4'h0;
    end else if(T2017) begin
      counts_327 <= T52;
    end else if(io_resetCounts) begin
      counts_327 <= 4'h0;
    end
    if(reset) begin
      counts_328 <= 4'h0;
    end else if(T2027) begin
      counts_328 <= T52;
    end else if(io_resetCounts) begin
      counts_328 <= 4'h0;
    end
    if(reset) begin
      counts_329 <= 4'h0;
    end else if(T2031) begin
      counts_329 <= T52;
    end else if(io_resetCounts) begin
      counts_329 <= 4'h0;
    end
    if(reset) begin
      counts_330 <= 4'h0;
    end else if(T2037) begin
      counts_330 <= T52;
    end else if(io_resetCounts) begin
      counts_330 <= 4'h0;
    end
    if(reset) begin
      counts_331 <= 4'h0;
    end else if(T2041) begin
      counts_331 <= T52;
    end else if(io_resetCounts) begin
      counts_331 <= 4'h0;
    end
    if(reset) begin
      counts_332 <= 4'h0;
    end else if(T2049) begin
      counts_332 <= T52;
    end else if(io_resetCounts) begin
      counts_332 <= 4'h0;
    end
    if(reset) begin
      counts_333 <= 4'h0;
    end else if(T2053) begin
      counts_333 <= T52;
    end else if(io_resetCounts) begin
      counts_333 <= 4'h0;
    end
    if(reset) begin
      counts_334 <= 4'h0;
    end else if(T2059) begin
      counts_334 <= T52;
    end else if(io_resetCounts) begin
      counts_334 <= 4'h0;
    end
    if(reset) begin
      counts_335 <= 4'h0;
    end else if(T2063) begin
      counts_335 <= T52;
    end else if(io_resetCounts) begin
      counts_335 <= 4'h0;
    end
    if(reset) begin
      counts_336 <= 4'h0;
    end else if(T2075) begin
      counts_336 <= T52;
    end else if(io_resetCounts) begin
      counts_336 <= 4'h0;
    end
    if(reset) begin
      counts_337 <= 4'h0;
    end else if(T2079) begin
      counts_337 <= T52;
    end else if(io_resetCounts) begin
      counts_337 <= 4'h0;
    end
    if(reset) begin
      counts_338 <= 4'h0;
    end else if(T2085) begin
      counts_338 <= T52;
    end else if(io_resetCounts) begin
      counts_338 <= 4'h0;
    end
    if(reset) begin
      counts_339 <= 4'h0;
    end else if(T2089) begin
      counts_339 <= T52;
    end else if(io_resetCounts) begin
      counts_339 <= 4'h0;
    end
    if(reset) begin
      counts_340 <= 4'h0;
    end else if(T2097) begin
      counts_340 <= T52;
    end else if(io_resetCounts) begin
      counts_340 <= 4'h0;
    end
    if(reset) begin
      counts_341 <= 4'h0;
    end else if(T2101) begin
      counts_341 <= T52;
    end else if(io_resetCounts) begin
      counts_341 <= 4'h0;
    end
    if(reset) begin
      counts_342 <= 4'h0;
    end else if(T2107) begin
      counts_342 <= T52;
    end else if(io_resetCounts) begin
      counts_342 <= 4'h0;
    end
    if(reset) begin
      counts_343 <= 4'h0;
    end else if(T2111) begin
      counts_343 <= T52;
    end else if(io_resetCounts) begin
      counts_343 <= 4'h0;
    end
    if(reset) begin
      counts_344 <= 4'h0;
    end else if(T2121) begin
      counts_344 <= T52;
    end else if(io_resetCounts) begin
      counts_344 <= 4'h0;
    end
    if(reset) begin
      counts_345 <= 4'h0;
    end else if(T2125) begin
      counts_345 <= T52;
    end else if(io_resetCounts) begin
      counts_345 <= 4'h0;
    end
    if(reset) begin
      counts_346 <= 4'h0;
    end else if(T2131) begin
      counts_346 <= T52;
    end else if(io_resetCounts) begin
      counts_346 <= 4'h0;
    end
    if(reset) begin
      counts_347 <= 4'h0;
    end else if(T2135) begin
      counts_347 <= T52;
    end else if(io_resetCounts) begin
      counts_347 <= 4'h0;
    end
    if(reset) begin
      counts_348 <= 4'h0;
    end else if(T2143) begin
      counts_348 <= T52;
    end else if(io_resetCounts) begin
      counts_348 <= 4'h0;
    end
    if(reset) begin
      counts_349 <= 4'h0;
    end else if(T2147) begin
      counts_349 <= T52;
    end else if(io_resetCounts) begin
      counts_349 <= 4'h0;
    end
    if(reset) begin
      counts_350 <= 4'h0;
    end else if(T2153) begin
      counts_350 <= T52;
    end else if(io_resetCounts) begin
      counts_350 <= 4'h0;
    end
    if(reset) begin
      counts_351 <= 4'h0;
    end else if(T2157) begin
      counts_351 <= T52;
    end else if(io_resetCounts) begin
      counts_351 <= 4'h0;
    end
    if(reset) begin
      counts_352 <= 4'h0;
    end else if(T2171) begin
      counts_352 <= T52;
    end else if(io_resetCounts) begin
      counts_352 <= 4'h0;
    end
    if(reset) begin
      counts_353 <= 4'h0;
    end else if(T2175) begin
      counts_353 <= T52;
    end else if(io_resetCounts) begin
      counts_353 <= 4'h0;
    end
    if(reset) begin
      counts_354 <= 4'h0;
    end else if(T2181) begin
      counts_354 <= T52;
    end else if(io_resetCounts) begin
      counts_354 <= 4'h0;
    end
    if(reset) begin
      counts_355 <= 4'h0;
    end else if(T2185) begin
      counts_355 <= T52;
    end else if(io_resetCounts) begin
      counts_355 <= 4'h0;
    end
    if(reset) begin
      counts_356 <= 4'h0;
    end else if(T2193) begin
      counts_356 <= T52;
    end else if(io_resetCounts) begin
      counts_356 <= 4'h0;
    end
    if(reset) begin
      counts_357 <= 4'h0;
    end else if(T2197) begin
      counts_357 <= T52;
    end else if(io_resetCounts) begin
      counts_357 <= 4'h0;
    end
    if(reset) begin
      counts_358 <= 4'h0;
    end else if(T2203) begin
      counts_358 <= T52;
    end else if(io_resetCounts) begin
      counts_358 <= 4'h0;
    end
    if(reset) begin
      counts_359 <= 4'h0;
    end else if(T2207) begin
      counts_359 <= T52;
    end else if(io_resetCounts) begin
      counts_359 <= 4'h0;
    end
    if(reset) begin
      counts_360 <= 4'h0;
    end else if(T2217) begin
      counts_360 <= T52;
    end else if(io_resetCounts) begin
      counts_360 <= 4'h0;
    end
    if(reset) begin
      counts_361 <= 4'h0;
    end else if(T2221) begin
      counts_361 <= T52;
    end else if(io_resetCounts) begin
      counts_361 <= 4'h0;
    end
    if(reset) begin
      counts_362 <= 4'h0;
    end else if(T2227) begin
      counts_362 <= T52;
    end else if(io_resetCounts) begin
      counts_362 <= 4'h0;
    end
    if(reset) begin
      counts_363 <= 4'h0;
    end else if(T2231) begin
      counts_363 <= T52;
    end else if(io_resetCounts) begin
      counts_363 <= 4'h0;
    end
    if(reset) begin
      counts_364 <= 4'h0;
    end else if(T2239) begin
      counts_364 <= T52;
    end else if(io_resetCounts) begin
      counts_364 <= 4'h0;
    end
    if(reset) begin
      counts_365 <= 4'h0;
    end else if(T2243) begin
      counts_365 <= T52;
    end else if(io_resetCounts) begin
      counts_365 <= 4'h0;
    end
    if(reset) begin
      counts_366 <= 4'h0;
    end else if(T2249) begin
      counts_366 <= T52;
    end else if(io_resetCounts) begin
      counts_366 <= 4'h0;
    end
    if(reset) begin
      counts_367 <= 4'h0;
    end else if(T2253) begin
      counts_367 <= T52;
    end else if(io_resetCounts) begin
      counts_367 <= 4'h0;
    end
    if(reset) begin
      counts_368 <= 4'h0;
    end else if(T2265) begin
      counts_368 <= T52;
    end else if(io_resetCounts) begin
      counts_368 <= 4'h0;
    end
    if(reset) begin
      counts_369 <= 4'h0;
    end else if(T2269) begin
      counts_369 <= T52;
    end else if(io_resetCounts) begin
      counts_369 <= 4'h0;
    end
    if(reset) begin
      counts_370 <= 4'h0;
    end else if(T2275) begin
      counts_370 <= T52;
    end else if(io_resetCounts) begin
      counts_370 <= 4'h0;
    end
    if(reset) begin
      counts_371 <= 4'h0;
    end else if(T2279) begin
      counts_371 <= T52;
    end else if(io_resetCounts) begin
      counts_371 <= 4'h0;
    end
    if(reset) begin
      counts_372 <= 4'h0;
    end else if(T2287) begin
      counts_372 <= T52;
    end else if(io_resetCounts) begin
      counts_372 <= 4'h0;
    end
    if(reset) begin
      counts_373 <= 4'h0;
    end else if(T2291) begin
      counts_373 <= T52;
    end else if(io_resetCounts) begin
      counts_373 <= 4'h0;
    end
    if(reset) begin
      counts_374 <= 4'h0;
    end else if(T2297) begin
      counts_374 <= T52;
    end else if(io_resetCounts) begin
      counts_374 <= 4'h0;
    end
    if(reset) begin
      counts_375 <= 4'h0;
    end else if(T2301) begin
      counts_375 <= T52;
    end else if(io_resetCounts) begin
      counts_375 <= 4'h0;
    end
    if(reset) begin
      counts_376 <= 4'h0;
    end else if(T2311) begin
      counts_376 <= T52;
    end else if(io_resetCounts) begin
      counts_376 <= 4'h0;
    end
    if(reset) begin
      counts_377 <= 4'h0;
    end else if(T2315) begin
      counts_377 <= T52;
    end else if(io_resetCounts) begin
      counts_377 <= 4'h0;
    end
    if(reset) begin
      counts_378 <= 4'h0;
    end else if(T2321) begin
      counts_378 <= T52;
    end else if(io_resetCounts) begin
      counts_378 <= 4'h0;
    end
    if(reset) begin
      counts_379 <= 4'h0;
    end else if(T2325) begin
      counts_379 <= T52;
    end else if(io_resetCounts) begin
      counts_379 <= 4'h0;
    end
    if(reset) begin
      counts_380 <= 4'h0;
    end else if(T2333) begin
      counts_380 <= T52;
    end else if(io_resetCounts) begin
      counts_380 <= 4'h0;
    end
    if(reset) begin
      counts_381 <= 4'h0;
    end else if(T2337) begin
      counts_381 <= T52;
    end else if(io_resetCounts) begin
      counts_381 <= 4'h0;
    end
    if(reset) begin
      counts_382 <= 4'h0;
    end else if(T2343) begin
      counts_382 <= T52;
    end else if(io_resetCounts) begin
      counts_382 <= 4'h0;
    end
    if(reset) begin
      counts_383 <= 4'h0;
    end else if(T2347) begin
      counts_383 <= T52;
    end else if(io_resetCounts) begin
      counts_383 <= 4'h0;
    end
    if(reset) begin
      counts_384 <= 4'h0;
    end else if(T2365) begin
      counts_384 <= T52;
    end else if(io_resetCounts) begin
      counts_384 <= 4'h0;
    end
    if(reset) begin
      counts_385 <= 4'h0;
    end else if(T2369) begin
      counts_385 <= T52;
    end else if(io_resetCounts) begin
      counts_385 <= 4'h0;
    end
    if(reset) begin
      counts_386 <= 4'h0;
    end else if(T2375) begin
      counts_386 <= T52;
    end else if(io_resetCounts) begin
      counts_386 <= 4'h0;
    end
    if(reset) begin
      counts_387 <= 4'h0;
    end else if(T2379) begin
      counts_387 <= T52;
    end else if(io_resetCounts) begin
      counts_387 <= 4'h0;
    end
    if(reset) begin
      counts_388 <= 4'h0;
    end else if(T2387) begin
      counts_388 <= T52;
    end else if(io_resetCounts) begin
      counts_388 <= 4'h0;
    end
    if(reset) begin
      counts_389 <= 4'h0;
    end else if(T2391) begin
      counts_389 <= T52;
    end else if(io_resetCounts) begin
      counts_389 <= 4'h0;
    end
    if(reset) begin
      counts_390 <= 4'h0;
    end else if(T2397) begin
      counts_390 <= T52;
    end else if(io_resetCounts) begin
      counts_390 <= 4'h0;
    end
    if(reset) begin
      counts_391 <= 4'h0;
    end else if(T2401) begin
      counts_391 <= T52;
    end else if(io_resetCounts) begin
      counts_391 <= 4'h0;
    end
    if(reset) begin
      counts_392 <= 4'h0;
    end else if(T2411) begin
      counts_392 <= T52;
    end else if(io_resetCounts) begin
      counts_392 <= 4'h0;
    end
    if(reset) begin
      counts_393 <= 4'h0;
    end else if(T2415) begin
      counts_393 <= T52;
    end else if(io_resetCounts) begin
      counts_393 <= 4'h0;
    end
    if(reset) begin
      counts_394 <= 4'h0;
    end else if(T2421) begin
      counts_394 <= T52;
    end else if(io_resetCounts) begin
      counts_394 <= 4'h0;
    end
    if(reset) begin
      counts_395 <= 4'h0;
    end else if(T2425) begin
      counts_395 <= T52;
    end else if(io_resetCounts) begin
      counts_395 <= 4'h0;
    end
    if(reset) begin
      counts_396 <= 4'h0;
    end else if(T2433) begin
      counts_396 <= T52;
    end else if(io_resetCounts) begin
      counts_396 <= 4'h0;
    end
    if(reset) begin
      counts_397 <= 4'h0;
    end else if(T2437) begin
      counts_397 <= T52;
    end else if(io_resetCounts) begin
      counts_397 <= 4'h0;
    end
    if(reset) begin
      counts_398 <= 4'h0;
    end else if(T2443) begin
      counts_398 <= T52;
    end else if(io_resetCounts) begin
      counts_398 <= 4'h0;
    end
    if(reset) begin
      counts_399 <= 4'h0;
    end else if(T2447) begin
      counts_399 <= T52;
    end else if(io_resetCounts) begin
      counts_399 <= 4'h0;
    end
    if(reset) begin
      counts_400 <= 4'h0;
    end else if(T2459) begin
      counts_400 <= T52;
    end else if(io_resetCounts) begin
      counts_400 <= 4'h0;
    end
    if(reset) begin
      counts_401 <= 4'h0;
    end else if(T2463) begin
      counts_401 <= T52;
    end else if(io_resetCounts) begin
      counts_401 <= 4'h0;
    end
    if(reset) begin
      counts_402 <= 4'h0;
    end else if(T2469) begin
      counts_402 <= T52;
    end else if(io_resetCounts) begin
      counts_402 <= 4'h0;
    end
    if(reset) begin
      counts_403 <= 4'h0;
    end else if(T2473) begin
      counts_403 <= T52;
    end else if(io_resetCounts) begin
      counts_403 <= 4'h0;
    end
    if(reset) begin
      counts_404 <= 4'h0;
    end else if(T2481) begin
      counts_404 <= T52;
    end else if(io_resetCounts) begin
      counts_404 <= 4'h0;
    end
    if(reset) begin
      counts_405 <= 4'h0;
    end else if(T2485) begin
      counts_405 <= T52;
    end else if(io_resetCounts) begin
      counts_405 <= 4'h0;
    end
    if(reset) begin
      counts_406 <= 4'h0;
    end else if(T2491) begin
      counts_406 <= T52;
    end else if(io_resetCounts) begin
      counts_406 <= 4'h0;
    end
    if(reset) begin
      counts_407 <= 4'h0;
    end else if(T2495) begin
      counts_407 <= T52;
    end else if(io_resetCounts) begin
      counts_407 <= 4'h0;
    end
    if(reset) begin
      counts_408 <= 4'h0;
    end else if(T2505) begin
      counts_408 <= T52;
    end else if(io_resetCounts) begin
      counts_408 <= 4'h0;
    end
    if(reset) begin
      counts_409 <= 4'h0;
    end else if(T2509) begin
      counts_409 <= T52;
    end else if(io_resetCounts) begin
      counts_409 <= 4'h0;
    end
    if(reset) begin
      counts_410 <= 4'h0;
    end else if(T2515) begin
      counts_410 <= T52;
    end else if(io_resetCounts) begin
      counts_410 <= 4'h0;
    end
    if(reset) begin
      counts_411 <= 4'h0;
    end else if(T2519) begin
      counts_411 <= T52;
    end else if(io_resetCounts) begin
      counts_411 <= 4'h0;
    end
    if(reset) begin
      counts_412 <= 4'h0;
    end else if(T2527) begin
      counts_412 <= T52;
    end else if(io_resetCounts) begin
      counts_412 <= 4'h0;
    end
    if(reset) begin
      counts_413 <= 4'h0;
    end else if(T2531) begin
      counts_413 <= T52;
    end else if(io_resetCounts) begin
      counts_413 <= 4'h0;
    end
    if(reset) begin
      counts_414 <= 4'h0;
    end else if(T2537) begin
      counts_414 <= T52;
    end else if(io_resetCounts) begin
      counts_414 <= 4'h0;
    end
    if(reset) begin
      counts_415 <= 4'h0;
    end else if(T2541) begin
      counts_415 <= T52;
    end else if(io_resetCounts) begin
      counts_415 <= 4'h0;
    end
    if(reset) begin
      counts_416 <= 4'h0;
    end else if(T2555) begin
      counts_416 <= T52;
    end else if(io_resetCounts) begin
      counts_416 <= 4'h0;
    end
    if(reset) begin
      counts_417 <= 4'h0;
    end else if(T2559) begin
      counts_417 <= T52;
    end else if(io_resetCounts) begin
      counts_417 <= 4'h0;
    end
    if(reset) begin
      counts_418 <= 4'h0;
    end else if(T2565) begin
      counts_418 <= T52;
    end else if(io_resetCounts) begin
      counts_418 <= 4'h0;
    end
    if(reset) begin
      counts_419 <= 4'h0;
    end else if(T2569) begin
      counts_419 <= T52;
    end else if(io_resetCounts) begin
      counts_419 <= 4'h0;
    end
    if(reset) begin
      counts_420 <= 4'h0;
    end else if(T2577) begin
      counts_420 <= T52;
    end else if(io_resetCounts) begin
      counts_420 <= 4'h0;
    end
    if(reset) begin
      counts_421 <= 4'h0;
    end else if(T2581) begin
      counts_421 <= T52;
    end else if(io_resetCounts) begin
      counts_421 <= 4'h0;
    end
    if(reset) begin
      counts_422 <= 4'h0;
    end else if(T2587) begin
      counts_422 <= T52;
    end else if(io_resetCounts) begin
      counts_422 <= 4'h0;
    end
    if(reset) begin
      counts_423 <= 4'h0;
    end else if(T2591) begin
      counts_423 <= T52;
    end else if(io_resetCounts) begin
      counts_423 <= 4'h0;
    end
    if(reset) begin
      counts_424 <= 4'h0;
    end else if(T2601) begin
      counts_424 <= T52;
    end else if(io_resetCounts) begin
      counts_424 <= 4'h0;
    end
    if(reset) begin
      counts_425 <= 4'h0;
    end else if(T2605) begin
      counts_425 <= T52;
    end else if(io_resetCounts) begin
      counts_425 <= 4'h0;
    end
    if(reset) begin
      counts_426 <= 4'h0;
    end else if(T2611) begin
      counts_426 <= T52;
    end else if(io_resetCounts) begin
      counts_426 <= 4'h0;
    end
    if(reset) begin
      counts_427 <= 4'h0;
    end else if(T2615) begin
      counts_427 <= T52;
    end else if(io_resetCounts) begin
      counts_427 <= 4'h0;
    end
    if(reset) begin
      counts_428 <= 4'h0;
    end else if(T2623) begin
      counts_428 <= T52;
    end else if(io_resetCounts) begin
      counts_428 <= 4'h0;
    end
    if(reset) begin
      counts_429 <= 4'h0;
    end else if(T2627) begin
      counts_429 <= T52;
    end else if(io_resetCounts) begin
      counts_429 <= 4'h0;
    end
    if(reset) begin
      counts_430 <= 4'h0;
    end else if(T2633) begin
      counts_430 <= T52;
    end else if(io_resetCounts) begin
      counts_430 <= 4'h0;
    end
    if(reset) begin
      counts_431 <= 4'h0;
    end else if(T2637) begin
      counts_431 <= T52;
    end else if(io_resetCounts) begin
      counts_431 <= 4'h0;
    end
    if(reset) begin
      counts_432 <= 4'h0;
    end else if(T2649) begin
      counts_432 <= T52;
    end else if(io_resetCounts) begin
      counts_432 <= 4'h0;
    end
    if(reset) begin
      counts_433 <= 4'h0;
    end else if(T2653) begin
      counts_433 <= T52;
    end else if(io_resetCounts) begin
      counts_433 <= 4'h0;
    end
    if(reset) begin
      counts_434 <= 4'h0;
    end else if(T2659) begin
      counts_434 <= T52;
    end else if(io_resetCounts) begin
      counts_434 <= 4'h0;
    end
    if(reset) begin
      counts_435 <= 4'h0;
    end else if(T2663) begin
      counts_435 <= T52;
    end else if(io_resetCounts) begin
      counts_435 <= 4'h0;
    end
    if(reset) begin
      counts_436 <= 4'h0;
    end else if(T2671) begin
      counts_436 <= T52;
    end else if(io_resetCounts) begin
      counts_436 <= 4'h0;
    end
    if(reset) begin
      counts_437 <= 4'h0;
    end else if(T2675) begin
      counts_437 <= T52;
    end else if(io_resetCounts) begin
      counts_437 <= 4'h0;
    end
    if(reset) begin
      counts_438 <= 4'h0;
    end else if(T2681) begin
      counts_438 <= T52;
    end else if(io_resetCounts) begin
      counts_438 <= 4'h0;
    end
    if(reset) begin
      counts_439 <= 4'h0;
    end else if(T2685) begin
      counts_439 <= T52;
    end else if(io_resetCounts) begin
      counts_439 <= 4'h0;
    end
    if(reset) begin
      counts_440 <= 4'h0;
    end else if(T2695) begin
      counts_440 <= T52;
    end else if(io_resetCounts) begin
      counts_440 <= 4'h0;
    end
    if(reset) begin
      counts_441 <= 4'h0;
    end else if(T2699) begin
      counts_441 <= T52;
    end else if(io_resetCounts) begin
      counts_441 <= 4'h0;
    end
    if(reset) begin
      counts_442 <= 4'h0;
    end else if(T2705) begin
      counts_442 <= T52;
    end else if(io_resetCounts) begin
      counts_442 <= 4'h0;
    end
    if(reset) begin
      counts_443 <= 4'h0;
    end else if(T2709) begin
      counts_443 <= T52;
    end else if(io_resetCounts) begin
      counts_443 <= 4'h0;
    end
    if(reset) begin
      counts_444 <= 4'h0;
    end else if(T2717) begin
      counts_444 <= T52;
    end else if(io_resetCounts) begin
      counts_444 <= 4'h0;
    end
    if(reset) begin
      counts_445 <= 4'h0;
    end else if(T2721) begin
      counts_445 <= T52;
    end else if(io_resetCounts) begin
      counts_445 <= 4'h0;
    end
    if(reset) begin
      counts_446 <= 4'h0;
    end else if(T2727) begin
      counts_446 <= T52;
    end else if(io_resetCounts) begin
      counts_446 <= 4'h0;
    end
    if(reset) begin
      counts_447 <= 4'h0;
    end else if(T2731) begin
      counts_447 <= T52;
    end else if(io_resetCounts) begin
      counts_447 <= 4'h0;
    end
    if(reset) begin
      counts_448 <= 4'h0;
    end else if(T2747) begin
      counts_448 <= T52;
    end else if(io_resetCounts) begin
      counts_448 <= 4'h0;
    end
    if(reset) begin
      counts_449 <= 4'h0;
    end else if(T2751) begin
      counts_449 <= T52;
    end else if(io_resetCounts) begin
      counts_449 <= 4'h0;
    end
    if(reset) begin
      counts_450 <= 4'h0;
    end else if(T2757) begin
      counts_450 <= T52;
    end else if(io_resetCounts) begin
      counts_450 <= 4'h0;
    end
    if(reset) begin
      counts_451 <= 4'h0;
    end else if(T2761) begin
      counts_451 <= T52;
    end else if(io_resetCounts) begin
      counts_451 <= 4'h0;
    end
    if(reset) begin
      counts_452 <= 4'h0;
    end else if(T2769) begin
      counts_452 <= T52;
    end else if(io_resetCounts) begin
      counts_452 <= 4'h0;
    end
    if(reset) begin
      counts_453 <= 4'h0;
    end else if(T2773) begin
      counts_453 <= T52;
    end else if(io_resetCounts) begin
      counts_453 <= 4'h0;
    end
    if(reset) begin
      counts_454 <= 4'h0;
    end else if(T2779) begin
      counts_454 <= T52;
    end else if(io_resetCounts) begin
      counts_454 <= 4'h0;
    end
    if(reset) begin
      counts_455 <= 4'h0;
    end else if(T2783) begin
      counts_455 <= T52;
    end else if(io_resetCounts) begin
      counts_455 <= 4'h0;
    end
    if(reset) begin
      counts_456 <= 4'h0;
    end else if(T2793) begin
      counts_456 <= T52;
    end else if(io_resetCounts) begin
      counts_456 <= 4'h0;
    end
    if(reset) begin
      counts_457 <= 4'h0;
    end else if(T2797) begin
      counts_457 <= T52;
    end else if(io_resetCounts) begin
      counts_457 <= 4'h0;
    end
    if(reset) begin
      counts_458 <= 4'h0;
    end else if(T2803) begin
      counts_458 <= T52;
    end else if(io_resetCounts) begin
      counts_458 <= 4'h0;
    end
    if(reset) begin
      counts_459 <= 4'h0;
    end else if(T2807) begin
      counts_459 <= T52;
    end else if(io_resetCounts) begin
      counts_459 <= 4'h0;
    end
    if(reset) begin
      counts_460 <= 4'h0;
    end else if(T2815) begin
      counts_460 <= T52;
    end else if(io_resetCounts) begin
      counts_460 <= 4'h0;
    end
    if(reset) begin
      counts_461 <= 4'h0;
    end else if(T2819) begin
      counts_461 <= T52;
    end else if(io_resetCounts) begin
      counts_461 <= 4'h0;
    end
    if(reset) begin
      counts_462 <= 4'h0;
    end else if(T2825) begin
      counts_462 <= T52;
    end else if(io_resetCounts) begin
      counts_462 <= 4'h0;
    end
    if(reset) begin
      counts_463 <= 4'h0;
    end else if(T2829) begin
      counts_463 <= T52;
    end else if(io_resetCounts) begin
      counts_463 <= 4'h0;
    end
    if(reset) begin
      counts_464 <= 4'h0;
    end else if(T2841) begin
      counts_464 <= T52;
    end else if(io_resetCounts) begin
      counts_464 <= 4'h0;
    end
    if(reset) begin
      counts_465 <= 4'h0;
    end else if(T2845) begin
      counts_465 <= T52;
    end else if(io_resetCounts) begin
      counts_465 <= 4'h0;
    end
    if(reset) begin
      counts_466 <= 4'h0;
    end else if(T2851) begin
      counts_466 <= T52;
    end else if(io_resetCounts) begin
      counts_466 <= 4'h0;
    end
    if(reset) begin
      counts_467 <= 4'h0;
    end else if(T2855) begin
      counts_467 <= T52;
    end else if(io_resetCounts) begin
      counts_467 <= 4'h0;
    end
    if(reset) begin
      counts_468 <= 4'h0;
    end else if(T2863) begin
      counts_468 <= T52;
    end else if(io_resetCounts) begin
      counts_468 <= 4'h0;
    end
    if(reset) begin
      counts_469 <= 4'h0;
    end else if(T2867) begin
      counts_469 <= T52;
    end else if(io_resetCounts) begin
      counts_469 <= 4'h0;
    end
    if(reset) begin
      counts_470 <= 4'h0;
    end else if(T2873) begin
      counts_470 <= T52;
    end else if(io_resetCounts) begin
      counts_470 <= 4'h0;
    end
    if(reset) begin
      counts_471 <= 4'h0;
    end else if(T2877) begin
      counts_471 <= T52;
    end else if(io_resetCounts) begin
      counts_471 <= 4'h0;
    end
    if(reset) begin
      counts_472 <= 4'h0;
    end else if(T2887) begin
      counts_472 <= T52;
    end else if(io_resetCounts) begin
      counts_472 <= 4'h0;
    end
    if(reset) begin
      counts_473 <= 4'h0;
    end else if(T2891) begin
      counts_473 <= T52;
    end else if(io_resetCounts) begin
      counts_473 <= 4'h0;
    end
    if(reset) begin
      counts_474 <= 4'h0;
    end else if(T2897) begin
      counts_474 <= T52;
    end else if(io_resetCounts) begin
      counts_474 <= 4'h0;
    end
    if(reset) begin
      counts_475 <= 4'h0;
    end else if(T2901) begin
      counts_475 <= T52;
    end else if(io_resetCounts) begin
      counts_475 <= 4'h0;
    end
    if(reset) begin
      counts_476 <= 4'h0;
    end else if(T2909) begin
      counts_476 <= T52;
    end else if(io_resetCounts) begin
      counts_476 <= 4'h0;
    end
    if(reset) begin
      counts_477 <= 4'h0;
    end else if(T2913) begin
      counts_477 <= T52;
    end else if(io_resetCounts) begin
      counts_477 <= 4'h0;
    end
    if(reset) begin
      counts_478 <= 4'h0;
    end else if(T2919) begin
      counts_478 <= T52;
    end else if(io_resetCounts) begin
      counts_478 <= 4'h0;
    end
    if(reset) begin
      counts_479 <= 4'h0;
    end else if(T2923) begin
      counts_479 <= T52;
    end else if(io_resetCounts) begin
      counts_479 <= 4'h0;
    end
    if(reset) begin
      counts_480 <= 4'h0;
    end else if(T2937) begin
      counts_480 <= T52;
    end else if(io_resetCounts) begin
      counts_480 <= 4'h0;
    end
    if(reset) begin
      counts_481 <= 4'h0;
    end else if(T2941) begin
      counts_481 <= T52;
    end else if(io_resetCounts) begin
      counts_481 <= 4'h0;
    end
    if(reset) begin
      counts_482 <= 4'h0;
    end else if(T2947) begin
      counts_482 <= T52;
    end else if(io_resetCounts) begin
      counts_482 <= 4'h0;
    end
    if(reset) begin
      counts_483 <= 4'h0;
    end else if(T2951) begin
      counts_483 <= T52;
    end else if(io_resetCounts) begin
      counts_483 <= 4'h0;
    end
    if(reset) begin
      counts_484 <= 4'h0;
    end else if(T2959) begin
      counts_484 <= T52;
    end else if(io_resetCounts) begin
      counts_484 <= 4'h0;
    end
    if(reset) begin
      counts_485 <= 4'h0;
    end else if(T2963) begin
      counts_485 <= T52;
    end else if(io_resetCounts) begin
      counts_485 <= 4'h0;
    end
    if(reset) begin
      counts_486 <= 4'h0;
    end else if(T2969) begin
      counts_486 <= T52;
    end else if(io_resetCounts) begin
      counts_486 <= 4'h0;
    end
    if(reset) begin
      counts_487 <= 4'h0;
    end else if(T2973) begin
      counts_487 <= T52;
    end else if(io_resetCounts) begin
      counts_487 <= 4'h0;
    end
    if(reset) begin
      counts_488 <= 4'h0;
    end else if(T2983) begin
      counts_488 <= T52;
    end else if(io_resetCounts) begin
      counts_488 <= 4'h0;
    end
    if(reset) begin
      counts_489 <= 4'h0;
    end else if(T2987) begin
      counts_489 <= T52;
    end else if(io_resetCounts) begin
      counts_489 <= 4'h0;
    end
    if(reset) begin
      counts_490 <= 4'h0;
    end else if(T2993) begin
      counts_490 <= T52;
    end else if(io_resetCounts) begin
      counts_490 <= 4'h0;
    end
    if(reset) begin
      counts_491 <= 4'h0;
    end else if(T2997) begin
      counts_491 <= T52;
    end else if(io_resetCounts) begin
      counts_491 <= 4'h0;
    end
    if(reset) begin
      counts_492 <= 4'h0;
    end else if(T3005) begin
      counts_492 <= T52;
    end else if(io_resetCounts) begin
      counts_492 <= 4'h0;
    end
    if(reset) begin
      counts_493 <= 4'h0;
    end else if(T3009) begin
      counts_493 <= T52;
    end else if(io_resetCounts) begin
      counts_493 <= 4'h0;
    end
    if(reset) begin
      counts_494 <= 4'h0;
    end else if(T3015) begin
      counts_494 <= T52;
    end else if(io_resetCounts) begin
      counts_494 <= 4'h0;
    end
    if(reset) begin
      counts_495 <= 4'h0;
    end else if(T3019) begin
      counts_495 <= T52;
    end else if(io_resetCounts) begin
      counts_495 <= 4'h0;
    end
    if(reset) begin
      counts_496 <= 4'h0;
    end else if(T3031) begin
      counts_496 <= T52;
    end else if(io_resetCounts) begin
      counts_496 <= 4'h0;
    end
    if(reset) begin
      counts_497 <= 4'h0;
    end else if(T3035) begin
      counts_497 <= T52;
    end else if(io_resetCounts) begin
      counts_497 <= 4'h0;
    end
    if(reset) begin
      counts_498 <= 4'h0;
    end else if(T3041) begin
      counts_498 <= T52;
    end else if(io_resetCounts) begin
      counts_498 <= 4'h0;
    end
    if(reset) begin
      counts_499 <= 4'h0;
    end else if(T3045) begin
      counts_499 <= T52;
    end else if(io_resetCounts) begin
      counts_499 <= 4'h0;
    end
    if(reset) begin
      counts_500 <= 4'h0;
    end else if(T3053) begin
      counts_500 <= T52;
    end else if(io_resetCounts) begin
      counts_500 <= 4'h0;
    end
    if(reset) begin
      counts_501 <= 4'h0;
    end else if(T3057) begin
      counts_501 <= T52;
    end else if(io_resetCounts) begin
      counts_501 <= 4'h0;
    end
    if(reset) begin
      counts_502 <= 4'h0;
    end else if(T3063) begin
      counts_502 <= T52;
    end else if(io_resetCounts) begin
      counts_502 <= 4'h0;
    end
    if(reset) begin
      counts_503 <= 4'h0;
    end else if(T3067) begin
      counts_503 <= T52;
    end else if(io_resetCounts) begin
      counts_503 <= 4'h0;
    end
    if(reset) begin
      counts_504 <= 4'h0;
    end else if(T3077) begin
      counts_504 <= T52;
    end else if(io_resetCounts) begin
      counts_504 <= 4'h0;
    end
    if(reset) begin
      counts_505 <= 4'h0;
    end else if(T3081) begin
      counts_505 <= T52;
    end else if(io_resetCounts) begin
      counts_505 <= 4'h0;
    end
    if(reset) begin
      counts_506 <= 4'h0;
    end else if(T3087) begin
      counts_506 <= T52;
    end else if(io_resetCounts) begin
      counts_506 <= 4'h0;
    end
    if(reset) begin
      counts_507 <= 4'h0;
    end else if(T3091) begin
      counts_507 <= T52;
    end else if(io_resetCounts) begin
      counts_507 <= 4'h0;
    end
    if(reset) begin
      counts_508 <= 4'h0;
    end else if(T3099) begin
      counts_508 <= T52;
    end else if(io_resetCounts) begin
      counts_508 <= 4'h0;
    end
    if(reset) begin
      counts_509 <= 4'h0;
    end else if(T3103) begin
      counts_509 <= T52;
    end else if(io_resetCounts) begin
      counts_509 <= 4'h0;
    end
    if(reset) begin
      counts_510 <= 4'h0;
    end else if(T3109) begin
      counts_510 <= T52;
    end else if(io_resetCounts) begin
      counts_510 <= 4'h0;
    end
    if(reset) begin
      counts_511 <= 4'h0;
    end else if(T3113) begin
      counts_511 <= T52;
    end else if(io_resetCounts) begin
      counts_511 <= 4'h0;
    end
    if(reset) begin
      counts_512 <= 4'h0;
    end else if(T3135) begin
      counts_512 <= T52;
    end else if(io_resetCounts) begin
      counts_512 <= 4'h0;
    end
    if(reset) begin
      counts_513 <= 4'h0;
    end else if(T3139) begin
      counts_513 <= T52;
    end else if(io_resetCounts) begin
      counts_513 <= 4'h0;
    end
    if(reset) begin
      counts_514 <= 4'h0;
    end else if(T3145) begin
      counts_514 <= T52;
    end else if(io_resetCounts) begin
      counts_514 <= 4'h0;
    end
    if(reset) begin
      counts_515 <= 4'h0;
    end else if(T3149) begin
      counts_515 <= T52;
    end else if(io_resetCounts) begin
      counts_515 <= 4'h0;
    end
    if(reset) begin
      counts_516 <= 4'h0;
    end else if(T3157) begin
      counts_516 <= T52;
    end else if(io_resetCounts) begin
      counts_516 <= 4'h0;
    end
    if(reset) begin
      counts_517 <= 4'h0;
    end else if(T3161) begin
      counts_517 <= T52;
    end else if(io_resetCounts) begin
      counts_517 <= 4'h0;
    end
    if(reset) begin
      counts_518 <= 4'h0;
    end else if(T3167) begin
      counts_518 <= T52;
    end else if(io_resetCounts) begin
      counts_518 <= 4'h0;
    end
    if(reset) begin
      counts_519 <= 4'h0;
    end else if(T3171) begin
      counts_519 <= T52;
    end else if(io_resetCounts) begin
      counts_519 <= 4'h0;
    end
    if(reset) begin
      counts_520 <= 4'h0;
    end else if(T3181) begin
      counts_520 <= T52;
    end else if(io_resetCounts) begin
      counts_520 <= 4'h0;
    end
    if(reset) begin
      counts_521 <= 4'h0;
    end else if(T3185) begin
      counts_521 <= T52;
    end else if(io_resetCounts) begin
      counts_521 <= 4'h0;
    end
    if(reset) begin
      counts_522 <= 4'h0;
    end else if(T3191) begin
      counts_522 <= T52;
    end else if(io_resetCounts) begin
      counts_522 <= 4'h0;
    end
    if(reset) begin
      counts_523 <= 4'h0;
    end else if(T3195) begin
      counts_523 <= T52;
    end else if(io_resetCounts) begin
      counts_523 <= 4'h0;
    end
    if(reset) begin
      counts_524 <= 4'h0;
    end else if(T3203) begin
      counts_524 <= T52;
    end else if(io_resetCounts) begin
      counts_524 <= 4'h0;
    end
    if(reset) begin
      counts_525 <= 4'h0;
    end else if(T3207) begin
      counts_525 <= T52;
    end else if(io_resetCounts) begin
      counts_525 <= 4'h0;
    end
    if(reset) begin
      counts_526 <= 4'h0;
    end else if(T3213) begin
      counts_526 <= T52;
    end else if(io_resetCounts) begin
      counts_526 <= 4'h0;
    end
    if(reset) begin
      counts_527 <= 4'h0;
    end else if(T3217) begin
      counts_527 <= T52;
    end else if(io_resetCounts) begin
      counts_527 <= 4'h0;
    end
    if(reset) begin
      counts_528 <= 4'h0;
    end else if(T3229) begin
      counts_528 <= T52;
    end else if(io_resetCounts) begin
      counts_528 <= 4'h0;
    end
    if(reset) begin
      counts_529 <= 4'h0;
    end else if(T3233) begin
      counts_529 <= T52;
    end else if(io_resetCounts) begin
      counts_529 <= 4'h0;
    end
    if(reset) begin
      counts_530 <= 4'h0;
    end else if(T3239) begin
      counts_530 <= T52;
    end else if(io_resetCounts) begin
      counts_530 <= 4'h0;
    end
    if(reset) begin
      counts_531 <= 4'h0;
    end else if(T3243) begin
      counts_531 <= T52;
    end else if(io_resetCounts) begin
      counts_531 <= 4'h0;
    end
    if(reset) begin
      counts_532 <= 4'h0;
    end else if(T3251) begin
      counts_532 <= T52;
    end else if(io_resetCounts) begin
      counts_532 <= 4'h0;
    end
    if(reset) begin
      counts_533 <= 4'h0;
    end else if(T3255) begin
      counts_533 <= T52;
    end else if(io_resetCounts) begin
      counts_533 <= 4'h0;
    end
    if(reset) begin
      counts_534 <= 4'h0;
    end else if(T3261) begin
      counts_534 <= T52;
    end else if(io_resetCounts) begin
      counts_534 <= 4'h0;
    end
    if(reset) begin
      counts_535 <= 4'h0;
    end else if(T3265) begin
      counts_535 <= T52;
    end else if(io_resetCounts) begin
      counts_535 <= 4'h0;
    end
    if(reset) begin
      counts_536 <= 4'h0;
    end else if(T3275) begin
      counts_536 <= T52;
    end else if(io_resetCounts) begin
      counts_536 <= 4'h0;
    end
    if(reset) begin
      counts_537 <= 4'h0;
    end else if(T3279) begin
      counts_537 <= T52;
    end else if(io_resetCounts) begin
      counts_537 <= 4'h0;
    end
    if(reset) begin
      counts_538 <= 4'h0;
    end else if(T3285) begin
      counts_538 <= T52;
    end else if(io_resetCounts) begin
      counts_538 <= 4'h0;
    end
    if(reset) begin
      counts_539 <= 4'h0;
    end else if(T3289) begin
      counts_539 <= T52;
    end else if(io_resetCounts) begin
      counts_539 <= 4'h0;
    end
    if(reset) begin
      counts_540 <= 4'h0;
    end else if(T3297) begin
      counts_540 <= T52;
    end else if(io_resetCounts) begin
      counts_540 <= 4'h0;
    end
    if(reset) begin
      counts_541 <= 4'h0;
    end else if(T3301) begin
      counts_541 <= T52;
    end else if(io_resetCounts) begin
      counts_541 <= 4'h0;
    end
    if(reset) begin
      counts_542 <= 4'h0;
    end else if(T3307) begin
      counts_542 <= T52;
    end else if(io_resetCounts) begin
      counts_542 <= 4'h0;
    end
    if(reset) begin
      counts_543 <= 4'h0;
    end else if(T3311) begin
      counts_543 <= T52;
    end else if(io_resetCounts) begin
      counts_543 <= 4'h0;
    end
    if(reset) begin
      counts_544 <= 4'h0;
    end else if(T3325) begin
      counts_544 <= T52;
    end else if(io_resetCounts) begin
      counts_544 <= 4'h0;
    end
    if(reset) begin
      counts_545 <= 4'h0;
    end else if(T3329) begin
      counts_545 <= T52;
    end else if(io_resetCounts) begin
      counts_545 <= 4'h0;
    end
    if(reset) begin
      counts_546 <= 4'h0;
    end else if(T3335) begin
      counts_546 <= T52;
    end else if(io_resetCounts) begin
      counts_546 <= 4'h0;
    end
    if(reset) begin
      counts_547 <= 4'h0;
    end else if(T3339) begin
      counts_547 <= T52;
    end else if(io_resetCounts) begin
      counts_547 <= 4'h0;
    end
    if(reset) begin
      counts_548 <= 4'h0;
    end else if(T3347) begin
      counts_548 <= T52;
    end else if(io_resetCounts) begin
      counts_548 <= 4'h0;
    end
    if(reset) begin
      counts_549 <= 4'h0;
    end else if(T3351) begin
      counts_549 <= T52;
    end else if(io_resetCounts) begin
      counts_549 <= 4'h0;
    end
    if(reset) begin
      counts_550 <= 4'h0;
    end else if(T3357) begin
      counts_550 <= T52;
    end else if(io_resetCounts) begin
      counts_550 <= 4'h0;
    end
    if(reset) begin
      counts_551 <= 4'h0;
    end else if(T3361) begin
      counts_551 <= T52;
    end else if(io_resetCounts) begin
      counts_551 <= 4'h0;
    end
    if(reset) begin
      counts_552 <= 4'h0;
    end else if(T3371) begin
      counts_552 <= T52;
    end else if(io_resetCounts) begin
      counts_552 <= 4'h0;
    end
    if(reset) begin
      counts_553 <= 4'h0;
    end else if(T3375) begin
      counts_553 <= T52;
    end else if(io_resetCounts) begin
      counts_553 <= 4'h0;
    end
    if(reset) begin
      counts_554 <= 4'h0;
    end else if(T3381) begin
      counts_554 <= T52;
    end else if(io_resetCounts) begin
      counts_554 <= 4'h0;
    end
    if(reset) begin
      counts_555 <= 4'h0;
    end else if(T3385) begin
      counts_555 <= T52;
    end else if(io_resetCounts) begin
      counts_555 <= 4'h0;
    end
    if(reset) begin
      counts_556 <= 4'h0;
    end else if(T3393) begin
      counts_556 <= T52;
    end else if(io_resetCounts) begin
      counts_556 <= 4'h0;
    end
    if(reset) begin
      counts_557 <= 4'h0;
    end else if(T3397) begin
      counts_557 <= T52;
    end else if(io_resetCounts) begin
      counts_557 <= 4'h0;
    end
    if(reset) begin
      counts_558 <= 4'h0;
    end else if(T3403) begin
      counts_558 <= T52;
    end else if(io_resetCounts) begin
      counts_558 <= 4'h0;
    end
    if(reset) begin
      counts_559 <= 4'h0;
    end else if(T3407) begin
      counts_559 <= T52;
    end else if(io_resetCounts) begin
      counts_559 <= 4'h0;
    end
    if(reset) begin
      counts_560 <= 4'h0;
    end else if(T3419) begin
      counts_560 <= T52;
    end else if(io_resetCounts) begin
      counts_560 <= 4'h0;
    end
    if(reset) begin
      counts_561 <= 4'h0;
    end else if(T3423) begin
      counts_561 <= T52;
    end else if(io_resetCounts) begin
      counts_561 <= 4'h0;
    end
    if(reset) begin
      counts_562 <= 4'h0;
    end else if(T3429) begin
      counts_562 <= T52;
    end else if(io_resetCounts) begin
      counts_562 <= 4'h0;
    end
    if(reset) begin
      counts_563 <= 4'h0;
    end else if(T3433) begin
      counts_563 <= T52;
    end else if(io_resetCounts) begin
      counts_563 <= 4'h0;
    end
    if(reset) begin
      counts_564 <= 4'h0;
    end else if(T3441) begin
      counts_564 <= T52;
    end else if(io_resetCounts) begin
      counts_564 <= 4'h0;
    end
    if(reset) begin
      counts_565 <= 4'h0;
    end else if(T3445) begin
      counts_565 <= T52;
    end else if(io_resetCounts) begin
      counts_565 <= 4'h0;
    end
    if(reset) begin
      counts_566 <= 4'h0;
    end else if(T3451) begin
      counts_566 <= T52;
    end else if(io_resetCounts) begin
      counts_566 <= 4'h0;
    end
    if(reset) begin
      counts_567 <= 4'h0;
    end else if(T3455) begin
      counts_567 <= T52;
    end else if(io_resetCounts) begin
      counts_567 <= 4'h0;
    end
    if(reset) begin
      counts_568 <= 4'h0;
    end else if(T3465) begin
      counts_568 <= T52;
    end else if(io_resetCounts) begin
      counts_568 <= 4'h0;
    end
    if(reset) begin
      counts_569 <= 4'h0;
    end else if(T3469) begin
      counts_569 <= T52;
    end else if(io_resetCounts) begin
      counts_569 <= 4'h0;
    end
    if(reset) begin
      counts_570 <= 4'h0;
    end else if(T3475) begin
      counts_570 <= T52;
    end else if(io_resetCounts) begin
      counts_570 <= 4'h0;
    end
    if(reset) begin
      counts_571 <= 4'h0;
    end else if(T3479) begin
      counts_571 <= T52;
    end else if(io_resetCounts) begin
      counts_571 <= 4'h0;
    end
    if(reset) begin
      counts_572 <= 4'h0;
    end else if(T3487) begin
      counts_572 <= T52;
    end else if(io_resetCounts) begin
      counts_572 <= 4'h0;
    end
    if(reset) begin
      counts_573 <= 4'h0;
    end else if(T3491) begin
      counts_573 <= T52;
    end else if(io_resetCounts) begin
      counts_573 <= 4'h0;
    end
    if(reset) begin
      counts_574 <= 4'h0;
    end else if(T3497) begin
      counts_574 <= T52;
    end else if(io_resetCounts) begin
      counts_574 <= 4'h0;
    end
    if(reset) begin
      counts_575 <= 4'h0;
    end else if(T3501) begin
      counts_575 <= T52;
    end else if(io_resetCounts) begin
      counts_575 <= 4'h0;
    end
    if(reset) begin
      counts_576 <= 4'h0;
    end else if(T3517) begin
      counts_576 <= T52;
    end else if(io_resetCounts) begin
      counts_576 <= 4'h0;
    end
    if(reset) begin
      counts_577 <= 4'h0;
    end else if(T3521) begin
      counts_577 <= T52;
    end else if(io_resetCounts) begin
      counts_577 <= 4'h0;
    end
    if(reset) begin
      counts_578 <= 4'h0;
    end else if(T3527) begin
      counts_578 <= T52;
    end else if(io_resetCounts) begin
      counts_578 <= 4'h0;
    end
    if(reset) begin
      counts_579 <= 4'h0;
    end else if(T3531) begin
      counts_579 <= T52;
    end else if(io_resetCounts) begin
      counts_579 <= 4'h0;
    end
    if(reset) begin
      counts_580 <= 4'h0;
    end else if(T3539) begin
      counts_580 <= T52;
    end else if(io_resetCounts) begin
      counts_580 <= 4'h0;
    end
    if(reset) begin
      counts_581 <= 4'h0;
    end else if(T3543) begin
      counts_581 <= T52;
    end else if(io_resetCounts) begin
      counts_581 <= 4'h0;
    end
    if(reset) begin
      counts_582 <= 4'h0;
    end else if(T3549) begin
      counts_582 <= T52;
    end else if(io_resetCounts) begin
      counts_582 <= 4'h0;
    end
    if(reset) begin
      counts_583 <= 4'h0;
    end else if(T3553) begin
      counts_583 <= T52;
    end else if(io_resetCounts) begin
      counts_583 <= 4'h0;
    end
    if(reset) begin
      counts_584 <= 4'h0;
    end else if(T3563) begin
      counts_584 <= T52;
    end else if(io_resetCounts) begin
      counts_584 <= 4'h0;
    end
    if(reset) begin
      counts_585 <= 4'h0;
    end else if(T3567) begin
      counts_585 <= T52;
    end else if(io_resetCounts) begin
      counts_585 <= 4'h0;
    end
    if(reset) begin
      counts_586 <= 4'h0;
    end else if(T3573) begin
      counts_586 <= T52;
    end else if(io_resetCounts) begin
      counts_586 <= 4'h0;
    end
    if(reset) begin
      counts_587 <= 4'h0;
    end else if(T3577) begin
      counts_587 <= T52;
    end else if(io_resetCounts) begin
      counts_587 <= 4'h0;
    end
    if(reset) begin
      counts_588 <= 4'h0;
    end else if(T3585) begin
      counts_588 <= T52;
    end else if(io_resetCounts) begin
      counts_588 <= 4'h0;
    end
    if(reset) begin
      counts_589 <= 4'h0;
    end else if(T3589) begin
      counts_589 <= T52;
    end else if(io_resetCounts) begin
      counts_589 <= 4'h0;
    end
    if(reset) begin
      counts_590 <= 4'h0;
    end else if(T3595) begin
      counts_590 <= T52;
    end else if(io_resetCounts) begin
      counts_590 <= 4'h0;
    end
    if(reset) begin
      counts_591 <= 4'h0;
    end else if(T3599) begin
      counts_591 <= T52;
    end else if(io_resetCounts) begin
      counts_591 <= 4'h0;
    end
    if(reset) begin
      counts_592 <= 4'h0;
    end else if(T3611) begin
      counts_592 <= T52;
    end else if(io_resetCounts) begin
      counts_592 <= 4'h0;
    end
    if(reset) begin
      counts_593 <= 4'h0;
    end else if(T3615) begin
      counts_593 <= T52;
    end else if(io_resetCounts) begin
      counts_593 <= 4'h0;
    end
    if(reset) begin
      counts_594 <= 4'h0;
    end else if(T3621) begin
      counts_594 <= T52;
    end else if(io_resetCounts) begin
      counts_594 <= 4'h0;
    end
    if(reset) begin
      counts_595 <= 4'h0;
    end else if(T3625) begin
      counts_595 <= T52;
    end else if(io_resetCounts) begin
      counts_595 <= 4'h0;
    end
    if(reset) begin
      counts_596 <= 4'h0;
    end else if(T3633) begin
      counts_596 <= T52;
    end else if(io_resetCounts) begin
      counts_596 <= 4'h0;
    end
    if(reset) begin
      counts_597 <= 4'h0;
    end else if(T3637) begin
      counts_597 <= T52;
    end else if(io_resetCounts) begin
      counts_597 <= 4'h0;
    end
    if(reset) begin
      counts_598 <= 4'h0;
    end else if(T3643) begin
      counts_598 <= T52;
    end else if(io_resetCounts) begin
      counts_598 <= 4'h0;
    end
    if(reset) begin
      counts_599 <= 4'h0;
    end else if(T3647) begin
      counts_599 <= T52;
    end else if(io_resetCounts) begin
      counts_599 <= 4'h0;
    end
    if(reset) begin
      counts_600 <= 4'h0;
    end else if(T3657) begin
      counts_600 <= T52;
    end else if(io_resetCounts) begin
      counts_600 <= 4'h0;
    end
    if(reset) begin
      counts_601 <= 4'h0;
    end else if(T3661) begin
      counts_601 <= T52;
    end else if(io_resetCounts) begin
      counts_601 <= 4'h0;
    end
    if(reset) begin
      counts_602 <= 4'h0;
    end else if(T3667) begin
      counts_602 <= T52;
    end else if(io_resetCounts) begin
      counts_602 <= 4'h0;
    end
    if(reset) begin
      counts_603 <= 4'h0;
    end else if(T3671) begin
      counts_603 <= T52;
    end else if(io_resetCounts) begin
      counts_603 <= 4'h0;
    end
    if(reset) begin
      counts_604 <= 4'h0;
    end else if(T3679) begin
      counts_604 <= T52;
    end else if(io_resetCounts) begin
      counts_604 <= 4'h0;
    end
    if(reset) begin
      counts_605 <= 4'h0;
    end else if(T3683) begin
      counts_605 <= T52;
    end else if(io_resetCounts) begin
      counts_605 <= 4'h0;
    end
    if(reset) begin
      counts_606 <= 4'h0;
    end else if(T3689) begin
      counts_606 <= T52;
    end else if(io_resetCounts) begin
      counts_606 <= 4'h0;
    end
    if(reset) begin
      counts_607 <= 4'h0;
    end else if(T3693) begin
      counts_607 <= T52;
    end else if(io_resetCounts) begin
      counts_607 <= 4'h0;
    end
    if(reset) begin
      counts_608 <= 4'h0;
    end else if(T3707) begin
      counts_608 <= T52;
    end else if(io_resetCounts) begin
      counts_608 <= 4'h0;
    end
    if(reset) begin
      counts_609 <= 4'h0;
    end else if(T3711) begin
      counts_609 <= T52;
    end else if(io_resetCounts) begin
      counts_609 <= 4'h0;
    end
    if(reset) begin
      counts_610 <= 4'h0;
    end else if(T3717) begin
      counts_610 <= T52;
    end else if(io_resetCounts) begin
      counts_610 <= 4'h0;
    end
    if(reset) begin
      counts_611 <= 4'h0;
    end else if(T3721) begin
      counts_611 <= T52;
    end else if(io_resetCounts) begin
      counts_611 <= 4'h0;
    end
    if(reset) begin
      counts_612 <= 4'h0;
    end else if(T3729) begin
      counts_612 <= T52;
    end else if(io_resetCounts) begin
      counts_612 <= 4'h0;
    end
    if(reset) begin
      counts_613 <= 4'h0;
    end else if(T3733) begin
      counts_613 <= T52;
    end else if(io_resetCounts) begin
      counts_613 <= 4'h0;
    end
    if(reset) begin
      counts_614 <= 4'h0;
    end else if(T3739) begin
      counts_614 <= T52;
    end else if(io_resetCounts) begin
      counts_614 <= 4'h0;
    end
    if(reset) begin
      counts_615 <= 4'h0;
    end else if(T3743) begin
      counts_615 <= T52;
    end else if(io_resetCounts) begin
      counts_615 <= 4'h0;
    end
    if(reset) begin
      counts_616 <= 4'h0;
    end else if(T3753) begin
      counts_616 <= T52;
    end else if(io_resetCounts) begin
      counts_616 <= 4'h0;
    end
    if(reset) begin
      counts_617 <= 4'h0;
    end else if(T3757) begin
      counts_617 <= T52;
    end else if(io_resetCounts) begin
      counts_617 <= 4'h0;
    end
    if(reset) begin
      counts_618 <= 4'h0;
    end else if(T3763) begin
      counts_618 <= T52;
    end else if(io_resetCounts) begin
      counts_618 <= 4'h0;
    end
    if(reset) begin
      counts_619 <= 4'h0;
    end else if(T3767) begin
      counts_619 <= T52;
    end else if(io_resetCounts) begin
      counts_619 <= 4'h0;
    end
    if(reset) begin
      counts_620 <= 4'h0;
    end else if(T3775) begin
      counts_620 <= T52;
    end else if(io_resetCounts) begin
      counts_620 <= 4'h0;
    end
    if(reset) begin
      counts_621 <= 4'h0;
    end else if(T3779) begin
      counts_621 <= T52;
    end else if(io_resetCounts) begin
      counts_621 <= 4'h0;
    end
    if(reset) begin
      counts_622 <= 4'h0;
    end else if(T3785) begin
      counts_622 <= T52;
    end else if(io_resetCounts) begin
      counts_622 <= 4'h0;
    end
    if(reset) begin
      counts_623 <= 4'h0;
    end else if(T3789) begin
      counts_623 <= T52;
    end else if(io_resetCounts) begin
      counts_623 <= 4'h0;
    end
    if(reset) begin
      counts_624 <= 4'h0;
    end else if(T3801) begin
      counts_624 <= T52;
    end else if(io_resetCounts) begin
      counts_624 <= 4'h0;
    end
    if(reset) begin
      counts_625 <= 4'h0;
    end else if(T3805) begin
      counts_625 <= T52;
    end else if(io_resetCounts) begin
      counts_625 <= 4'h0;
    end
    if(reset) begin
      counts_626 <= 4'h0;
    end else if(T3811) begin
      counts_626 <= T52;
    end else if(io_resetCounts) begin
      counts_626 <= 4'h0;
    end
    if(reset) begin
      counts_627 <= 4'h0;
    end else if(T3815) begin
      counts_627 <= T52;
    end else if(io_resetCounts) begin
      counts_627 <= 4'h0;
    end
    if(reset) begin
      counts_628 <= 4'h0;
    end else if(T3823) begin
      counts_628 <= T52;
    end else if(io_resetCounts) begin
      counts_628 <= 4'h0;
    end
    if(reset) begin
      counts_629 <= 4'h0;
    end else if(T3827) begin
      counts_629 <= T52;
    end else if(io_resetCounts) begin
      counts_629 <= 4'h0;
    end
    if(reset) begin
      counts_630 <= 4'h0;
    end else if(T3833) begin
      counts_630 <= T52;
    end else if(io_resetCounts) begin
      counts_630 <= 4'h0;
    end
    if(reset) begin
      counts_631 <= 4'h0;
    end else if(T3837) begin
      counts_631 <= T52;
    end else if(io_resetCounts) begin
      counts_631 <= 4'h0;
    end
    if(reset) begin
      counts_632 <= 4'h0;
    end else if(T3847) begin
      counts_632 <= T52;
    end else if(io_resetCounts) begin
      counts_632 <= 4'h0;
    end
    if(reset) begin
      counts_633 <= 4'h0;
    end else if(T3851) begin
      counts_633 <= T52;
    end else if(io_resetCounts) begin
      counts_633 <= 4'h0;
    end
    if(reset) begin
      counts_634 <= 4'h0;
    end else if(T3857) begin
      counts_634 <= T52;
    end else if(io_resetCounts) begin
      counts_634 <= 4'h0;
    end
    if(reset) begin
      counts_635 <= 4'h0;
    end else if(T3861) begin
      counts_635 <= T52;
    end else if(io_resetCounts) begin
      counts_635 <= 4'h0;
    end
    if(reset) begin
      counts_636 <= 4'h0;
    end else if(T3869) begin
      counts_636 <= T52;
    end else if(io_resetCounts) begin
      counts_636 <= 4'h0;
    end
    if(reset) begin
      counts_637 <= 4'h0;
    end else if(T3873) begin
      counts_637 <= T52;
    end else if(io_resetCounts) begin
      counts_637 <= 4'h0;
    end
    if(reset) begin
      counts_638 <= 4'h0;
    end else if(T3879) begin
      counts_638 <= T52;
    end else if(io_resetCounts) begin
      counts_638 <= 4'h0;
    end
    if(reset) begin
      counts_639 <= 4'h0;
    end else if(T3883) begin
      counts_639 <= T52;
    end else if(io_resetCounts) begin
      counts_639 <= 4'h0;
    end
    if(reset) begin
      counts_640 <= 4'h0;
    end else if(T3901) begin
      counts_640 <= T52;
    end else if(io_resetCounts) begin
      counts_640 <= 4'h0;
    end
    if(reset) begin
      counts_641 <= 4'h0;
    end else if(T3905) begin
      counts_641 <= T52;
    end else if(io_resetCounts) begin
      counts_641 <= 4'h0;
    end
    if(reset) begin
      counts_642 <= 4'h0;
    end else if(T3911) begin
      counts_642 <= T52;
    end else if(io_resetCounts) begin
      counts_642 <= 4'h0;
    end
    if(reset) begin
      counts_643 <= 4'h0;
    end else if(T3915) begin
      counts_643 <= T52;
    end else if(io_resetCounts) begin
      counts_643 <= 4'h0;
    end
    if(reset) begin
      counts_644 <= 4'h0;
    end else if(T3923) begin
      counts_644 <= T52;
    end else if(io_resetCounts) begin
      counts_644 <= 4'h0;
    end
    if(reset) begin
      counts_645 <= 4'h0;
    end else if(T3927) begin
      counts_645 <= T52;
    end else if(io_resetCounts) begin
      counts_645 <= 4'h0;
    end
    if(reset) begin
      counts_646 <= 4'h0;
    end else if(T3933) begin
      counts_646 <= T52;
    end else if(io_resetCounts) begin
      counts_646 <= 4'h0;
    end
    if(reset) begin
      counts_647 <= 4'h0;
    end else if(T3937) begin
      counts_647 <= T52;
    end else if(io_resetCounts) begin
      counts_647 <= 4'h0;
    end
    if(reset) begin
      counts_648 <= 4'h0;
    end else if(T3947) begin
      counts_648 <= T52;
    end else if(io_resetCounts) begin
      counts_648 <= 4'h0;
    end
    if(reset) begin
      counts_649 <= 4'h0;
    end else if(T3951) begin
      counts_649 <= T52;
    end else if(io_resetCounts) begin
      counts_649 <= 4'h0;
    end
    if(reset) begin
      counts_650 <= 4'h0;
    end else if(T3957) begin
      counts_650 <= T52;
    end else if(io_resetCounts) begin
      counts_650 <= 4'h0;
    end
    if(reset) begin
      counts_651 <= 4'h0;
    end else if(T3961) begin
      counts_651 <= T52;
    end else if(io_resetCounts) begin
      counts_651 <= 4'h0;
    end
    if(reset) begin
      counts_652 <= 4'h0;
    end else if(T3969) begin
      counts_652 <= T52;
    end else if(io_resetCounts) begin
      counts_652 <= 4'h0;
    end
    if(reset) begin
      counts_653 <= 4'h0;
    end else if(T3973) begin
      counts_653 <= T52;
    end else if(io_resetCounts) begin
      counts_653 <= 4'h0;
    end
    if(reset) begin
      counts_654 <= 4'h0;
    end else if(T3979) begin
      counts_654 <= T52;
    end else if(io_resetCounts) begin
      counts_654 <= 4'h0;
    end
    if(reset) begin
      counts_655 <= 4'h0;
    end else if(T3983) begin
      counts_655 <= T52;
    end else if(io_resetCounts) begin
      counts_655 <= 4'h0;
    end
    if(reset) begin
      counts_656 <= 4'h0;
    end else if(T3995) begin
      counts_656 <= T52;
    end else if(io_resetCounts) begin
      counts_656 <= 4'h0;
    end
    if(reset) begin
      counts_657 <= 4'h0;
    end else if(T3999) begin
      counts_657 <= T52;
    end else if(io_resetCounts) begin
      counts_657 <= 4'h0;
    end
    if(reset) begin
      counts_658 <= 4'h0;
    end else if(T4005) begin
      counts_658 <= T52;
    end else if(io_resetCounts) begin
      counts_658 <= 4'h0;
    end
    if(reset) begin
      counts_659 <= 4'h0;
    end else if(T4009) begin
      counts_659 <= T52;
    end else if(io_resetCounts) begin
      counts_659 <= 4'h0;
    end
    if(reset) begin
      counts_660 <= 4'h0;
    end else if(T4017) begin
      counts_660 <= T52;
    end else if(io_resetCounts) begin
      counts_660 <= 4'h0;
    end
    if(reset) begin
      counts_661 <= 4'h0;
    end else if(T4021) begin
      counts_661 <= T52;
    end else if(io_resetCounts) begin
      counts_661 <= 4'h0;
    end
    if(reset) begin
      counts_662 <= 4'h0;
    end else if(T4027) begin
      counts_662 <= T52;
    end else if(io_resetCounts) begin
      counts_662 <= 4'h0;
    end
    if(reset) begin
      counts_663 <= 4'h0;
    end else if(T4031) begin
      counts_663 <= T52;
    end else if(io_resetCounts) begin
      counts_663 <= 4'h0;
    end
    if(reset) begin
      counts_664 <= 4'h0;
    end else if(T4041) begin
      counts_664 <= T52;
    end else if(io_resetCounts) begin
      counts_664 <= 4'h0;
    end
    if(reset) begin
      counts_665 <= 4'h0;
    end else if(T4045) begin
      counts_665 <= T52;
    end else if(io_resetCounts) begin
      counts_665 <= 4'h0;
    end
    if(reset) begin
      counts_666 <= 4'h0;
    end else if(T4051) begin
      counts_666 <= T52;
    end else if(io_resetCounts) begin
      counts_666 <= 4'h0;
    end
    if(reset) begin
      counts_667 <= 4'h0;
    end else if(T4055) begin
      counts_667 <= T52;
    end else if(io_resetCounts) begin
      counts_667 <= 4'h0;
    end
    if(reset) begin
      counts_668 <= 4'h0;
    end else if(T4063) begin
      counts_668 <= T52;
    end else if(io_resetCounts) begin
      counts_668 <= 4'h0;
    end
    if(reset) begin
      counts_669 <= 4'h0;
    end else if(T4067) begin
      counts_669 <= T52;
    end else if(io_resetCounts) begin
      counts_669 <= 4'h0;
    end
    if(reset) begin
      counts_670 <= 4'h0;
    end else if(T4073) begin
      counts_670 <= T52;
    end else if(io_resetCounts) begin
      counts_670 <= 4'h0;
    end
    if(reset) begin
      counts_671 <= 4'h0;
    end else if(T4077) begin
      counts_671 <= T52;
    end else if(io_resetCounts) begin
      counts_671 <= 4'h0;
    end
    if(reset) begin
      counts_672 <= 4'h0;
    end else if(T4091) begin
      counts_672 <= T52;
    end else if(io_resetCounts) begin
      counts_672 <= 4'h0;
    end
    if(reset) begin
      counts_673 <= 4'h0;
    end else if(T4095) begin
      counts_673 <= T52;
    end else if(io_resetCounts) begin
      counts_673 <= 4'h0;
    end
    if(reset) begin
      counts_674 <= 4'h0;
    end else if(T4101) begin
      counts_674 <= T52;
    end else if(io_resetCounts) begin
      counts_674 <= 4'h0;
    end
    if(reset) begin
      counts_675 <= 4'h0;
    end else if(T4105) begin
      counts_675 <= T52;
    end else if(io_resetCounts) begin
      counts_675 <= 4'h0;
    end
    if(reset) begin
      counts_676 <= 4'h0;
    end else if(T4113) begin
      counts_676 <= T52;
    end else if(io_resetCounts) begin
      counts_676 <= 4'h0;
    end
    if(reset) begin
      counts_677 <= 4'h0;
    end else if(T4117) begin
      counts_677 <= T52;
    end else if(io_resetCounts) begin
      counts_677 <= 4'h0;
    end
    if(reset) begin
      counts_678 <= 4'h0;
    end else if(T4123) begin
      counts_678 <= T52;
    end else if(io_resetCounts) begin
      counts_678 <= 4'h0;
    end
    if(reset) begin
      counts_679 <= 4'h0;
    end else if(T4127) begin
      counts_679 <= T52;
    end else if(io_resetCounts) begin
      counts_679 <= 4'h0;
    end
    if(reset) begin
      counts_680 <= 4'h0;
    end else if(T4137) begin
      counts_680 <= T52;
    end else if(io_resetCounts) begin
      counts_680 <= 4'h0;
    end
    if(reset) begin
      counts_681 <= 4'h0;
    end else if(T4141) begin
      counts_681 <= T52;
    end else if(io_resetCounts) begin
      counts_681 <= 4'h0;
    end
    if(reset) begin
      counts_682 <= 4'h0;
    end else if(T4147) begin
      counts_682 <= T52;
    end else if(io_resetCounts) begin
      counts_682 <= 4'h0;
    end
    if(reset) begin
      counts_683 <= 4'h0;
    end else if(T4151) begin
      counts_683 <= T52;
    end else if(io_resetCounts) begin
      counts_683 <= 4'h0;
    end
    if(reset) begin
      counts_684 <= 4'h0;
    end else if(T4159) begin
      counts_684 <= T52;
    end else if(io_resetCounts) begin
      counts_684 <= 4'h0;
    end
    if(reset) begin
      counts_685 <= 4'h0;
    end else if(T4163) begin
      counts_685 <= T52;
    end else if(io_resetCounts) begin
      counts_685 <= 4'h0;
    end
    if(reset) begin
      counts_686 <= 4'h0;
    end else if(T4169) begin
      counts_686 <= T52;
    end else if(io_resetCounts) begin
      counts_686 <= 4'h0;
    end
    if(reset) begin
      counts_687 <= 4'h0;
    end else if(T4173) begin
      counts_687 <= T52;
    end else if(io_resetCounts) begin
      counts_687 <= 4'h0;
    end
    if(reset) begin
      counts_688 <= 4'h0;
    end else if(T4185) begin
      counts_688 <= T52;
    end else if(io_resetCounts) begin
      counts_688 <= 4'h0;
    end
    if(reset) begin
      counts_689 <= 4'h0;
    end else if(T4189) begin
      counts_689 <= T52;
    end else if(io_resetCounts) begin
      counts_689 <= 4'h0;
    end
    if(reset) begin
      counts_690 <= 4'h0;
    end else if(T4195) begin
      counts_690 <= T52;
    end else if(io_resetCounts) begin
      counts_690 <= 4'h0;
    end
    if(reset) begin
      counts_691 <= 4'h0;
    end else if(T4199) begin
      counts_691 <= T52;
    end else if(io_resetCounts) begin
      counts_691 <= 4'h0;
    end
    if(reset) begin
      counts_692 <= 4'h0;
    end else if(T4207) begin
      counts_692 <= T52;
    end else if(io_resetCounts) begin
      counts_692 <= 4'h0;
    end
    if(reset) begin
      counts_693 <= 4'h0;
    end else if(T4211) begin
      counts_693 <= T52;
    end else if(io_resetCounts) begin
      counts_693 <= 4'h0;
    end
    if(reset) begin
      counts_694 <= 4'h0;
    end else if(T4217) begin
      counts_694 <= T52;
    end else if(io_resetCounts) begin
      counts_694 <= 4'h0;
    end
    if(reset) begin
      counts_695 <= 4'h0;
    end else if(T4221) begin
      counts_695 <= T52;
    end else if(io_resetCounts) begin
      counts_695 <= 4'h0;
    end
    if(reset) begin
      counts_696 <= 4'h0;
    end else if(T4231) begin
      counts_696 <= T52;
    end else if(io_resetCounts) begin
      counts_696 <= 4'h0;
    end
    if(reset) begin
      counts_697 <= 4'h0;
    end else if(T4235) begin
      counts_697 <= T52;
    end else if(io_resetCounts) begin
      counts_697 <= 4'h0;
    end
    if(reset) begin
      counts_698 <= 4'h0;
    end else if(T4241) begin
      counts_698 <= T52;
    end else if(io_resetCounts) begin
      counts_698 <= 4'h0;
    end
    if(reset) begin
      counts_699 <= 4'h0;
    end else if(T4245) begin
      counts_699 <= T52;
    end else if(io_resetCounts) begin
      counts_699 <= 4'h0;
    end
    if(reset) begin
      counts_700 <= 4'h0;
    end else if(T4253) begin
      counts_700 <= T52;
    end else if(io_resetCounts) begin
      counts_700 <= 4'h0;
    end
    if(reset) begin
      counts_701 <= 4'h0;
    end else if(T4257) begin
      counts_701 <= T52;
    end else if(io_resetCounts) begin
      counts_701 <= 4'h0;
    end
    if(reset) begin
      counts_702 <= 4'h0;
    end else if(T4263) begin
      counts_702 <= T52;
    end else if(io_resetCounts) begin
      counts_702 <= 4'h0;
    end
    if(reset) begin
      counts_703 <= 4'h0;
    end else if(T4267) begin
      counts_703 <= T52;
    end else if(io_resetCounts) begin
      counts_703 <= 4'h0;
    end
    if(reset) begin
      counts_704 <= 4'h0;
    end else if(T4283) begin
      counts_704 <= T52;
    end else if(io_resetCounts) begin
      counts_704 <= 4'h0;
    end
    if(reset) begin
      counts_705 <= 4'h0;
    end else if(T4287) begin
      counts_705 <= T52;
    end else if(io_resetCounts) begin
      counts_705 <= 4'h0;
    end
    if(reset) begin
      counts_706 <= 4'h0;
    end else if(T4293) begin
      counts_706 <= T52;
    end else if(io_resetCounts) begin
      counts_706 <= 4'h0;
    end
    if(reset) begin
      counts_707 <= 4'h0;
    end else if(T4297) begin
      counts_707 <= T52;
    end else if(io_resetCounts) begin
      counts_707 <= 4'h0;
    end
    if(reset) begin
      counts_708 <= 4'h0;
    end else if(T4305) begin
      counts_708 <= T52;
    end else if(io_resetCounts) begin
      counts_708 <= 4'h0;
    end
    if(reset) begin
      counts_709 <= 4'h0;
    end else if(T4309) begin
      counts_709 <= T52;
    end else if(io_resetCounts) begin
      counts_709 <= 4'h0;
    end
    if(reset) begin
      counts_710 <= 4'h0;
    end else if(T4315) begin
      counts_710 <= T52;
    end else if(io_resetCounts) begin
      counts_710 <= 4'h0;
    end
    if(reset) begin
      counts_711 <= 4'h0;
    end else if(T4319) begin
      counts_711 <= T52;
    end else if(io_resetCounts) begin
      counts_711 <= 4'h0;
    end
    if(reset) begin
      counts_712 <= 4'h0;
    end else if(T4329) begin
      counts_712 <= T52;
    end else if(io_resetCounts) begin
      counts_712 <= 4'h0;
    end
    if(reset) begin
      counts_713 <= 4'h0;
    end else if(T4333) begin
      counts_713 <= T52;
    end else if(io_resetCounts) begin
      counts_713 <= 4'h0;
    end
    if(reset) begin
      counts_714 <= 4'h0;
    end else if(T4339) begin
      counts_714 <= T52;
    end else if(io_resetCounts) begin
      counts_714 <= 4'h0;
    end
    if(reset) begin
      counts_715 <= 4'h0;
    end else if(T4343) begin
      counts_715 <= T52;
    end else if(io_resetCounts) begin
      counts_715 <= 4'h0;
    end
    if(reset) begin
      counts_716 <= 4'h0;
    end else if(T4351) begin
      counts_716 <= T52;
    end else if(io_resetCounts) begin
      counts_716 <= 4'h0;
    end
    if(reset) begin
      counts_717 <= 4'h0;
    end else if(T4355) begin
      counts_717 <= T52;
    end else if(io_resetCounts) begin
      counts_717 <= 4'h0;
    end
    if(reset) begin
      counts_718 <= 4'h0;
    end else if(T4361) begin
      counts_718 <= T52;
    end else if(io_resetCounts) begin
      counts_718 <= 4'h0;
    end
    if(reset) begin
      counts_719 <= 4'h0;
    end else if(T4365) begin
      counts_719 <= T52;
    end else if(io_resetCounts) begin
      counts_719 <= 4'h0;
    end
    if(reset) begin
      counts_720 <= 4'h0;
    end else if(T4377) begin
      counts_720 <= T52;
    end else if(io_resetCounts) begin
      counts_720 <= 4'h0;
    end
    if(reset) begin
      counts_721 <= 4'h0;
    end else if(T4381) begin
      counts_721 <= T52;
    end else if(io_resetCounts) begin
      counts_721 <= 4'h0;
    end
    if(reset) begin
      counts_722 <= 4'h0;
    end else if(T4387) begin
      counts_722 <= T52;
    end else if(io_resetCounts) begin
      counts_722 <= 4'h0;
    end
    if(reset) begin
      counts_723 <= 4'h0;
    end else if(T4391) begin
      counts_723 <= T52;
    end else if(io_resetCounts) begin
      counts_723 <= 4'h0;
    end
    if(reset) begin
      counts_724 <= 4'h0;
    end else if(T4399) begin
      counts_724 <= T52;
    end else if(io_resetCounts) begin
      counts_724 <= 4'h0;
    end
    if(reset) begin
      counts_725 <= 4'h0;
    end else if(T4403) begin
      counts_725 <= T52;
    end else if(io_resetCounts) begin
      counts_725 <= 4'h0;
    end
    if(reset) begin
      counts_726 <= 4'h0;
    end else if(T4409) begin
      counts_726 <= T52;
    end else if(io_resetCounts) begin
      counts_726 <= 4'h0;
    end
    if(reset) begin
      counts_727 <= 4'h0;
    end else if(T4413) begin
      counts_727 <= T52;
    end else if(io_resetCounts) begin
      counts_727 <= 4'h0;
    end
    if(reset) begin
      counts_728 <= 4'h0;
    end else if(T4423) begin
      counts_728 <= T52;
    end else if(io_resetCounts) begin
      counts_728 <= 4'h0;
    end
    if(reset) begin
      counts_729 <= 4'h0;
    end else if(T4427) begin
      counts_729 <= T52;
    end else if(io_resetCounts) begin
      counts_729 <= 4'h0;
    end
    if(reset) begin
      counts_730 <= 4'h0;
    end else if(T4433) begin
      counts_730 <= T52;
    end else if(io_resetCounts) begin
      counts_730 <= 4'h0;
    end
    if(reset) begin
      counts_731 <= 4'h0;
    end else if(T4437) begin
      counts_731 <= T52;
    end else if(io_resetCounts) begin
      counts_731 <= 4'h0;
    end
    if(reset) begin
      counts_732 <= 4'h0;
    end else if(T4445) begin
      counts_732 <= T52;
    end else if(io_resetCounts) begin
      counts_732 <= 4'h0;
    end
    if(reset) begin
      counts_733 <= 4'h0;
    end else if(T4449) begin
      counts_733 <= T52;
    end else if(io_resetCounts) begin
      counts_733 <= 4'h0;
    end
    if(reset) begin
      counts_734 <= 4'h0;
    end else if(T4455) begin
      counts_734 <= T52;
    end else if(io_resetCounts) begin
      counts_734 <= 4'h0;
    end
    if(reset) begin
      counts_735 <= 4'h0;
    end else if(T4459) begin
      counts_735 <= T52;
    end else if(io_resetCounts) begin
      counts_735 <= 4'h0;
    end
    if(reset) begin
      counts_736 <= 4'h0;
    end else if(T4473) begin
      counts_736 <= T52;
    end else if(io_resetCounts) begin
      counts_736 <= 4'h0;
    end
    if(reset) begin
      counts_737 <= 4'h0;
    end else if(T4477) begin
      counts_737 <= T52;
    end else if(io_resetCounts) begin
      counts_737 <= 4'h0;
    end
    if(reset) begin
      counts_738 <= 4'h0;
    end else if(T4483) begin
      counts_738 <= T52;
    end else if(io_resetCounts) begin
      counts_738 <= 4'h0;
    end
    if(reset) begin
      counts_739 <= 4'h0;
    end else if(T4487) begin
      counts_739 <= T52;
    end else if(io_resetCounts) begin
      counts_739 <= 4'h0;
    end
    if(reset) begin
      counts_740 <= 4'h0;
    end else if(T4495) begin
      counts_740 <= T52;
    end else if(io_resetCounts) begin
      counts_740 <= 4'h0;
    end
    if(reset) begin
      counts_741 <= 4'h0;
    end else if(T4499) begin
      counts_741 <= T52;
    end else if(io_resetCounts) begin
      counts_741 <= 4'h0;
    end
    if(reset) begin
      counts_742 <= 4'h0;
    end else if(T4505) begin
      counts_742 <= T52;
    end else if(io_resetCounts) begin
      counts_742 <= 4'h0;
    end
    if(reset) begin
      counts_743 <= 4'h0;
    end else if(T4509) begin
      counts_743 <= T52;
    end else if(io_resetCounts) begin
      counts_743 <= 4'h0;
    end
    if(reset) begin
      counts_744 <= 4'h0;
    end else if(T4519) begin
      counts_744 <= T52;
    end else if(io_resetCounts) begin
      counts_744 <= 4'h0;
    end
    if(reset) begin
      counts_745 <= 4'h0;
    end else if(T4523) begin
      counts_745 <= T52;
    end else if(io_resetCounts) begin
      counts_745 <= 4'h0;
    end
    if(reset) begin
      counts_746 <= 4'h0;
    end else if(T4529) begin
      counts_746 <= T52;
    end else if(io_resetCounts) begin
      counts_746 <= 4'h0;
    end
    if(reset) begin
      counts_747 <= 4'h0;
    end else if(T4533) begin
      counts_747 <= T52;
    end else if(io_resetCounts) begin
      counts_747 <= 4'h0;
    end
    if(reset) begin
      counts_748 <= 4'h0;
    end else if(T4541) begin
      counts_748 <= T52;
    end else if(io_resetCounts) begin
      counts_748 <= 4'h0;
    end
    if(reset) begin
      counts_749 <= 4'h0;
    end else if(T4545) begin
      counts_749 <= T52;
    end else if(io_resetCounts) begin
      counts_749 <= 4'h0;
    end
    if(reset) begin
      counts_750 <= 4'h0;
    end else if(T4551) begin
      counts_750 <= T52;
    end else if(io_resetCounts) begin
      counts_750 <= 4'h0;
    end
    if(reset) begin
      counts_751 <= 4'h0;
    end else if(T4555) begin
      counts_751 <= T52;
    end else if(io_resetCounts) begin
      counts_751 <= 4'h0;
    end
    if(reset) begin
      counts_752 <= 4'h0;
    end else if(T4567) begin
      counts_752 <= T52;
    end else if(io_resetCounts) begin
      counts_752 <= 4'h0;
    end
    if(reset) begin
      counts_753 <= 4'h0;
    end else if(T4571) begin
      counts_753 <= T52;
    end else if(io_resetCounts) begin
      counts_753 <= 4'h0;
    end
    if(reset) begin
      counts_754 <= 4'h0;
    end else if(T4577) begin
      counts_754 <= T52;
    end else if(io_resetCounts) begin
      counts_754 <= 4'h0;
    end
    if(reset) begin
      counts_755 <= 4'h0;
    end else if(T4581) begin
      counts_755 <= T52;
    end else if(io_resetCounts) begin
      counts_755 <= 4'h0;
    end
    if(reset) begin
      counts_756 <= 4'h0;
    end else if(T4589) begin
      counts_756 <= T52;
    end else if(io_resetCounts) begin
      counts_756 <= 4'h0;
    end
    if(reset) begin
      counts_757 <= 4'h0;
    end else if(T4593) begin
      counts_757 <= T52;
    end else if(io_resetCounts) begin
      counts_757 <= 4'h0;
    end
    if(reset) begin
      counts_758 <= 4'h0;
    end else if(T4599) begin
      counts_758 <= T52;
    end else if(io_resetCounts) begin
      counts_758 <= 4'h0;
    end
    if(reset) begin
      counts_759 <= 4'h0;
    end else if(T4603) begin
      counts_759 <= T52;
    end else if(io_resetCounts) begin
      counts_759 <= 4'h0;
    end
    if(reset) begin
      counts_760 <= 4'h0;
    end else if(T4613) begin
      counts_760 <= T52;
    end else if(io_resetCounts) begin
      counts_760 <= 4'h0;
    end
    if(reset) begin
      counts_761 <= 4'h0;
    end else if(T4617) begin
      counts_761 <= T52;
    end else if(io_resetCounts) begin
      counts_761 <= 4'h0;
    end
    if(reset) begin
      counts_762 <= 4'h0;
    end else if(T4623) begin
      counts_762 <= T52;
    end else if(io_resetCounts) begin
      counts_762 <= 4'h0;
    end
    if(reset) begin
      counts_763 <= 4'h0;
    end else if(T4627) begin
      counts_763 <= T52;
    end else if(io_resetCounts) begin
      counts_763 <= 4'h0;
    end
    if(reset) begin
      counts_764 <= 4'h0;
    end else if(T4635) begin
      counts_764 <= T52;
    end else if(io_resetCounts) begin
      counts_764 <= 4'h0;
    end
    if(reset) begin
      counts_765 <= 4'h0;
    end else if(T4639) begin
      counts_765 <= T52;
    end else if(io_resetCounts) begin
      counts_765 <= 4'h0;
    end
    if(reset) begin
      counts_766 <= 4'h0;
    end else if(T4645) begin
      counts_766 <= T52;
    end else if(io_resetCounts) begin
      counts_766 <= 4'h0;
    end
    if(reset) begin
      counts_767 <= 4'h0;
    end else if(T4649) begin
      counts_767 <= T52;
    end else if(io_resetCounts) begin
      counts_767 <= 4'h0;
    end
    if(reset) begin
      counts_768 <= 4'h0;
    end else if(T4669) begin
      counts_768 <= T52;
    end else if(io_resetCounts) begin
      counts_768 <= 4'h0;
    end
    if(reset) begin
      counts_769 <= 4'h0;
    end else if(T4673) begin
      counts_769 <= T52;
    end else if(io_resetCounts) begin
      counts_769 <= 4'h0;
    end
    if(reset) begin
      counts_770 <= 4'h0;
    end else if(T4679) begin
      counts_770 <= T52;
    end else if(io_resetCounts) begin
      counts_770 <= 4'h0;
    end
    if(reset) begin
      counts_771 <= 4'h0;
    end else if(T4683) begin
      counts_771 <= T52;
    end else if(io_resetCounts) begin
      counts_771 <= 4'h0;
    end
    if(reset) begin
      counts_772 <= 4'h0;
    end else if(T4691) begin
      counts_772 <= T52;
    end else if(io_resetCounts) begin
      counts_772 <= 4'h0;
    end
    if(reset) begin
      counts_773 <= 4'h0;
    end else if(T4695) begin
      counts_773 <= T52;
    end else if(io_resetCounts) begin
      counts_773 <= 4'h0;
    end
    if(reset) begin
      counts_774 <= 4'h0;
    end else if(T4701) begin
      counts_774 <= T52;
    end else if(io_resetCounts) begin
      counts_774 <= 4'h0;
    end
    if(reset) begin
      counts_775 <= 4'h0;
    end else if(T4705) begin
      counts_775 <= T52;
    end else if(io_resetCounts) begin
      counts_775 <= 4'h0;
    end
    if(reset) begin
      counts_776 <= 4'h0;
    end else if(T4715) begin
      counts_776 <= T52;
    end else if(io_resetCounts) begin
      counts_776 <= 4'h0;
    end
    if(reset) begin
      counts_777 <= 4'h0;
    end else if(T4719) begin
      counts_777 <= T52;
    end else if(io_resetCounts) begin
      counts_777 <= 4'h0;
    end
    if(reset) begin
      counts_778 <= 4'h0;
    end else if(T4725) begin
      counts_778 <= T52;
    end else if(io_resetCounts) begin
      counts_778 <= 4'h0;
    end
    if(reset) begin
      counts_779 <= 4'h0;
    end else if(T4729) begin
      counts_779 <= T52;
    end else if(io_resetCounts) begin
      counts_779 <= 4'h0;
    end
    if(reset) begin
      counts_780 <= 4'h0;
    end else if(T4737) begin
      counts_780 <= T52;
    end else if(io_resetCounts) begin
      counts_780 <= 4'h0;
    end
    if(reset) begin
      counts_781 <= 4'h0;
    end else if(T4741) begin
      counts_781 <= T52;
    end else if(io_resetCounts) begin
      counts_781 <= 4'h0;
    end
    if(reset) begin
      counts_782 <= 4'h0;
    end else if(T4747) begin
      counts_782 <= T52;
    end else if(io_resetCounts) begin
      counts_782 <= 4'h0;
    end
    if(reset) begin
      counts_783 <= 4'h0;
    end else if(T4751) begin
      counts_783 <= T52;
    end else if(io_resetCounts) begin
      counts_783 <= 4'h0;
    end
    if(reset) begin
      counts_784 <= 4'h0;
    end else if(T4763) begin
      counts_784 <= T52;
    end else if(io_resetCounts) begin
      counts_784 <= 4'h0;
    end
    if(reset) begin
      counts_785 <= 4'h0;
    end else if(T4767) begin
      counts_785 <= T52;
    end else if(io_resetCounts) begin
      counts_785 <= 4'h0;
    end
    if(reset) begin
      counts_786 <= 4'h0;
    end else if(T4773) begin
      counts_786 <= T52;
    end else if(io_resetCounts) begin
      counts_786 <= 4'h0;
    end
    if(reset) begin
      counts_787 <= 4'h0;
    end else if(T4777) begin
      counts_787 <= T52;
    end else if(io_resetCounts) begin
      counts_787 <= 4'h0;
    end
    if(reset) begin
      counts_788 <= 4'h0;
    end else if(T4785) begin
      counts_788 <= T52;
    end else if(io_resetCounts) begin
      counts_788 <= 4'h0;
    end
    if(reset) begin
      counts_789 <= 4'h0;
    end else if(T4789) begin
      counts_789 <= T52;
    end else if(io_resetCounts) begin
      counts_789 <= 4'h0;
    end
    if(reset) begin
      counts_790 <= 4'h0;
    end else if(T4795) begin
      counts_790 <= T52;
    end else if(io_resetCounts) begin
      counts_790 <= 4'h0;
    end
    if(reset) begin
      counts_791 <= 4'h0;
    end else if(T4799) begin
      counts_791 <= T52;
    end else if(io_resetCounts) begin
      counts_791 <= 4'h0;
    end
    if(reset) begin
      counts_792 <= 4'h0;
    end else if(T4809) begin
      counts_792 <= T52;
    end else if(io_resetCounts) begin
      counts_792 <= 4'h0;
    end
    if(reset) begin
      counts_793 <= 4'h0;
    end else if(T4813) begin
      counts_793 <= T52;
    end else if(io_resetCounts) begin
      counts_793 <= 4'h0;
    end
    if(reset) begin
      counts_794 <= 4'h0;
    end else if(T4819) begin
      counts_794 <= T52;
    end else if(io_resetCounts) begin
      counts_794 <= 4'h0;
    end
    if(reset) begin
      counts_795 <= 4'h0;
    end else if(T4823) begin
      counts_795 <= T52;
    end else if(io_resetCounts) begin
      counts_795 <= 4'h0;
    end
    if(reset) begin
      counts_796 <= 4'h0;
    end else if(T4831) begin
      counts_796 <= T52;
    end else if(io_resetCounts) begin
      counts_796 <= 4'h0;
    end
    if(reset) begin
      counts_797 <= 4'h0;
    end else if(T4835) begin
      counts_797 <= T52;
    end else if(io_resetCounts) begin
      counts_797 <= 4'h0;
    end
    if(reset) begin
      counts_798 <= 4'h0;
    end else if(T4841) begin
      counts_798 <= T52;
    end else if(io_resetCounts) begin
      counts_798 <= 4'h0;
    end
    if(reset) begin
      counts_799 <= 4'h0;
    end else if(T4845) begin
      counts_799 <= T52;
    end else if(io_resetCounts) begin
      counts_799 <= 4'h0;
    end
    if(reset) begin
      counts_800 <= 4'h0;
    end else if(T4859) begin
      counts_800 <= T52;
    end else if(io_resetCounts) begin
      counts_800 <= 4'h0;
    end
    if(reset) begin
      counts_801 <= 4'h0;
    end else if(T4863) begin
      counts_801 <= T52;
    end else if(io_resetCounts) begin
      counts_801 <= 4'h0;
    end
    if(reset) begin
      counts_802 <= 4'h0;
    end else if(T4869) begin
      counts_802 <= T52;
    end else if(io_resetCounts) begin
      counts_802 <= 4'h0;
    end
    if(reset) begin
      counts_803 <= 4'h0;
    end else if(T4873) begin
      counts_803 <= T52;
    end else if(io_resetCounts) begin
      counts_803 <= 4'h0;
    end
    if(reset) begin
      counts_804 <= 4'h0;
    end else if(T4881) begin
      counts_804 <= T52;
    end else if(io_resetCounts) begin
      counts_804 <= 4'h0;
    end
    if(reset) begin
      counts_805 <= 4'h0;
    end else if(T4885) begin
      counts_805 <= T52;
    end else if(io_resetCounts) begin
      counts_805 <= 4'h0;
    end
    if(reset) begin
      counts_806 <= 4'h0;
    end else if(T4891) begin
      counts_806 <= T52;
    end else if(io_resetCounts) begin
      counts_806 <= 4'h0;
    end
    if(reset) begin
      counts_807 <= 4'h0;
    end else if(T4895) begin
      counts_807 <= T52;
    end else if(io_resetCounts) begin
      counts_807 <= 4'h0;
    end
    if(reset) begin
      counts_808 <= 4'h0;
    end else if(T4905) begin
      counts_808 <= T52;
    end else if(io_resetCounts) begin
      counts_808 <= 4'h0;
    end
    if(reset) begin
      counts_809 <= 4'h0;
    end else if(T4909) begin
      counts_809 <= T52;
    end else if(io_resetCounts) begin
      counts_809 <= 4'h0;
    end
    if(reset) begin
      counts_810 <= 4'h0;
    end else if(T4915) begin
      counts_810 <= T52;
    end else if(io_resetCounts) begin
      counts_810 <= 4'h0;
    end
    if(reset) begin
      counts_811 <= 4'h0;
    end else if(T4919) begin
      counts_811 <= T52;
    end else if(io_resetCounts) begin
      counts_811 <= 4'h0;
    end
    if(reset) begin
      counts_812 <= 4'h0;
    end else if(T4927) begin
      counts_812 <= T52;
    end else if(io_resetCounts) begin
      counts_812 <= 4'h0;
    end
    if(reset) begin
      counts_813 <= 4'h0;
    end else if(T4931) begin
      counts_813 <= T52;
    end else if(io_resetCounts) begin
      counts_813 <= 4'h0;
    end
    if(reset) begin
      counts_814 <= 4'h0;
    end else if(T4937) begin
      counts_814 <= T52;
    end else if(io_resetCounts) begin
      counts_814 <= 4'h0;
    end
    if(reset) begin
      counts_815 <= 4'h0;
    end else if(T4941) begin
      counts_815 <= T52;
    end else if(io_resetCounts) begin
      counts_815 <= 4'h0;
    end
    if(reset) begin
      counts_816 <= 4'h0;
    end else if(T4953) begin
      counts_816 <= T52;
    end else if(io_resetCounts) begin
      counts_816 <= 4'h0;
    end
    if(reset) begin
      counts_817 <= 4'h0;
    end else if(T4957) begin
      counts_817 <= T52;
    end else if(io_resetCounts) begin
      counts_817 <= 4'h0;
    end
    if(reset) begin
      counts_818 <= 4'h0;
    end else if(T4963) begin
      counts_818 <= T52;
    end else if(io_resetCounts) begin
      counts_818 <= 4'h0;
    end
    if(reset) begin
      counts_819 <= 4'h0;
    end else if(T4967) begin
      counts_819 <= T52;
    end else if(io_resetCounts) begin
      counts_819 <= 4'h0;
    end
    if(reset) begin
      counts_820 <= 4'h0;
    end else if(T4975) begin
      counts_820 <= T52;
    end else if(io_resetCounts) begin
      counts_820 <= 4'h0;
    end
    if(reset) begin
      counts_821 <= 4'h0;
    end else if(T4979) begin
      counts_821 <= T52;
    end else if(io_resetCounts) begin
      counts_821 <= 4'h0;
    end
    if(reset) begin
      counts_822 <= 4'h0;
    end else if(T4985) begin
      counts_822 <= T52;
    end else if(io_resetCounts) begin
      counts_822 <= 4'h0;
    end
    if(reset) begin
      counts_823 <= 4'h0;
    end else if(T4989) begin
      counts_823 <= T52;
    end else if(io_resetCounts) begin
      counts_823 <= 4'h0;
    end
    if(reset) begin
      counts_824 <= 4'h0;
    end else if(T4999) begin
      counts_824 <= T52;
    end else if(io_resetCounts) begin
      counts_824 <= 4'h0;
    end
    if(reset) begin
      counts_825 <= 4'h0;
    end else if(T5003) begin
      counts_825 <= T52;
    end else if(io_resetCounts) begin
      counts_825 <= 4'h0;
    end
    if(reset) begin
      counts_826 <= 4'h0;
    end else if(T5009) begin
      counts_826 <= T52;
    end else if(io_resetCounts) begin
      counts_826 <= 4'h0;
    end
    if(reset) begin
      counts_827 <= 4'h0;
    end else if(T5013) begin
      counts_827 <= T52;
    end else if(io_resetCounts) begin
      counts_827 <= 4'h0;
    end
    if(reset) begin
      counts_828 <= 4'h0;
    end else if(T5021) begin
      counts_828 <= T52;
    end else if(io_resetCounts) begin
      counts_828 <= 4'h0;
    end
    if(reset) begin
      counts_829 <= 4'h0;
    end else if(T5025) begin
      counts_829 <= T52;
    end else if(io_resetCounts) begin
      counts_829 <= 4'h0;
    end
    if(reset) begin
      counts_830 <= 4'h0;
    end else if(T5031) begin
      counts_830 <= T52;
    end else if(io_resetCounts) begin
      counts_830 <= 4'h0;
    end
    if(reset) begin
      counts_831 <= 4'h0;
    end else if(T5035) begin
      counts_831 <= T52;
    end else if(io_resetCounts) begin
      counts_831 <= 4'h0;
    end
    if(reset) begin
      counts_832 <= 4'h0;
    end else if(T5051) begin
      counts_832 <= T52;
    end else if(io_resetCounts) begin
      counts_832 <= 4'h0;
    end
    if(reset) begin
      counts_833 <= 4'h0;
    end else if(T5055) begin
      counts_833 <= T52;
    end else if(io_resetCounts) begin
      counts_833 <= 4'h0;
    end
    if(reset) begin
      counts_834 <= 4'h0;
    end else if(T5061) begin
      counts_834 <= T52;
    end else if(io_resetCounts) begin
      counts_834 <= 4'h0;
    end
    if(reset) begin
      counts_835 <= 4'h0;
    end else if(T5065) begin
      counts_835 <= T52;
    end else if(io_resetCounts) begin
      counts_835 <= 4'h0;
    end
    if(reset) begin
      counts_836 <= 4'h0;
    end else if(T5073) begin
      counts_836 <= T52;
    end else if(io_resetCounts) begin
      counts_836 <= 4'h0;
    end
    if(reset) begin
      counts_837 <= 4'h0;
    end else if(T5077) begin
      counts_837 <= T52;
    end else if(io_resetCounts) begin
      counts_837 <= 4'h0;
    end
    if(reset) begin
      counts_838 <= 4'h0;
    end else if(T5083) begin
      counts_838 <= T52;
    end else if(io_resetCounts) begin
      counts_838 <= 4'h0;
    end
    if(reset) begin
      counts_839 <= 4'h0;
    end else if(T5087) begin
      counts_839 <= T52;
    end else if(io_resetCounts) begin
      counts_839 <= 4'h0;
    end
    if(reset) begin
      counts_840 <= 4'h0;
    end else if(T5097) begin
      counts_840 <= T52;
    end else if(io_resetCounts) begin
      counts_840 <= 4'h0;
    end
    if(reset) begin
      counts_841 <= 4'h0;
    end else if(T5101) begin
      counts_841 <= T52;
    end else if(io_resetCounts) begin
      counts_841 <= 4'h0;
    end
    if(reset) begin
      counts_842 <= 4'h0;
    end else if(T5107) begin
      counts_842 <= T52;
    end else if(io_resetCounts) begin
      counts_842 <= 4'h0;
    end
    if(reset) begin
      counts_843 <= 4'h0;
    end else if(T5111) begin
      counts_843 <= T52;
    end else if(io_resetCounts) begin
      counts_843 <= 4'h0;
    end
    if(reset) begin
      counts_844 <= 4'h0;
    end else if(T5119) begin
      counts_844 <= T52;
    end else if(io_resetCounts) begin
      counts_844 <= 4'h0;
    end
    if(reset) begin
      counts_845 <= 4'h0;
    end else if(T5123) begin
      counts_845 <= T52;
    end else if(io_resetCounts) begin
      counts_845 <= 4'h0;
    end
    if(reset) begin
      counts_846 <= 4'h0;
    end else if(T5129) begin
      counts_846 <= T52;
    end else if(io_resetCounts) begin
      counts_846 <= 4'h0;
    end
    if(reset) begin
      counts_847 <= 4'h0;
    end else if(T5133) begin
      counts_847 <= T52;
    end else if(io_resetCounts) begin
      counts_847 <= 4'h0;
    end
    if(reset) begin
      counts_848 <= 4'h0;
    end else if(T5145) begin
      counts_848 <= T52;
    end else if(io_resetCounts) begin
      counts_848 <= 4'h0;
    end
    if(reset) begin
      counts_849 <= 4'h0;
    end else if(T5149) begin
      counts_849 <= T52;
    end else if(io_resetCounts) begin
      counts_849 <= 4'h0;
    end
    if(reset) begin
      counts_850 <= 4'h0;
    end else if(T5155) begin
      counts_850 <= T52;
    end else if(io_resetCounts) begin
      counts_850 <= 4'h0;
    end
    if(reset) begin
      counts_851 <= 4'h0;
    end else if(T5159) begin
      counts_851 <= T52;
    end else if(io_resetCounts) begin
      counts_851 <= 4'h0;
    end
    if(reset) begin
      counts_852 <= 4'h0;
    end else if(T5167) begin
      counts_852 <= T52;
    end else if(io_resetCounts) begin
      counts_852 <= 4'h0;
    end
    if(reset) begin
      counts_853 <= 4'h0;
    end else if(T5171) begin
      counts_853 <= T52;
    end else if(io_resetCounts) begin
      counts_853 <= 4'h0;
    end
    if(reset) begin
      counts_854 <= 4'h0;
    end else if(T5177) begin
      counts_854 <= T52;
    end else if(io_resetCounts) begin
      counts_854 <= 4'h0;
    end
    if(reset) begin
      counts_855 <= 4'h0;
    end else if(T5181) begin
      counts_855 <= T52;
    end else if(io_resetCounts) begin
      counts_855 <= 4'h0;
    end
    if(reset) begin
      counts_856 <= 4'h0;
    end else if(T5191) begin
      counts_856 <= T52;
    end else if(io_resetCounts) begin
      counts_856 <= 4'h0;
    end
    if(reset) begin
      counts_857 <= 4'h0;
    end else if(T5195) begin
      counts_857 <= T52;
    end else if(io_resetCounts) begin
      counts_857 <= 4'h0;
    end
    if(reset) begin
      counts_858 <= 4'h0;
    end else if(T5201) begin
      counts_858 <= T52;
    end else if(io_resetCounts) begin
      counts_858 <= 4'h0;
    end
    if(reset) begin
      counts_859 <= 4'h0;
    end else if(T5205) begin
      counts_859 <= T52;
    end else if(io_resetCounts) begin
      counts_859 <= 4'h0;
    end
    if(reset) begin
      counts_860 <= 4'h0;
    end else if(T5213) begin
      counts_860 <= T52;
    end else if(io_resetCounts) begin
      counts_860 <= 4'h0;
    end
    if(reset) begin
      counts_861 <= 4'h0;
    end else if(T5217) begin
      counts_861 <= T52;
    end else if(io_resetCounts) begin
      counts_861 <= 4'h0;
    end
    if(reset) begin
      counts_862 <= 4'h0;
    end else if(T5223) begin
      counts_862 <= T52;
    end else if(io_resetCounts) begin
      counts_862 <= 4'h0;
    end
    if(reset) begin
      counts_863 <= 4'h0;
    end else if(T5227) begin
      counts_863 <= T52;
    end else if(io_resetCounts) begin
      counts_863 <= 4'h0;
    end
    if(reset) begin
      counts_864 <= 4'h0;
    end else if(T5241) begin
      counts_864 <= T52;
    end else if(io_resetCounts) begin
      counts_864 <= 4'h0;
    end
    if(reset) begin
      counts_865 <= 4'h0;
    end else if(T5245) begin
      counts_865 <= T52;
    end else if(io_resetCounts) begin
      counts_865 <= 4'h0;
    end
    if(reset) begin
      counts_866 <= 4'h0;
    end else if(T5251) begin
      counts_866 <= T52;
    end else if(io_resetCounts) begin
      counts_866 <= 4'h0;
    end
    if(reset) begin
      counts_867 <= 4'h0;
    end else if(T5255) begin
      counts_867 <= T52;
    end else if(io_resetCounts) begin
      counts_867 <= 4'h0;
    end
    if(reset) begin
      counts_868 <= 4'h0;
    end else if(T5263) begin
      counts_868 <= T52;
    end else if(io_resetCounts) begin
      counts_868 <= 4'h0;
    end
    if(reset) begin
      counts_869 <= 4'h0;
    end else if(T5267) begin
      counts_869 <= T52;
    end else if(io_resetCounts) begin
      counts_869 <= 4'h0;
    end
    if(reset) begin
      counts_870 <= 4'h0;
    end else if(T5273) begin
      counts_870 <= T52;
    end else if(io_resetCounts) begin
      counts_870 <= 4'h0;
    end
    if(reset) begin
      counts_871 <= 4'h0;
    end else if(T5277) begin
      counts_871 <= T52;
    end else if(io_resetCounts) begin
      counts_871 <= 4'h0;
    end
    if(reset) begin
      counts_872 <= 4'h0;
    end else if(T5287) begin
      counts_872 <= T52;
    end else if(io_resetCounts) begin
      counts_872 <= 4'h0;
    end
    if(reset) begin
      counts_873 <= 4'h0;
    end else if(T5291) begin
      counts_873 <= T52;
    end else if(io_resetCounts) begin
      counts_873 <= 4'h0;
    end
    if(reset) begin
      counts_874 <= 4'h0;
    end else if(T5297) begin
      counts_874 <= T52;
    end else if(io_resetCounts) begin
      counts_874 <= 4'h0;
    end
    if(reset) begin
      counts_875 <= 4'h0;
    end else if(T5301) begin
      counts_875 <= T52;
    end else if(io_resetCounts) begin
      counts_875 <= 4'h0;
    end
    if(reset) begin
      counts_876 <= 4'h0;
    end else if(T5309) begin
      counts_876 <= T52;
    end else if(io_resetCounts) begin
      counts_876 <= 4'h0;
    end
    if(reset) begin
      counts_877 <= 4'h0;
    end else if(T5313) begin
      counts_877 <= T52;
    end else if(io_resetCounts) begin
      counts_877 <= 4'h0;
    end
    if(reset) begin
      counts_878 <= 4'h0;
    end else if(T5319) begin
      counts_878 <= T52;
    end else if(io_resetCounts) begin
      counts_878 <= 4'h0;
    end
    if(reset) begin
      counts_879 <= 4'h0;
    end else if(T5323) begin
      counts_879 <= T52;
    end else if(io_resetCounts) begin
      counts_879 <= 4'h0;
    end
    if(reset) begin
      counts_880 <= 4'h0;
    end else if(T5335) begin
      counts_880 <= T52;
    end else if(io_resetCounts) begin
      counts_880 <= 4'h0;
    end
    if(reset) begin
      counts_881 <= 4'h0;
    end else if(T5339) begin
      counts_881 <= T52;
    end else if(io_resetCounts) begin
      counts_881 <= 4'h0;
    end
    if(reset) begin
      counts_882 <= 4'h0;
    end else if(T5345) begin
      counts_882 <= T52;
    end else if(io_resetCounts) begin
      counts_882 <= 4'h0;
    end
    if(reset) begin
      counts_883 <= 4'h0;
    end else if(T5349) begin
      counts_883 <= T52;
    end else if(io_resetCounts) begin
      counts_883 <= 4'h0;
    end
    if(reset) begin
      counts_884 <= 4'h0;
    end else if(T5357) begin
      counts_884 <= T52;
    end else if(io_resetCounts) begin
      counts_884 <= 4'h0;
    end
    if(reset) begin
      counts_885 <= 4'h0;
    end else if(T5361) begin
      counts_885 <= T52;
    end else if(io_resetCounts) begin
      counts_885 <= 4'h0;
    end
    if(reset) begin
      counts_886 <= 4'h0;
    end else if(T5367) begin
      counts_886 <= T52;
    end else if(io_resetCounts) begin
      counts_886 <= 4'h0;
    end
    if(reset) begin
      counts_887 <= 4'h0;
    end else if(T5371) begin
      counts_887 <= T52;
    end else if(io_resetCounts) begin
      counts_887 <= 4'h0;
    end
    if(reset) begin
      counts_888 <= 4'h0;
    end else if(T5381) begin
      counts_888 <= T52;
    end else if(io_resetCounts) begin
      counts_888 <= 4'h0;
    end
    if(reset) begin
      counts_889 <= 4'h0;
    end else if(T5385) begin
      counts_889 <= T52;
    end else if(io_resetCounts) begin
      counts_889 <= 4'h0;
    end
    if(reset) begin
      counts_890 <= 4'h0;
    end else if(T5391) begin
      counts_890 <= T52;
    end else if(io_resetCounts) begin
      counts_890 <= 4'h0;
    end
    if(reset) begin
      counts_891 <= 4'h0;
    end else if(T5395) begin
      counts_891 <= T52;
    end else if(io_resetCounts) begin
      counts_891 <= 4'h0;
    end
    if(reset) begin
      counts_892 <= 4'h0;
    end else if(T5403) begin
      counts_892 <= T52;
    end else if(io_resetCounts) begin
      counts_892 <= 4'h0;
    end
    if(reset) begin
      counts_893 <= 4'h0;
    end else if(T5407) begin
      counts_893 <= T52;
    end else if(io_resetCounts) begin
      counts_893 <= 4'h0;
    end
    if(reset) begin
      counts_894 <= 4'h0;
    end else if(T5413) begin
      counts_894 <= T52;
    end else if(io_resetCounts) begin
      counts_894 <= 4'h0;
    end
    if(reset) begin
      counts_895 <= 4'h0;
    end else if(T5417) begin
      counts_895 <= T52;
    end else if(io_resetCounts) begin
      counts_895 <= 4'h0;
    end
    if(reset) begin
      counts_896 <= 4'h0;
    end else if(T5435) begin
      counts_896 <= T52;
    end else if(io_resetCounts) begin
      counts_896 <= 4'h0;
    end
    if(reset) begin
      counts_897 <= 4'h0;
    end else if(T5439) begin
      counts_897 <= T52;
    end else if(io_resetCounts) begin
      counts_897 <= 4'h0;
    end
    if(reset) begin
      counts_898 <= 4'h0;
    end else if(T5445) begin
      counts_898 <= T52;
    end else if(io_resetCounts) begin
      counts_898 <= 4'h0;
    end
    if(reset) begin
      counts_899 <= 4'h0;
    end else if(T5449) begin
      counts_899 <= T52;
    end else if(io_resetCounts) begin
      counts_899 <= 4'h0;
    end
    if(reset) begin
      counts_900 <= 4'h0;
    end else if(T5457) begin
      counts_900 <= T52;
    end else if(io_resetCounts) begin
      counts_900 <= 4'h0;
    end
    if(reset) begin
      counts_901 <= 4'h0;
    end else if(T5461) begin
      counts_901 <= T52;
    end else if(io_resetCounts) begin
      counts_901 <= 4'h0;
    end
    if(reset) begin
      counts_902 <= 4'h0;
    end else if(T5467) begin
      counts_902 <= T52;
    end else if(io_resetCounts) begin
      counts_902 <= 4'h0;
    end
    if(reset) begin
      counts_903 <= 4'h0;
    end else if(T5471) begin
      counts_903 <= T52;
    end else if(io_resetCounts) begin
      counts_903 <= 4'h0;
    end
    if(reset) begin
      counts_904 <= 4'h0;
    end else if(T5481) begin
      counts_904 <= T52;
    end else if(io_resetCounts) begin
      counts_904 <= 4'h0;
    end
    if(reset) begin
      counts_905 <= 4'h0;
    end else if(T5485) begin
      counts_905 <= T52;
    end else if(io_resetCounts) begin
      counts_905 <= 4'h0;
    end
    if(reset) begin
      counts_906 <= 4'h0;
    end else if(T5491) begin
      counts_906 <= T52;
    end else if(io_resetCounts) begin
      counts_906 <= 4'h0;
    end
    if(reset) begin
      counts_907 <= 4'h0;
    end else if(T5495) begin
      counts_907 <= T52;
    end else if(io_resetCounts) begin
      counts_907 <= 4'h0;
    end
    if(reset) begin
      counts_908 <= 4'h0;
    end else if(T5503) begin
      counts_908 <= T52;
    end else if(io_resetCounts) begin
      counts_908 <= 4'h0;
    end
    if(reset) begin
      counts_909 <= 4'h0;
    end else if(T5507) begin
      counts_909 <= T52;
    end else if(io_resetCounts) begin
      counts_909 <= 4'h0;
    end
    if(reset) begin
      counts_910 <= 4'h0;
    end else if(T5513) begin
      counts_910 <= T52;
    end else if(io_resetCounts) begin
      counts_910 <= 4'h0;
    end
    if(reset) begin
      counts_911 <= 4'h0;
    end else if(T5517) begin
      counts_911 <= T52;
    end else if(io_resetCounts) begin
      counts_911 <= 4'h0;
    end
    if(reset) begin
      counts_912 <= 4'h0;
    end else if(T5529) begin
      counts_912 <= T52;
    end else if(io_resetCounts) begin
      counts_912 <= 4'h0;
    end
    if(reset) begin
      counts_913 <= 4'h0;
    end else if(T5533) begin
      counts_913 <= T52;
    end else if(io_resetCounts) begin
      counts_913 <= 4'h0;
    end
    if(reset) begin
      counts_914 <= 4'h0;
    end else if(T5539) begin
      counts_914 <= T52;
    end else if(io_resetCounts) begin
      counts_914 <= 4'h0;
    end
    if(reset) begin
      counts_915 <= 4'h0;
    end else if(T5543) begin
      counts_915 <= T52;
    end else if(io_resetCounts) begin
      counts_915 <= 4'h0;
    end
    if(reset) begin
      counts_916 <= 4'h0;
    end else if(T5551) begin
      counts_916 <= T52;
    end else if(io_resetCounts) begin
      counts_916 <= 4'h0;
    end
    if(reset) begin
      counts_917 <= 4'h0;
    end else if(T5555) begin
      counts_917 <= T52;
    end else if(io_resetCounts) begin
      counts_917 <= 4'h0;
    end
    if(reset) begin
      counts_918 <= 4'h0;
    end else if(T5561) begin
      counts_918 <= T52;
    end else if(io_resetCounts) begin
      counts_918 <= 4'h0;
    end
    if(reset) begin
      counts_919 <= 4'h0;
    end else if(T5565) begin
      counts_919 <= T52;
    end else if(io_resetCounts) begin
      counts_919 <= 4'h0;
    end
    if(reset) begin
      counts_920 <= 4'h0;
    end else if(T5575) begin
      counts_920 <= T52;
    end else if(io_resetCounts) begin
      counts_920 <= 4'h0;
    end
    if(reset) begin
      counts_921 <= 4'h0;
    end else if(T5579) begin
      counts_921 <= T52;
    end else if(io_resetCounts) begin
      counts_921 <= 4'h0;
    end
    if(reset) begin
      counts_922 <= 4'h0;
    end else if(T5585) begin
      counts_922 <= T52;
    end else if(io_resetCounts) begin
      counts_922 <= 4'h0;
    end
    if(reset) begin
      counts_923 <= 4'h0;
    end else if(T5589) begin
      counts_923 <= T52;
    end else if(io_resetCounts) begin
      counts_923 <= 4'h0;
    end
    if(reset) begin
      counts_924 <= 4'h0;
    end else if(T5597) begin
      counts_924 <= T52;
    end else if(io_resetCounts) begin
      counts_924 <= 4'h0;
    end
    if(reset) begin
      counts_925 <= 4'h0;
    end else if(T5601) begin
      counts_925 <= T52;
    end else if(io_resetCounts) begin
      counts_925 <= 4'h0;
    end
    if(reset) begin
      counts_926 <= 4'h0;
    end else if(T5607) begin
      counts_926 <= T52;
    end else if(io_resetCounts) begin
      counts_926 <= 4'h0;
    end
    if(reset) begin
      counts_927 <= 4'h0;
    end else if(T5611) begin
      counts_927 <= T52;
    end else if(io_resetCounts) begin
      counts_927 <= 4'h0;
    end
    if(reset) begin
      counts_928 <= 4'h0;
    end else if(T5625) begin
      counts_928 <= T52;
    end else if(io_resetCounts) begin
      counts_928 <= 4'h0;
    end
    if(reset) begin
      counts_929 <= 4'h0;
    end else if(T5629) begin
      counts_929 <= T52;
    end else if(io_resetCounts) begin
      counts_929 <= 4'h0;
    end
    if(reset) begin
      counts_930 <= 4'h0;
    end else if(T5635) begin
      counts_930 <= T52;
    end else if(io_resetCounts) begin
      counts_930 <= 4'h0;
    end
    if(reset) begin
      counts_931 <= 4'h0;
    end else if(T5639) begin
      counts_931 <= T52;
    end else if(io_resetCounts) begin
      counts_931 <= 4'h0;
    end
    if(reset) begin
      counts_932 <= 4'h0;
    end else if(T5647) begin
      counts_932 <= T52;
    end else if(io_resetCounts) begin
      counts_932 <= 4'h0;
    end
    if(reset) begin
      counts_933 <= 4'h0;
    end else if(T5651) begin
      counts_933 <= T52;
    end else if(io_resetCounts) begin
      counts_933 <= 4'h0;
    end
    if(reset) begin
      counts_934 <= 4'h0;
    end else if(T5657) begin
      counts_934 <= T52;
    end else if(io_resetCounts) begin
      counts_934 <= 4'h0;
    end
    if(reset) begin
      counts_935 <= 4'h0;
    end else if(T5661) begin
      counts_935 <= T52;
    end else if(io_resetCounts) begin
      counts_935 <= 4'h0;
    end
    if(reset) begin
      counts_936 <= 4'h0;
    end else if(T5671) begin
      counts_936 <= T52;
    end else if(io_resetCounts) begin
      counts_936 <= 4'h0;
    end
    if(reset) begin
      counts_937 <= 4'h0;
    end else if(T5675) begin
      counts_937 <= T52;
    end else if(io_resetCounts) begin
      counts_937 <= 4'h0;
    end
    if(reset) begin
      counts_938 <= 4'h0;
    end else if(T5681) begin
      counts_938 <= T52;
    end else if(io_resetCounts) begin
      counts_938 <= 4'h0;
    end
    if(reset) begin
      counts_939 <= 4'h0;
    end else if(T5685) begin
      counts_939 <= T52;
    end else if(io_resetCounts) begin
      counts_939 <= 4'h0;
    end
    if(reset) begin
      counts_940 <= 4'h0;
    end else if(T5693) begin
      counts_940 <= T52;
    end else if(io_resetCounts) begin
      counts_940 <= 4'h0;
    end
    if(reset) begin
      counts_941 <= 4'h0;
    end else if(T5697) begin
      counts_941 <= T52;
    end else if(io_resetCounts) begin
      counts_941 <= 4'h0;
    end
    if(reset) begin
      counts_942 <= 4'h0;
    end else if(T5703) begin
      counts_942 <= T52;
    end else if(io_resetCounts) begin
      counts_942 <= 4'h0;
    end
    if(reset) begin
      counts_943 <= 4'h0;
    end else if(T5707) begin
      counts_943 <= T52;
    end else if(io_resetCounts) begin
      counts_943 <= 4'h0;
    end
    if(reset) begin
      counts_944 <= 4'h0;
    end else if(T5719) begin
      counts_944 <= T52;
    end else if(io_resetCounts) begin
      counts_944 <= 4'h0;
    end
    if(reset) begin
      counts_945 <= 4'h0;
    end else if(T5723) begin
      counts_945 <= T52;
    end else if(io_resetCounts) begin
      counts_945 <= 4'h0;
    end
    if(reset) begin
      counts_946 <= 4'h0;
    end else if(T5729) begin
      counts_946 <= T52;
    end else if(io_resetCounts) begin
      counts_946 <= 4'h0;
    end
    if(reset) begin
      counts_947 <= 4'h0;
    end else if(T5733) begin
      counts_947 <= T52;
    end else if(io_resetCounts) begin
      counts_947 <= 4'h0;
    end
    if(reset) begin
      counts_948 <= 4'h0;
    end else if(T5741) begin
      counts_948 <= T52;
    end else if(io_resetCounts) begin
      counts_948 <= 4'h0;
    end
    if(reset) begin
      counts_949 <= 4'h0;
    end else if(T5745) begin
      counts_949 <= T52;
    end else if(io_resetCounts) begin
      counts_949 <= 4'h0;
    end
    if(reset) begin
      counts_950 <= 4'h0;
    end else if(T5751) begin
      counts_950 <= T52;
    end else if(io_resetCounts) begin
      counts_950 <= 4'h0;
    end
    if(reset) begin
      counts_951 <= 4'h0;
    end else if(T5755) begin
      counts_951 <= T52;
    end else if(io_resetCounts) begin
      counts_951 <= 4'h0;
    end
    if(reset) begin
      counts_952 <= 4'h0;
    end else if(T5765) begin
      counts_952 <= T52;
    end else if(io_resetCounts) begin
      counts_952 <= 4'h0;
    end
    if(reset) begin
      counts_953 <= 4'h0;
    end else if(T5769) begin
      counts_953 <= T52;
    end else if(io_resetCounts) begin
      counts_953 <= 4'h0;
    end
    if(reset) begin
      counts_954 <= 4'h0;
    end else if(T5775) begin
      counts_954 <= T52;
    end else if(io_resetCounts) begin
      counts_954 <= 4'h0;
    end
    if(reset) begin
      counts_955 <= 4'h0;
    end else if(T5779) begin
      counts_955 <= T52;
    end else if(io_resetCounts) begin
      counts_955 <= 4'h0;
    end
    if(reset) begin
      counts_956 <= 4'h0;
    end else if(T5787) begin
      counts_956 <= T52;
    end else if(io_resetCounts) begin
      counts_956 <= 4'h0;
    end
    if(reset) begin
      counts_957 <= 4'h0;
    end else if(T5791) begin
      counts_957 <= T52;
    end else if(io_resetCounts) begin
      counts_957 <= 4'h0;
    end
    if(reset) begin
      counts_958 <= 4'h0;
    end else if(T5797) begin
      counts_958 <= T52;
    end else if(io_resetCounts) begin
      counts_958 <= 4'h0;
    end
    if(reset) begin
      counts_959 <= 4'h0;
    end else if(T5801) begin
      counts_959 <= T52;
    end else if(io_resetCounts) begin
      counts_959 <= 4'h0;
    end
    if(reset) begin
      counts_960 <= 4'h0;
    end else if(T5817) begin
      counts_960 <= T52;
    end else if(io_resetCounts) begin
      counts_960 <= 4'h0;
    end
    if(reset) begin
      counts_961 <= 4'h0;
    end else if(T5821) begin
      counts_961 <= T52;
    end else if(io_resetCounts) begin
      counts_961 <= 4'h0;
    end
    if(reset) begin
      counts_962 <= 4'h0;
    end else if(T5827) begin
      counts_962 <= T52;
    end else if(io_resetCounts) begin
      counts_962 <= 4'h0;
    end
    if(reset) begin
      counts_963 <= 4'h0;
    end else if(T5831) begin
      counts_963 <= T52;
    end else if(io_resetCounts) begin
      counts_963 <= 4'h0;
    end
    if(reset) begin
      counts_964 <= 4'h0;
    end else if(T5839) begin
      counts_964 <= T52;
    end else if(io_resetCounts) begin
      counts_964 <= 4'h0;
    end
    if(reset) begin
      counts_965 <= 4'h0;
    end else if(T5843) begin
      counts_965 <= T52;
    end else if(io_resetCounts) begin
      counts_965 <= 4'h0;
    end
    if(reset) begin
      counts_966 <= 4'h0;
    end else if(T5849) begin
      counts_966 <= T52;
    end else if(io_resetCounts) begin
      counts_966 <= 4'h0;
    end
    if(reset) begin
      counts_967 <= 4'h0;
    end else if(T5853) begin
      counts_967 <= T52;
    end else if(io_resetCounts) begin
      counts_967 <= 4'h0;
    end
    if(reset) begin
      counts_968 <= 4'h0;
    end else if(T5863) begin
      counts_968 <= T52;
    end else if(io_resetCounts) begin
      counts_968 <= 4'h0;
    end
    if(reset) begin
      counts_969 <= 4'h0;
    end else if(T5867) begin
      counts_969 <= T52;
    end else if(io_resetCounts) begin
      counts_969 <= 4'h0;
    end
    if(reset) begin
      counts_970 <= 4'h0;
    end else if(T5873) begin
      counts_970 <= T52;
    end else if(io_resetCounts) begin
      counts_970 <= 4'h0;
    end
    if(reset) begin
      counts_971 <= 4'h0;
    end else if(T5877) begin
      counts_971 <= T52;
    end else if(io_resetCounts) begin
      counts_971 <= 4'h0;
    end
    if(reset) begin
      counts_972 <= 4'h0;
    end else if(T5885) begin
      counts_972 <= T52;
    end else if(io_resetCounts) begin
      counts_972 <= 4'h0;
    end
    if(reset) begin
      counts_973 <= 4'h0;
    end else if(T5889) begin
      counts_973 <= T52;
    end else if(io_resetCounts) begin
      counts_973 <= 4'h0;
    end
    if(reset) begin
      counts_974 <= 4'h0;
    end else if(T5895) begin
      counts_974 <= T52;
    end else if(io_resetCounts) begin
      counts_974 <= 4'h0;
    end
    if(reset) begin
      counts_975 <= 4'h0;
    end else if(T5899) begin
      counts_975 <= T52;
    end else if(io_resetCounts) begin
      counts_975 <= 4'h0;
    end
    if(reset) begin
      counts_976 <= 4'h0;
    end else if(T5911) begin
      counts_976 <= T52;
    end else if(io_resetCounts) begin
      counts_976 <= 4'h0;
    end
    if(reset) begin
      counts_977 <= 4'h0;
    end else if(T5915) begin
      counts_977 <= T52;
    end else if(io_resetCounts) begin
      counts_977 <= 4'h0;
    end
    if(reset) begin
      counts_978 <= 4'h0;
    end else if(T5921) begin
      counts_978 <= T52;
    end else if(io_resetCounts) begin
      counts_978 <= 4'h0;
    end
    if(reset) begin
      counts_979 <= 4'h0;
    end else if(T5925) begin
      counts_979 <= T52;
    end else if(io_resetCounts) begin
      counts_979 <= 4'h0;
    end
    if(reset) begin
      counts_980 <= 4'h0;
    end else if(T5933) begin
      counts_980 <= T52;
    end else if(io_resetCounts) begin
      counts_980 <= 4'h0;
    end
    if(reset) begin
      counts_981 <= 4'h0;
    end else if(T5937) begin
      counts_981 <= T52;
    end else if(io_resetCounts) begin
      counts_981 <= 4'h0;
    end
    if(reset) begin
      counts_982 <= 4'h0;
    end else if(T5943) begin
      counts_982 <= T52;
    end else if(io_resetCounts) begin
      counts_982 <= 4'h0;
    end
    if(reset) begin
      counts_983 <= 4'h0;
    end else if(T5947) begin
      counts_983 <= T52;
    end else if(io_resetCounts) begin
      counts_983 <= 4'h0;
    end
    if(reset) begin
      counts_984 <= 4'h0;
    end else if(T5957) begin
      counts_984 <= T52;
    end else if(io_resetCounts) begin
      counts_984 <= 4'h0;
    end
    if(reset) begin
      counts_985 <= 4'h0;
    end else if(T5961) begin
      counts_985 <= T52;
    end else if(io_resetCounts) begin
      counts_985 <= 4'h0;
    end
    if(reset) begin
      counts_986 <= 4'h0;
    end else if(T5967) begin
      counts_986 <= T52;
    end else if(io_resetCounts) begin
      counts_986 <= 4'h0;
    end
    if(reset) begin
      counts_987 <= 4'h0;
    end else if(T5971) begin
      counts_987 <= T52;
    end else if(io_resetCounts) begin
      counts_987 <= 4'h0;
    end
    if(reset) begin
      counts_988 <= 4'h0;
    end else if(T5979) begin
      counts_988 <= T52;
    end else if(io_resetCounts) begin
      counts_988 <= 4'h0;
    end
    if(reset) begin
      counts_989 <= 4'h0;
    end else if(T5983) begin
      counts_989 <= T52;
    end else if(io_resetCounts) begin
      counts_989 <= 4'h0;
    end
    if(reset) begin
      counts_990 <= 4'h0;
    end else if(T5989) begin
      counts_990 <= T52;
    end else if(io_resetCounts) begin
      counts_990 <= 4'h0;
    end
    if(reset) begin
      counts_991 <= 4'h0;
    end else if(T5993) begin
      counts_991 <= T52;
    end else if(io_resetCounts) begin
      counts_991 <= 4'h0;
    end
    if(reset) begin
      counts_992 <= 4'h0;
    end else if(T6007) begin
      counts_992 <= T52;
    end else if(io_resetCounts) begin
      counts_992 <= 4'h0;
    end
    if(reset) begin
      counts_993 <= 4'h0;
    end else if(T6011) begin
      counts_993 <= T52;
    end else if(io_resetCounts) begin
      counts_993 <= 4'h0;
    end
    if(reset) begin
      counts_994 <= 4'h0;
    end else if(T6017) begin
      counts_994 <= T52;
    end else if(io_resetCounts) begin
      counts_994 <= 4'h0;
    end
    if(reset) begin
      counts_995 <= 4'h0;
    end else if(T6021) begin
      counts_995 <= T52;
    end else if(io_resetCounts) begin
      counts_995 <= 4'h0;
    end
    if(reset) begin
      counts_996 <= 4'h0;
    end else if(T6029) begin
      counts_996 <= T52;
    end else if(io_resetCounts) begin
      counts_996 <= 4'h0;
    end
    if(reset) begin
      counts_997 <= 4'h0;
    end else if(T6033) begin
      counts_997 <= T52;
    end else if(io_resetCounts) begin
      counts_997 <= 4'h0;
    end
    if(reset) begin
      counts_998 <= 4'h0;
    end else if(T6039) begin
      counts_998 <= T52;
    end else if(io_resetCounts) begin
      counts_998 <= 4'h0;
    end
    if(reset) begin
      counts_999 <= 4'h0;
    end else if(T6043) begin
      counts_999 <= T52;
    end else if(io_resetCounts) begin
      counts_999 <= 4'h0;
    end
    if(reset) begin
      counts_1000 <= 4'h0;
    end else if(T6053) begin
      counts_1000 <= T52;
    end else if(io_resetCounts) begin
      counts_1000 <= 4'h0;
    end
    if(reset) begin
      counts_1001 <= 4'h0;
    end else if(T6057) begin
      counts_1001 <= T52;
    end else if(io_resetCounts) begin
      counts_1001 <= 4'h0;
    end
    if(reset) begin
      counts_1002 <= 4'h0;
    end else if(T6063) begin
      counts_1002 <= T52;
    end else if(io_resetCounts) begin
      counts_1002 <= 4'h0;
    end
    if(reset) begin
      counts_1003 <= 4'h0;
    end else if(T6067) begin
      counts_1003 <= T52;
    end else if(io_resetCounts) begin
      counts_1003 <= 4'h0;
    end
    if(reset) begin
      counts_1004 <= 4'h0;
    end else if(T6075) begin
      counts_1004 <= T52;
    end else if(io_resetCounts) begin
      counts_1004 <= 4'h0;
    end
    if(reset) begin
      counts_1005 <= 4'h0;
    end else if(T6079) begin
      counts_1005 <= T52;
    end else if(io_resetCounts) begin
      counts_1005 <= 4'h0;
    end
    if(reset) begin
      counts_1006 <= 4'h0;
    end else if(T6085) begin
      counts_1006 <= T52;
    end else if(io_resetCounts) begin
      counts_1006 <= 4'h0;
    end
    if(reset) begin
      counts_1007 <= 4'h0;
    end else if(T6089) begin
      counts_1007 <= T52;
    end else if(io_resetCounts) begin
      counts_1007 <= 4'h0;
    end
    if(reset) begin
      counts_1008 <= 4'h0;
    end else if(T6101) begin
      counts_1008 <= T52;
    end else if(io_resetCounts) begin
      counts_1008 <= 4'h0;
    end
    if(reset) begin
      counts_1009 <= 4'h0;
    end else if(T6105) begin
      counts_1009 <= T52;
    end else if(io_resetCounts) begin
      counts_1009 <= 4'h0;
    end
    if(reset) begin
      counts_1010 <= 4'h0;
    end else if(T6111) begin
      counts_1010 <= T52;
    end else if(io_resetCounts) begin
      counts_1010 <= 4'h0;
    end
    if(reset) begin
      counts_1011 <= 4'h0;
    end else if(T6115) begin
      counts_1011 <= T52;
    end else if(io_resetCounts) begin
      counts_1011 <= 4'h0;
    end
    if(reset) begin
      counts_1012 <= 4'h0;
    end else if(T6123) begin
      counts_1012 <= T52;
    end else if(io_resetCounts) begin
      counts_1012 <= 4'h0;
    end
    if(reset) begin
      counts_1013 <= 4'h0;
    end else if(T6127) begin
      counts_1013 <= T52;
    end else if(io_resetCounts) begin
      counts_1013 <= 4'h0;
    end
    if(reset) begin
      counts_1014 <= 4'h0;
    end else if(T6133) begin
      counts_1014 <= T52;
    end else if(io_resetCounts) begin
      counts_1014 <= 4'h0;
    end
    if(reset) begin
      counts_1015 <= 4'h0;
    end else if(T6137) begin
      counts_1015 <= T52;
    end else if(io_resetCounts) begin
      counts_1015 <= 4'h0;
    end
    if(reset) begin
      counts_1016 <= 4'h0;
    end else if(T6147) begin
      counts_1016 <= T52;
    end else if(io_resetCounts) begin
      counts_1016 <= 4'h0;
    end
    if(reset) begin
      counts_1017 <= 4'h0;
    end else if(T6151) begin
      counts_1017 <= T52;
    end else if(io_resetCounts) begin
      counts_1017 <= 4'h0;
    end
    if(reset) begin
      counts_1018 <= 4'h0;
    end else if(T6157) begin
      counts_1018 <= T52;
    end else if(io_resetCounts) begin
      counts_1018 <= 4'h0;
    end
    if(reset) begin
      counts_1019 <= 4'h0;
    end else if(T6161) begin
      counts_1019 <= T52;
    end else if(io_resetCounts) begin
      counts_1019 <= 4'h0;
    end
    if(reset) begin
      counts_1020 <= 4'h0;
    end else if(T6169) begin
      counts_1020 <= T52;
    end else if(io_resetCounts) begin
      counts_1020 <= 4'h0;
    end
    if(reset) begin
      counts_1021 <= 4'h0;
    end else if(T6173) begin
      counts_1021 <= T52;
    end else if(io_resetCounts) begin
      counts_1021 <= 4'h0;
    end
    if(reset) begin
      counts_1022 <= 4'h0;
    end else if(T6179) begin
      counts_1022 <= T52;
    end else if(io_resetCounts) begin
      counts_1022 <= 4'h0;
    end
    if(reset) begin
      counts_1023 <= 4'h0;
    end else if(T6183) begin
      counts_1023 <= T52;
    end else if(io_resetCounts) begin
      counts_1023 <= 4'h0;
    end
    if(reset) begin
      counts_1 <= 4'h0;
    end else if(T6200) begin
      counts_1 <= T52;
    end else if(io_resetCounts) begin
      counts_1 <= 4'h0;
    end
    if(reset) begin
      hashCount1 <= 4'h0;
    end else if(T21) begin
      hashCount1 <= T8240;
    end
    if(T10303) begin
      delayCount <= T10302;
    end else if(T22) begin
      delayCount <= 1'h1;
    end
    delayedIndex <= R10323;
    R10323 <= index;
    if(T10329) begin
      index <= T10328;
    end else if(T10303) begin
      index <= T10327;
    end else if(T22) begin
      index <= 6'h0;
    end
    if(T20) begin
      curInfo_tag <= io_hashIn_bits_tag;
    end
  end
endmodule

module KeyCopier(input clk, input reset,
    output[5:0] io_curKeyAddr,
    input [31:0] io_curKeyData,
    output[15:0] io_allKeyAddr,
    output[31:0] io_allKeyData,
    output io_allKeyWrite,
    output io_copyReq_ready,
    input  io_copyReq_valid,
    input [9:0] io_copyReq_bits_hash,
    input [7:0] io_copyReq_bits_len,
    output io_selCopy
);

  wire T0;
  reg  state;
  wire T23;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[7:0] nextlen;
  wire[7:0] T7;
  reg [7:0] len;
  wire[7:0] T8;
  wire[7:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[5:0] T13;
  wire T14;
  wire T15;
  reg  delayedWrite;
  reg  R16;
  wire write;
  wire[15:0] T17;
  reg [5:0] delayedIndex;
  reg [5:0] R18;
  reg [5:0] index;
  wire[5:0] T19;
  wire[5:0] T20;
  wire[5:0] T21;
  reg [9:0] hash;
  wire[9:0] T22;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    len = {1{$random}};
    delayedWrite = {1{$random}};
    R16 = {1{$random}};
    delayedIndex = {1{$random}};
    R18 = {1{$random}};
    index = {1{$random}};
    hash = {1{$random}};
  end
`endif

  assign io_selCopy = T0;
  assign T0 = state == 1'h1;
  assign T23 = reset ? 1'h0 : T1;
  assign T1 = T5 ? 1'h0 : T2;
  assign T2 = T3 ? 1'h1 : state;
  assign T3 = T4 & io_copyReq_valid;
  assign T4 = 1'h0 == state;
  assign T5 = T14 & T6;
  assign T6 = nextlen == 8'h0;
  assign nextlen = T12 ? 8'h0 : T7;
  assign T7 = len - 8'h4;
  assign T8 = T10 ? nextlen : T9;
  assign T9 = T3 ? io_copyReq_bits_len : len;
  assign T10 = T14 & T11;
  assign T11 = T6 ^ 1'h1;
  assign T12 = T13 == 6'h0;
  assign T13 = len[3'h7:2'h2];
  assign T14 = 1'h1 == state;
  assign io_copyReq_ready = T15;
  assign T15 = state == 1'h0;
  assign io_allKeyWrite = delayedWrite;
  assign write = state == 1'h1;
  assign io_allKeyData = io_curKeyData;
  assign io_allKeyAddr = T17;
  assign T17 = {hash, delayedIndex};
  assign T19 = T10 ? T21 : T20;
  assign T20 = T3 ? 6'h0 : index;
  assign T21 = index + 6'h1;
  assign T22 = T3 ? io_copyReq_bits_hash : hash;
  assign io_curKeyAddr = index;

  always @(posedge clk) begin
    if(reset) begin
      state <= 1'h0;
    end else if(T5) begin
      state <= 1'h0;
    end else if(T3) begin
      state <= 1'h1;
    end
    if(T10) begin
      len <= nextlen;
    end else if(T3) begin
      len <= io_copyReq_bits_len;
    end
    delayedWrite <= R16;
    R16 <= write;
    delayedIndex <= R18;
    R18 <= index;
    if(T10) begin
      index <= T21;
    end else if(T3) begin
      index <= 6'h0;
    end
    if(T3) begin
      hash <= io_copyReq_bits_hash;
    end
  end
endmodule

module UnbankedMem_0(input clk,
    input [6:0] io_readAddr,
    output[31:0] io_readData,
    input  io_readEn,
    input [6:0] io_writeAddr,
    input [31:0] io_writeData,
    input  io_writeEn
);

  reg [31:0] readDataReg;
  wire[31:0] T0;
  wire[31:0] readData;
  wire[31:0] T1;
  reg [31:0] writeDataReg;
  reg  writeEnReg;
  reg [6:0] writeAddrReg;
  reg [6:0] readAddrReg;
  wire[6:0] T2;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    readDataReg = {1{$random}};
    writeDataReg = {1{$random}};
    writeEnReg = {1{$random}};
    writeAddrReg = {1{$random}};
    readAddrReg = {1{$random}};
  end
`endif

  assign io_readData = readDataReg;
  assign T0 = io_readEn ? readData : readDataReg;
  UnbankedMem_mem mem (
    .CLK(clk),
    .W0A(writeAddrReg),
    .W0E(writeEnReg),
    .W0I(writeDataReg),
    .R1A(io_readAddr),
    .R1E(io_readEn),
    .R1O(readData)
  );
  assign T2 = io_readEn ? io_readAddr : readAddrReg;

  always @(posedge clk) begin
    if(io_readEn) begin
      readDataReg <= readData;
    end
    writeDataReg <= io_writeData;
    writeEnReg <= io_writeEn;
    writeAddrReg <= io_writeAddr;
    if(io_readEn) begin
      readAddrReg <= io_readAddr;
    end
  end
endmodule

module UnbankedMem_1(input clk,
    input [15:0] io_readAddr,
    output[31:0] io_readData,
    input  io_readEn,
    input [15:0] io_writeAddr,
    input [31:0] io_writeData,
    input  io_writeEn
);

  reg [31:0] readDataReg;
  wire[31:0] T0;
  wire[31:0] readData;
  wire[31:0] T1;
  reg [31:0] writeDataReg;
  reg  writeEnReg;
  reg [15:0] writeAddrReg;
  reg [15:0] readAddrReg;
  wire[15:0] T2;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    readDataReg = {1{$random}};
    writeDataReg = {1{$random}};
    writeEnReg = {1{$random}};
    writeAddrReg = {1{$random}};
    readAddrReg = {1{$random}};
  end
`endif

  assign io_readData = readDataReg;
  assign T0 = io_readEn ? readData : readDataReg;
  UnbankedMem_mem_1 mem (
    .CLK(clk),
    .W0A(writeAddrReg),
    .W0E(writeEnReg),
    .W0I(writeDataReg),
    .R1A(io_readAddr),
    .R1E(io_readEn),
    .R1O(readData)
  );
  assign T2 = io_readEn ? io_readAddr : readAddrReg;

  always @(posedge clk) begin
    if(io_readEn) begin
      readDataReg <= readData;
    end
    writeDataReg <= io_writeData;
    writeEnReg <= io_writeEn;
    writeAddrReg <= io_writeAddr;
    if(io_readEn) begin
      readAddrReg <= io_readAddr;
    end
  end
endmodule

module UnbankedMem_2(input clk,
    input [18:0] io_readAddr,
    output[7:0] io_readData,
    input  io_readEn,
    input [18:0] io_writeAddr,
    input [7:0] io_writeData,
    input  io_writeEn
);

  reg [7:0] readDataReg;
  wire[7:0] T0;
  wire[7:0] readData;
  wire[7:0] T1;
  reg [7:0] writeDataReg;
  reg  writeEnReg;
  reg [18:0] writeAddrReg;
  reg [18:0] readAddrReg;
  wire[18:0] T2;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    readDataReg = {1{$random}};
    writeDataReg = {1{$random}};
    writeEnReg = {1{$random}};
    writeAddrReg = {1{$random}};
    readAddrReg = {1{$random}};
  end
`endif

  assign io_readData = readDataReg;
  assign T0 = io_readEn ? readData : readDataReg;
  UnbankedMem_mem_2 mem (
    .CLK(clk),
    .W0A(writeAddrReg),
    .W0E(writeEnReg),
    .W0I(writeDataReg),
    .R1A(io_readAddr),
    .R1E(io_readEn),
    .R1O(readData)
  );
  assign T2 = io_readEn ? io_readAddr : readAddrReg;

  always @(posedge clk) begin
    if(io_readEn) begin
      readDataReg <= readData;
    end
    writeDataReg <= io_writeData;
    writeEnReg <= io_writeEn;
    writeAddrReg <= io_writeAddr;
    if(io_readEn) begin
      readAddrReg <= io_readAddr;
    end
  end
endmodule

module UnbankedMem_3(input clk,
    input [9:0] io_readAddr,
    output[18:0] io_readData,
    input  io_readEn,
    input [9:0] io_writeAddr,
    input [18:0] io_writeData,
    input  io_writeEn
);

  reg [18:0] readDataReg;
  wire[18:0] T0;
  wire[18:0] readData;
  wire[18:0] T1;
  reg [18:0] writeDataReg;
  reg  writeEnReg;
  reg [9:0] writeAddrReg;
  reg [9:0] readAddrReg;
  wire[9:0] T2;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    readDataReg = {1{$random}};
    writeDataReg = {1{$random}};
    writeEnReg = {1{$random}};
    writeAddrReg = {1{$random}};
    readAddrReg = {1{$random}};
  end
`endif

  assign io_readData = readDataReg;
  assign T0 = io_readEn ? readData : readDataReg;
  UnbankedMem_mem_3 mem (
    .CLK(clk),
    .W0A(writeAddrReg),
    .W0E(writeEnReg),
    .W0I(writeDataReg),
    .R1A(io_readAddr),
    .R1E(io_readEn),
    .R1O(readData)
  );
  assign T2 = io_readEn ? io_readAddr : readAddrReg;

  always @(posedge clk) begin
    if(io_readEn) begin
      readDataReg <= readData;
    end
    writeDataReg <= io_writeData;
    writeEnReg <= io_writeEn;
    writeAddrReg <= io_writeAddr;
    if(io_readEn) begin
      readAddrReg <= io_readAddr;
    end
  end
endmodule

module ValueCache(input clk, input reset,
    output io_hashIn_ready,
    input  io_hashIn_valid,
    input [3:0] io_hashIn_bits_tag,
    input [9:0] io_hashIn_bits_hash,
    input  io_hashIn_bits_found,
    input  io_resultInfo_ready,
    output io_resultInfo_valid,
    output[18:0] io_resultInfo_bits_len,
    output[3:0] io_resultInfo_bits_tag,
    input  io_resultData_ready,
    output io_resultData_valid,
    output[7:0] io_resultData_bits,
    input [18:0] io_cacheWriteAddr,
    input [7:0] io_cacheWriteData,
    input  io_cacheWriteEn,
    input [9:0] io_addrLenAddr,
    input [18:0] io_addrLenWriteData_addr,
    input [18:0] io_addrLenWriteData_len,
    input  io_addrLenWriteEn_1,
    input  io_addrLenWriteEn_0,
    output[18:0] io_addrLenReadData_addr,
    output[18:0] io_addrLenReadData_len,
    input  io_addrLenReadEn
);

  wire[9:0] realAddrLenAddr;
  reg [9:0] addrLenAddr;
  wire[9:0] T53;
  wire T9;
  wire T10;
  wire T11;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  delayCount;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg [18:0] len;
  wire[18:0] T37;
  wire[18:0] T38;
  wire[18:0] T39;
  wire[18:0] T40;
  wire[18:0] addrLenData_len;
  wire[18:0] T41;
  wire[18:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg  cacheReadEn;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  reg [18:0] cacheAddr;
  wire[18:0] T60;
  wire[18:0] T61;
  wire[18:0] T62;
  wire[18:0] addrLenData_addr;
  wire[18:0] T63;
  wire[18:0] T64;
  wire T0;
  reg [3:0] tag;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[7:0] cacheMem_io_readData;
  wire[18:0] addrTable_io_readData;
  wire[18:0] lenTable_io_readData;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    addrLenAddr = {1{$random}};
    state = {1{$random}};
    delayCount = {1{$random}};
    len = {1{$random}};
    cacheReadEn = {1{$random}};
    cacheAddr = {1{$random}};
    tag = {1{$random}};
  end
`endif

  assign realAddrLenAddr = io_addrLenReadEn ? io_addrLenAddr : addrLenAddr;
  assign T53 = T9 ? io_hashIn_bits_hash : addrLenAddr;
  assign T9 = T10 & io_hashIn_bits_found;
  assign T10 = T11 & io_hashIn_valid;
  assign T11 = 3'h0 == state;
  assign T52 = reset ? 3'h0 : T1;
  assign T1 = T35 ? 3'h0 : T2;
  assign T2 = T34 ? 3'h6 : T3;
  assign T3 = T32 ? 3'h5 : T4;
  assign T4 = T31 ? 3'h4 : T5;
  assign T5 = T16 ? 3'h3 : T6;
  assign T6 = T14 ? 3'h0 : T7;
  assign T7 = T12 ? 3'h1 : T8;
  assign T8 = T9 ? 3'h2 : state;
  assign T12 = T10 & T13;
  assign T13 = io_hashIn_bits_found ^ 1'h1;
  assign T14 = T15 & io_resultInfo_ready;
  assign T15 = 3'h1 == state;
  assign T16 = T30 & T17;
  assign T17 = delayCount == 1'h0;
  assign T18 = T26 ? T25 : T19;
  assign T19 = T32 ? 1'h1 : T20;
  assign T20 = T23 ? T22 : T21;
  assign T21 = T9 ? 1'h1 : delayCount;
  assign T22 = delayCount - 1'h1;
  assign T23 = T30 & T24;
  assign T24 = T17 ^ 1'h1;
  assign T25 = delayCount - 1'h1;
  assign T26 = T29 & T27;
  assign T27 = T28 ^ 1'h1;
  assign T28 = delayCount == 1'h0;
  assign T29 = 3'h5 == state;
  assign T30 = 3'h2 == state;
  assign T31 = 3'h3 == state;
  assign T32 = T33 & io_resultInfo_ready;
  assign T33 = 3'h4 == state;
  assign T34 = T29 & T28;
  assign T35 = T45 & T36;
  assign T36 = len == 19'h0;
  assign T37 = T43 ? T42 : T38;
  assign T38 = T34 ? T41 : T39;
  assign T39 = T31 ? addrLenData_len : T40;
  assign T40 = T12 ? 19'h0 : len;
  assign addrLenData_len = lenTable_io_readData;
  assign T41 = len - 19'h1;
  assign T42 = len - 19'h1;
  assign T43 = T45 & T44;
  assign T44 = T36 ^ 1'h1;
  assign T45 = T46 & io_resultData_ready;
  assign T46 = 3'h6 == state;
  assign T54 = reset ? 1'h0 : T55;
  assign T55 = T43 ? 1'h1 : T56;
  assign T56 = T35 ? 1'h0 : T57;
  assign T57 = T46 ? 1'h0 : T58;
  assign T58 = T29 ? 1'h1 : T59;
  assign T59 = T32 ? 1'h1 : cacheReadEn;
  assign T60 = T43 ? T64 : T61;
  assign T61 = T29 ? T63 : T62;
  assign T62 = T31 ? addrLenData_addr : cacheAddr;
  assign addrLenData_addr = addrTable_io_readData;
  assign T63 = cacheAddr + 19'h1;
  assign T64 = cacheAddr + 19'h1;
  assign io_addrLenReadData_len = lenTable_io_readData;
  assign io_addrLenReadData_addr = addrTable_io_readData;
  assign io_resultData_bits = cacheMem_io_readData;
  assign io_resultData_valid = T0;
  assign T0 = state == 3'h6;
  assign io_resultInfo_bits_tag = tag;
  assign T47 = T10 ? io_hashIn_bits_tag : tag;
  assign io_resultInfo_bits_len = len;
  assign io_resultInfo_valid = T48;
  assign T48 = T50 | T49;
  assign T49 = state == 3'h1;
  assign T50 = state == 3'h4;
  assign io_hashIn_ready = T51;
  assign T51 = state == 3'h0;
  UnbankedMem_2 cacheMem(.clk(clk),
       .io_readAddr( cacheAddr ),
       .io_readData( cacheMem_io_readData ),
       .io_readEn( cacheReadEn ),
       .io_writeAddr( io_cacheWriteAddr ),
       .io_writeData( io_cacheWriteData ),
       .io_writeEn( io_cacheWriteEn )
  );
  UnbankedMem_3 addrTable(.clk(clk),
       .io_readAddr( realAddrLenAddr ),
       .io_readData( addrTable_io_readData ),
       .io_readEn( 1'h1 ),
       .io_writeAddr( io_addrLenAddr ),
       .io_writeData( io_addrLenWriteData_addr ),
       .io_writeEn( io_addrLenWriteEn_0 )
  );
  UnbankedMem_3 lenTable(.clk(clk),
       .io_readAddr( realAddrLenAddr ),
       .io_readData( lenTable_io_readData ),
       .io_readEn( 1'h1 ),
       .io_writeAddr( io_addrLenAddr ),
       .io_writeData( io_addrLenWriteData_len ),
       .io_writeEn( io_addrLenWriteEn_1 )
  );

  always @(posedge clk) begin
    if(T9) begin
      addrLenAddr <= io_hashIn_bits_hash;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h6;
    end else if(T32) begin
      state <= 3'h5;
    end else if(T31) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= 3'h3;
    end else if(T14) begin
      state <= 3'h0;
    end else if(T12) begin
      state <= 3'h1;
    end else if(T9) begin
      state <= 3'h2;
    end
    if(T26) begin
      delayCount <= T25;
    end else if(T32) begin
      delayCount <= 1'h1;
    end else if(T23) begin
      delayCount <= T22;
    end else if(T9) begin
      delayCount <= 1'h1;
    end
    if(T43) begin
      len <= T42;
    end else if(T34) begin
      len <= T41;
    end else if(T31) begin
      len <= addrLenData_len;
    end else if(T12) begin
      len <= 19'h0;
    end
    if(reset) begin
      cacheReadEn <= 1'h0;
    end else if(T43) begin
      cacheReadEn <= 1'h1;
    end else if(T35) begin
      cacheReadEn <= 1'h0;
    end else if(T46) begin
      cacheReadEn <= 1'h0;
    end else if(T29) begin
      cacheReadEn <= 1'h1;
    end else if(T32) begin
      cacheReadEn <= 1'h1;
    end
    if(T43) begin
      cacheAddr <= T64;
    end else if(T29) begin
      cacheAddr <= T63;
    end else if(T31) begin
      cacheAddr <= addrLenData_addr;
    end
    if(T10) begin
      tag <= io_hashIn_bits_tag;
    end
  end
endmodule

module LookupPipeline(input clk, input reset,
    input  io_lock,
    output io_halted,
    input  io_writemode,
    input  io_findAvailable,
    input  io_resetCounts,
    output io_readKeyInfo_ready,
    input  io_readKeyInfo_valid,
    input [7:0] io_readKeyInfo_bits_len,
    input [3:0] io_readKeyInfo_bits_tag,
    output io_readKeyData_ready,
    input  io_readKeyData_valid,
    input [7:0] io_readKeyData_bits,
    output io_writeKeyInfo_ready,
    input  io_writeKeyInfo_valid,
    input [7:0] io_writeKeyInfo_bits_len,
    input [3:0] io_writeKeyInfo_bits_tag,
    output io_writeKeyData_ready,
    input  io_writeKeyData_valid,
    input [7:0] io_writeKeyData_bits,
    input  io_hashSel_ready,
    output io_hashSel_valid,
    output[3:0] io_hashSel_bits_tag,
    output[9:0] io_hashSel_bits_hash,
    output io_hashSel_bits_found,
    output io_copyReq_ready,
    input  io_copyReq_valid,
    input [9:0] io_copyReq_bits_hash,
    input [7:0] io_copyReq_bits_len,
    input  io_resultInfo_ready,
    output io_resultInfo_valid,
    output[18:0] io_resultInfo_bits_len,
    output[3:0] io_resultInfo_bits_tag,
    input  io_resultData_ready,
    output io_resultData_valid,
    output[7:0] io_resultData_bits,
    input [18:0] io_cacheWriteAddr,
    input [7:0] io_cacheWriteData,
    input  io_cacheWriteEn,
    input [9:0] io_addrLenAddr,
    input [18:0] io_addrLenWriteData_addr,
    input [18:0] io_addrLenWriteData_len,
    input  io_addrLenWriteEn_1,
    input  io_addrLenWriteEn_0,
    output[18:0] io_addrLenReadData_addr,
    output[18:0] io_addrLenReadData_len,
    input  io_addrLenReadEn,
    input [9:0] io_keyLenAddr,
    input [7:0] io_keyLenData,
    input  io_keyLenWrite
);

  wire T9;
  wire T10;
  wire[6:0] hwWriteAddr;
  reg  swapped;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire[6:0] curReadAddrExt;
  wire[5:0] curReadAddrRaw;
  wire T15;
  wire T16;
  wire[7:0] T17;
  wire[7:0] T18;
  reg [9:0] lenAddr;
  wire[3:0] T19;
  wire[7:0] T20;
  wire T21;
  wire[7:0] T22;
  wire T23;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[5:0] keycompare_io_curKeyAddr;
  wire[15:0] keycompare_io_allKeyAddr;
  wire[9:0] keycompare_io_lenAddr;
  wire keycompare_io_hashIn_ready;
  wire keycompare_io_hashOut_valid;
  wire[3:0] keycompare_io_hashOut_bits_tag;
  wire[9:0] keycompare_io_hashOut_bits_hash;
  wire keycompare_io_hashOut_bits_found;
  wire[5:0] keycopy_io_curKeyAddr;
  wire[15:0] keycopy_io_allKeyAddr;
  wire[31:0] keycopy_io_allKeyData;
  wire keycopy_io_allKeyWrite;
  wire keycopy_io_copyReq_ready;
  wire keycopy_io_selCopy;
  wire[31:0] curKeyMem_io_readData;
  wire[31:0] allKeyMem_io_readData;
  wire[5:0] hasherwriter_io_keyWriteAddr;
  wire[31:0] hasherwriter_io_keyWriteData;
  wire hasherwriter_io_keyWrite;
  wire hasherwriter_io_keyData_ready;
  wire hasherwriter_io_keyInfo_ready;
  wire hasherwriter_io_hashOut_valid;
  wire[9:0] hasherwriter_io_hashOut_bits_hash1;
  wire[9:0] hasherwriter_io_hashOut_bits_hash2;
  wire[7:0] hasherwriter_io_hashOut_bits_len;
  wire[3:0] hasherwriter_io_hashOut_bits_tag;
  wire hasherwriter_io_halted;
  wire valcache_io_hashIn_ready;
  wire valcache_io_resultInfo_valid;
  wire[18:0] valcache_io_resultInfo_bits_len;
  wire[3:0] valcache_io_resultInfo_bits_tag;
  wire valcache_io_resultData_valid;
  wire[7:0] valcache_io_resultData_bits;
  wire[18:0] valcache_io_addrLenReadData_addr;
  wire[18:0] valcache_io_addrLenReadData_len;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    swapped = {1{$random}};
    lenAddr = {1{$random}};
  end
`endif

  assign T9 = keycompare_io_hashOut_valid & T10;
  assign T10 = io_writemode ^ 1'h1;
  assign hwWriteAddr = {swapped, hasherwriter_io_keyWriteAddr};
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = T14 ? T13 : swapped;
  assign T13 = swapped ^ 1'h1;
  assign T14 = hasherwriter_io_hashOut_valid & keycompare_io_hashIn_ready;
  assign curReadAddrExt = {T15, curReadAddrRaw};
  assign curReadAddrRaw = keycopy_io_selCopy ? keycopy_io_curKeyAddr : keycompare_io_curKeyAddr;
  assign T15 = swapped ^ 1'h1;
  assign T16 = io_writemode ? io_hashSel_ready : valcache_io_hashIn_ready;
  LookupPipeline_lenMem lenMem (
    .CLK(clk),
    .W0A(io_keyLenAddr),
    .W0E(io_keyLenWrite),
    .W0I(io_keyLenData),
    .R1A(keycompare_io_lenAddr),
    .R1E(1'h1),
    .R1O(T17)
  );
  assign T19 = io_writemode ? io_writeKeyInfo_bits_tag : io_readKeyInfo_bits_tag;
  assign T20 = io_writemode ? io_writeKeyInfo_bits_len : io_readKeyInfo_bits_len;
  assign T21 = io_writemode ? io_writeKeyInfo_valid : io_readKeyInfo_valid;
  assign T22 = io_writemode ? io_writeKeyData_bits : io_readKeyData_bits;
  assign T23 = io_writemode ? io_writeKeyData_valid : io_readKeyData_valid;
  assign io_addrLenReadData_len = valcache_io_addrLenReadData_len;
  assign io_addrLenReadData_addr = valcache_io_addrLenReadData_addr;
  assign io_resultData_bits = valcache_io_resultData_bits;
  assign io_resultData_valid = valcache_io_resultData_valid;
  assign io_resultInfo_bits_tag = valcache_io_resultInfo_bits_tag;
  assign io_resultInfo_bits_len = valcache_io_resultInfo_bits_len;
  assign io_resultInfo_valid = valcache_io_resultInfo_valid;
  assign io_copyReq_ready = keycopy_io_copyReq_ready;
  assign io_hashSel_bits_found = keycompare_io_hashOut_bits_found;
  assign io_hashSel_bits_hash = keycompare_io_hashOut_bits_hash;
  assign io_hashSel_bits_tag = keycompare_io_hashOut_bits_tag;
  assign io_hashSel_valid = T0;
  assign T0 = keycompare_io_hashOut_valid & io_writemode;
  assign io_writeKeyData_ready = T1;
  assign T1 = hasherwriter_io_keyData_ready & io_writemode;
  assign io_writeKeyInfo_ready = T2;
  assign T2 = hasherwriter_io_keyInfo_ready & io_writemode;
  assign io_readKeyData_ready = T3;
  assign T3 = hasherwriter_io_keyData_ready & T4;
  assign T4 = io_writemode ^ 1'h1;
  assign io_readKeyInfo_ready = T5;
  assign T5 = hasherwriter_io_keyInfo_ready & T6;
  assign T6 = io_writemode ^ 1'h1;
  assign io_halted = T7;
  assign T7 = T8 & valcache_io_hashIn_ready;
  assign T8 = hasherwriter_io_halted & keycompare_io_hashIn_ready;
  HasherWriter hasherwriter(.clk(clk), .reset(reset),
       .io_keyWriteAddr( hasherwriter_io_keyWriteAddr ),
       .io_keyWriteData( hasherwriter_io_keyWriteData ),
       .io_keyWrite( hasherwriter_io_keyWrite ),
       .io_keyData_ready( hasherwriter_io_keyData_ready ),
       .io_keyData_valid( T23 ),
       .io_keyData_bits( T22 ),
       .io_keyInfo_ready( hasherwriter_io_keyInfo_ready ),
       .io_keyInfo_valid( T21 ),
       .io_keyInfo_bits_len( T20 ),
       .io_keyInfo_bits_tag( T19 ),
       .io_hashOut_ready( keycompare_io_hashIn_ready ),
       .io_hashOut_valid( hasherwriter_io_hashOut_valid ),
       .io_hashOut_bits_hash1( hasherwriter_io_hashOut_bits_hash1 ),
       .io_hashOut_bits_hash2( hasherwriter_io_hashOut_bits_hash2 ),
       .io_hashOut_bits_len( hasherwriter_io_hashOut_bits_len ),
       .io_hashOut_bits_tag( hasherwriter_io_hashOut_bits_tag ),
       .io_lock( io_lock ),
       .io_halted( hasherwriter_io_halted )
  );
  KeyCompare keycompare(.clk(clk), .reset(reset),
       .io_curKeyAddr( keycompare_io_curKeyAddr ),
       .io_curKeyData( curKeyMem_io_readData ),
       .io_allKeyAddr( keycompare_io_allKeyAddr ),
       .io_allKeyData( allKeyMem_io_readData ),
       .io_lenAddr( keycompare_io_lenAddr ),
       .io_lenData( T17 ),
       .io_hashIn_ready( keycompare_io_hashIn_ready ),
       .io_hashIn_valid( hasherwriter_io_hashOut_valid ),
       .io_hashIn_bits_hash1( hasherwriter_io_hashOut_bits_hash1 ),
       .io_hashIn_bits_hash2( hasherwriter_io_hashOut_bits_hash2 ),
       .io_hashIn_bits_len( hasherwriter_io_hashOut_bits_len ),
       .io_hashIn_bits_tag( hasherwriter_io_hashOut_bits_tag ),
       .io_hashOut_ready( T16 ),
       .io_hashOut_valid( keycompare_io_hashOut_valid ),
       .io_hashOut_bits_tag( keycompare_io_hashOut_bits_tag ),
       .io_hashOut_bits_hash( keycompare_io_hashOut_bits_hash ),
       .io_hashOut_bits_found( keycompare_io_hashOut_bits_found ),
       .io_findAvailable( io_findAvailable ),
       .io_resetCounts( io_resetCounts )
  );
  KeyCopier keycopy(.clk(clk), .reset(reset),
       .io_curKeyAddr( keycopy_io_curKeyAddr ),
       .io_curKeyData( curKeyMem_io_readData ),
       .io_allKeyAddr( keycopy_io_allKeyAddr ),
       .io_allKeyData( keycopy_io_allKeyData ),
       .io_allKeyWrite( keycopy_io_allKeyWrite ),
       .io_copyReq_ready( keycopy_io_copyReq_ready ),
       .io_copyReq_valid( io_copyReq_valid ),
       .io_copyReq_bits_hash( io_copyReq_bits_hash ),
       .io_copyReq_bits_len( io_copyReq_bits_len ),
       .io_selCopy( keycopy_io_selCopy )
  );
  UnbankedMem_0 curKeyMem(.clk(clk),
       .io_readAddr( curReadAddrExt ),
       .io_readData( curKeyMem_io_readData ),
       .io_readEn( 1'h1 ),
       .io_writeAddr( hwWriteAddr ),
       .io_writeData( hasherwriter_io_keyWriteData ),
       .io_writeEn( hasherwriter_io_keyWrite )
  );
  UnbankedMem_1 allKeyMem(.clk(clk),
       .io_readAddr( keycompare_io_allKeyAddr ),
       .io_readData( allKeyMem_io_readData ),
       .io_readEn( 1'h1 ),
       .io_writeAddr( keycopy_io_allKeyAddr ),
       .io_writeData( keycopy_io_allKeyData ),
       .io_writeEn( keycopy_io_allKeyWrite )
  );
  ValueCache valcache(.clk(clk), .reset(reset),
       .io_hashIn_ready( valcache_io_hashIn_ready ),
       .io_hashIn_valid( T9 ),
       .io_hashIn_bits_tag( keycompare_io_hashOut_bits_tag ),
       .io_hashIn_bits_hash( keycompare_io_hashOut_bits_hash ),
       .io_hashIn_bits_found( keycompare_io_hashOut_bits_found ),
       .io_resultInfo_ready( io_resultInfo_ready ),
       .io_resultInfo_valid( valcache_io_resultInfo_valid ),
       .io_resultInfo_bits_len( valcache_io_resultInfo_bits_len ),
       .io_resultInfo_bits_tag( valcache_io_resultInfo_bits_tag ),
       .io_resultData_ready( io_resultData_ready ),
       .io_resultData_valid( valcache_io_resultData_valid ),
       .io_resultData_bits( valcache_io_resultData_bits ),
       .io_cacheWriteAddr( io_cacheWriteAddr ),
       .io_cacheWriteData( io_cacheWriteData ),
       .io_cacheWriteEn( io_cacheWriteEn ),
       .io_addrLenAddr( io_addrLenAddr ),
       .io_addrLenWriteData_addr( io_addrLenWriteData_addr ),
       .io_addrLenWriteData_len( io_addrLenWriteData_len ),
       .io_addrLenWriteEn_1( io_addrLenWriteEn_1 ),
       .io_addrLenWriteEn_0( io_addrLenWriteEn_0 ),
       .io_addrLenReadData_addr( valcache_io_addrLenReadData_addr ),
       .io_addrLenReadData_len( valcache_io_addrLenReadData_len ),
       .io_addrLenReadEn( io_addrLenReadEn )
  );

  always @(posedge clk) begin
    if(reset) begin
      swapped <= 1'h0;
    end else if(T14) begin
      swapped <= T13;
    end
    lenAddr <= keycompare_io_lenAddr;
  end
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [7:0] io_enq_bits_len,
    input [3:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[7:0] io_deq_bits_len,
    output[3:0] io_deq_bits_tag
);

  wire[3:0] T0;
  wire[11:0] T1;
  reg [11:0] ram [1:0];
  wire[11:0] T2;
  wire[11:0] T3;
  wire[11:0] T4;
  wire do_enq;
  reg  R5;
  wire T17;
  wire T6;
  wire T7;
  reg  R8;
  wire T18;
  wire T9;
  wire T10;
  wire do_deq;
  wire[7:0] T11;
  wire T12;
  wire empty;
  wire T13;
  reg  maybe_full;
  wire T19;
  wire T14;
  wire T15;
  wire ptr_match;
  wire T16;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R5 = {1{$random}};
    R8 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[R8];
  assign T3 = T4;
  assign T4 = {io_enq_bits_len, io_enq_bits_tag};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T17 = reset ? 1'h0 : T6;
  assign T6 = do_enq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign T18 = reset ? 1'h0 : T9;
  assign T9 = do_deq ? T10 : R8;
  assign T10 = R8 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_len = T11;
  assign T11 = T1[4'hb:3'h4];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign T19 = reset ? 1'h0 : T14;
  assign T14 = T15 ? do_enq : maybe_full;
  assign T15 = do_enq != do_deq;
  assign ptr_match = R5 == R8;
  assign io_enq_ready = T16;
  assign T16 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R5] <= T3;
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_enq) begin
      R5 <= T7;
    end
    if(reset) begin
      R8 <= 1'h0;
    end else if(do_deq) begin
      R8 <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T15) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [7:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[7:0] io_deq_bits
);

  wire[7:0] T0;
  reg [7:0] ram [1:0];
  wire[7:0] T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [18:0] io_enq_bits_len,
    input [3:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[18:0] io_deq_bits_len,
    output[3:0] io_deq_bits_tag
);

  wire[3:0] T0;
  wire[22:0] T1;
  reg [22:0] ram [1:0];
  wire[22:0] T2;
  wire[22:0] T3;
  wire[22:0] T4;
  wire do_enq;
  reg  R5;
  wire T17;
  wire T6;
  wire T7;
  reg  R8;
  wire T18;
  wire T9;
  wire T10;
  wire do_deq;
  wire[18:0] T11;
  wire T12;
  wire empty;
  wire T13;
  reg  maybe_full;
  wire T19;
  wire T14;
  wire T15;
  wire ptr_match;
  wire T16;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R5 = {1{$random}};
    R8 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[R8];
  assign T3 = T4;
  assign T4 = {io_enq_bits_len, io_enq_bits_tag};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T17 = reset ? 1'h0 : T6;
  assign T6 = do_enq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign T18 = reset ? 1'h0 : T9;
  assign T9 = do_deq ? T10 : R8;
  assign T10 = R8 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_len = T11;
  assign T11 = T1[5'h16:3'h4];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign T19 = reset ? 1'h0 : T14;
  assign T14 = T15 ? do_enq : maybe_full;
  assign T15 = do_enq != do_deq;
  assign ptr_match = R5 == R8;
  assign io_enq_ready = T16;
  assign T16 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R5] <= T3;
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_enq) begin
      R5 <= T7;
    end
    if(reset) begin
      R8 <= 1'h0;
    end else if(do_deq) begin
      R8 <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T15) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module MemoryHandler(input clk, input reset,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[42:0] io_mem_req_bits_addr,
    //output[63:0] io_mem_req_bits_data
    //output[8:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [8:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [42:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input  io_keyData_ready,
    output io_keyData_valid,
    output[7:0] io_keyData_bits,
    output[18:0] io_cacheWriteAddr,
    output[7:0] io_cacheWriteData,
    output io_cacheWriteEn,
    output io_cmd_ready,
    input  io_cmd_valid,
    input  io_cmd_bits_action,
    input [63:0] io_cmd_bits_readstart,
    input [18:0] io_cmd_bits_writestart,
    input [63:0] io_cmd_bits_len
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T55;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[18:0] T19;
  reg [18:0] len;
  wire[18:0] T56;
  wire[63:0] T20;
  wire[63:0] T57;
  reg [18:0] bytesread;
  wire[18:0] T21;
  wire[18:0] T22;
  wire[18:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[2:0] byteOff;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg [1:0] outputMask;
  wire[1:0] T37;
  wire[1:0] T38;
  wire shifting;
  wire[7:0] T39;
  reg [63:0] word;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[63:0] T42;
  wire[55:0] T43;
  reg [18:0] writeaddr;
  wire[18:0] T44;
  wire[18:0] T45;
  wire[18:0] T46;
  wire[7:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[42:0] T58;
  reg [63:0] readaddr;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire T54;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    len = {1{$random}};
    bytesread = {1{$random}};
    outputMask = {1{$random}};
    word = {2{$random}};
    writeaddr = {1{$random}};
    readaddr = {2{$random}};
  end
`endif

  assign io_cmd_ready = T0;
  assign T0 = state == 3'h0;
  assign T55 = reset ? 3'h0 : T1;
  assign T1 = T33 ? 3'h0 : T2;
  assign T2 = T31 ? 3'h2 : T3;
  assign T3 = T29 ? 3'h4 : T4;
  assign T4 = T25 ? 3'h3 : T5;
  assign T5 = T17 ? 3'h5 : T6;
  assign T6 = T15 ? 3'h3 : T7;
  assign T7 = T13 ? 3'h3 : T8;
  assign T8 = T9 ? 3'h1 : state;
  assign T9 = T11 & T10;
  assign T10 = 1'h0 == io_cmd_bits_action;
  assign T11 = T12 & io_cmd_valid;
  assign T12 = 3'h0 == state;
  assign T13 = T11 & T14;
  assign T14 = 1'h1 == io_cmd_bits_action;
  assign T15 = T16 & io_keyData_ready;
  assign T16 = 3'h1 == state;
  assign T17 = T24 & T18;
  assign T18 = bytesread == T19;
  assign T19 = len - 19'h1;
  assign T56 = T20[5'h12:1'h0];
  assign T20 = T11 ? io_cmd_bits_len : T57;
  assign T57 = {45'h0, len};
  assign T21 = T24 ? T23 : T22;
  assign T22 = T11 ? 19'h0 : bytesread;
  assign T23 = bytesread + 19'h1;
  assign T24 = 3'h2 == state;
  assign T25 = T24 & T26;
  assign T26 = T28 & T27;
  assign T27 = byteOff == 3'h7;
  assign byteOff = bytesread[2'h2:1'h0];
  assign T28 = T18 ^ 1'h1;
  assign T29 = T30 & io_mem_req_ready;
  assign T30 = 3'h3 == state;
  assign T31 = T32 & io_mem_resp_valid;
  assign T32 = 3'h4 == state;
  assign T33 = 3'h5 == state;
  assign io_cacheWriteEn = T34;
  assign T34 = shifting & T35;
  assign T35 = T36;
  assign T36 = outputMask[1'h1:1'h1];
  assign T37 = T13 ? 2'h2 : T38;
  assign T38 = T9 ? 2'h1 : outputMask;
  assign shifting = state == 3'h2;
  assign io_cacheWriteData = T39;
  assign T39 = word[3'h7:1'h0];
  assign T40 = T31 ? io_mem_resp_bits_data : T41;
  assign T41 = T24 ? T42 : word;
  assign T42 = {8'h0, T43};
  assign T43 = word[6'h3f:4'h8];
  assign io_cacheWriteAddr = writeaddr;
  assign T44 = T24 ? T46 : T45;
  assign T45 = T11 ? io_cmd_bits_writestart : writeaddr;
  assign T46 = writeaddr + 19'h1;
  assign io_keyData_bits = T47;
  assign T47 = word[3'h7:1'h0];
  assign io_keyData_valid = T48;
  assign T48 = shifting & T49;
  assign T49 = T50;
  assign T50 = outputMask[1'h0:1'h0];
  assign io_mem_req_bits_cmd = 5'h0;
  assign io_mem_req_bits_addr = T58;
  assign T58 = readaddr[6'h2a:1'h0];
  assign T51 = T29 ? T53 : T52;
  assign T52 = T11 ? io_cmd_bits_readstart : readaddr;
  assign T53 = readaddr + 64'h8;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T54;
  assign T54 = state == 3'h3;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T33) begin
      state <= 3'h0;
    end else if(T31) begin
      state <= 3'h2;
    end else if(T29) begin
      state <= 3'h4;
    end else if(T25) begin
      state <= 3'h3;
    end else if(T17) begin
      state <= 3'h5;
    end else if(T15) begin
      state <= 3'h3;
    end else if(T13) begin
      state <= 3'h3;
    end else if(T9) begin
      state <= 3'h1;
    end
    len <= T56;
    if(T24) begin
      bytesread <= T23;
    end else if(T11) begin
      bytesread <= 19'h0;
    end
    if(T13) begin
      outputMask <= 2'h2;
    end else if(T9) begin
      outputMask <= 2'h1;
    end
    if(T31) begin
      word <= io_mem_resp_bits_data;
    end else if(T24) begin
      word <= T42;
    end
    if(T24) begin
      writeaddr <= T46;
    end else if(T11) begin
      writeaddr <= io_cmd_bits_writestart;
    end
    if(T29) begin
      readaddr <= T53;
    end else if(T11) begin
      readaddr <= io_cmd_bits_readstart;
    end
  end
endmodule

module CtrlModule(input clk, input reset,
    output io_rocc_cmd_ready,
    input  io_rocc_cmd_valid,
    input [6:0] io_rocc_cmd_bits_inst_funct,
    input [4:0] io_rocc_cmd_bits_inst_rs2,
    input [4:0] io_rocc_cmd_bits_inst_rs1,
    input  io_rocc_cmd_bits_inst_xd,
    input  io_rocc_cmd_bits_inst_xs1,
    input  io_rocc_cmd_bits_inst_xs2,
    input [4:0] io_rocc_cmd_bits_inst_rd,
    input [6:0] io_rocc_cmd_bits_inst_opcode,
    input [63:0] io_rocc_cmd_bits_rs1,
    input [63:0] io_rocc_cmd_bits_rs2,
    input  io_rocc_resp_ready,
    output io_rocc_resp_valid,
    output[4:0] io_rocc_resp_bits_rd,
    output[63:0] io_rocc_resp_bits_data,
    input  io_rocc_mem_req_ready,
    output io_rocc_mem_req_valid,
    output io_rocc_mem_req_bits_kill,
    output[2:0] io_rocc_mem_req_bits_typ,
    output io_rocc_mem_req_bits_phys,
    output[42:0] io_rocc_mem_req_bits_addr,
    //output[63:0] io_rocc_mem_req_bits_data
    //output[8:0] io_rocc_mem_req_bits_tag
    output[4:0] io_rocc_mem_req_bits_cmd,
    input  io_rocc_mem_resp_valid,
    input  io_rocc_mem_resp_bits_nack,
    input  io_rocc_mem_resp_bits_replay,
    input [2:0] io_rocc_mem_resp_bits_typ,
    input  io_rocc_mem_resp_bits_has_data,
    input [63:0] io_rocc_mem_resp_bits_data,
    input [63:0] io_rocc_mem_resp_bits_data_subword,
    input [8:0] io_rocc_mem_resp_bits_tag,
    input [3:0] io_rocc_mem_resp_bits_cmd,
    input [42:0] io_rocc_mem_resp_bits_addr,
    input [63:0] io_rocc_mem_resp_bits_store_data,
    input  io_rocc_mem_replay_next_valid,
    input [8:0] io_rocc_mem_replay_next_bits,
    input  io_rocc_mem_xcpt_ma_ld,
    input  io_rocc_mem_xcpt_ma_st,
    input  io_rocc_mem_xcpt_pf_ld,
    input  io_rocc_mem_xcpt_pf_st,
    //output io_rocc_mem_ptw_req_ready
    input  io_rocc_mem_ptw_req_valid,
    input [29:0] io_rocc_mem_ptw_req_bits,
    //output io_rocc_mem_ptw_resp_valid
    //output io_rocc_mem_ptw_resp_bits_error
    //output[18:0] io_rocc_mem_ptw_resp_bits_ppn
    //output[5:0] io_rocc_mem_ptw_resp_bits_perm
    //output[7:0] io_rocc_mem_ptw_status_ip
    //output[7:0] io_rocc_mem_ptw_status_im
    //output[6:0] io_rocc_mem_ptw_status_zero
    //output io_rocc_mem_ptw_status_er
    //output io_rocc_mem_ptw_status_vm
    //output io_rocc_mem_ptw_status_s64
    //output io_rocc_mem_ptw_status_u64
    //output io_rocc_mem_ptw_status_ef
    //output io_rocc_mem_ptw_status_pei
    //output io_rocc_mem_ptw_status_ei
    //output io_rocc_mem_ptw_status_ps
    //output io_rocc_mem_ptw_status_s
    //output io_rocc_mem_ptw_invalidate
    //output io_rocc_mem_ptw_sret
    input  io_rocc_mem_ordered,
    output io_rocc_busy,
    input  io_rocc_s,
    output io_rocc_interrupt,
    input  io_rocc_imem_acquire_ready,
    output io_rocc_imem_acquire_valid,
    //output[1:0] io_rocc_imem_acquire_bits_header_src
    //output[1:0] io_rocc_imem_acquire_bits_header_dst
    //output[25:0] io_rocc_imem_acquire_bits_payload_addr
    //output[2:0] io_rocc_imem_acquire_bits_payload_client_xact_id
    //output[511:0] io_rocc_imem_acquire_bits_payload_data
    //output[9:0] io_rocc_imem_acquire_bits_payload_a_type
    //output[5:0] io_rocc_imem_acquire_bits_payload_write_mask
    //output[2:0] io_rocc_imem_acquire_bits_payload_subword_addr
    //output[3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode
    output io_rocc_imem_grant_ready,
    input  io_rocc_imem_grant_valid,
    input [1:0] io_rocc_imem_grant_bits_header_src,
    input [1:0] io_rocc_imem_grant_bits_header_dst,
    input [511:0] io_rocc_imem_grant_bits_payload_data,
    input [2:0] io_rocc_imem_grant_bits_payload_client_xact_id,
    input [2:0] io_rocc_imem_grant_bits_payload_master_xact_id,
    input [4:0] io_rocc_imem_grant_bits_payload_g_type,
    input  io_rocc_imem_finish_ready,
    output io_rocc_imem_finish_valid,
    //output[1:0] io_rocc_imem_finish_bits_header_src
    //output[1:0] io_rocc_imem_finish_bits_header_dst
    //output[2:0] io_rocc_imem_finish_bits_payload_master_xact_id
    input  io_rocc_iptw_req_ready,
    output io_rocc_iptw_req_valid,
    //output[29:0] io_rocc_iptw_req_bits
    input  io_rocc_iptw_resp_valid,
    input  io_rocc_iptw_resp_bits_error,
    input [18:0] io_rocc_iptw_resp_bits_ppn,
    input [5:0] io_rocc_iptw_resp_bits_perm,
    input [7:0] io_rocc_iptw_status_ip,
    input [7:0] io_rocc_iptw_status_im,
    input [6:0] io_rocc_iptw_status_zero,
    input  io_rocc_iptw_status_er,
    input  io_rocc_iptw_status_vm,
    input  io_rocc_iptw_status_s64,
    input  io_rocc_iptw_status_u64,
    input  io_rocc_iptw_status_ef,
    input  io_rocc_iptw_status_pei,
    input  io_rocc_iptw_status_ei,
    input  io_rocc_iptw_status_ps,
    input  io_rocc_iptw_status_s,
    input  io_rocc_iptw_invalidate,
    input  io_rocc_iptw_sret,
    input  io_rocc_dptw_req_ready,
    output io_rocc_dptw_req_valid,
    //output[29:0] io_rocc_dptw_req_bits
    input  io_rocc_dptw_resp_valid,
    input  io_rocc_dptw_resp_bits_error,
    input [18:0] io_rocc_dptw_resp_bits_ppn,
    input [5:0] io_rocc_dptw_resp_bits_perm,
    input [7:0] io_rocc_dptw_status_ip,
    input [7:0] io_rocc_dptw_status_im,
    input [6:0] io_rocc_dptw_status_zero,
    input  io_rocc_dptw_status_er,
    input  io_rocc_dptw_status_vm,
    input  io_rocc_dptw_status_s64,
    input  io_rocc_dptw_status_u64,
    input  io_rocc_dptw_status_ef,
    input  io_rocc_dptw_status_pei,
    input  io_rocc_dptw_status_ei,
    input  io_rocc_dptw_status_ps,
    input  io_rocc_dptw_status_s,
    input  io_rocc_dptw_invalidate,
    input  io_rocc_dptw_sret,
    input  io_rocc_pptw_req_ready,
    output io_rocc_pptw_req_valid,
    //output[29:0] io_rocc_pptw_req_bits
    input  io_rocc_pptw_resp_valid,
    input  io_rocc_pptw_resp_bits_error,
    input [18:0] io_rocc_pptw_resp_bits_ppn,
    input [5:0] io_rocc_pptw_resp_bits_perm,
    input [7:0] io_rocc_pptw_status_ip,
    input [7:0] io_rocc_pptw_status_im,
    input [6:0] io_rocc_pptw_status_zero,
    input  io_rocc_pptw_status_er,
    input  io_rocc_pptw_status_vm,
    input  io_rocc_pptw_status_s64,
    input  io_rocc_pptw_status_u64,
    input  io_rocc_pptw_status_ef,
    input  io_rocc_pptw_status_pei,
    input  io_rocc_pptw_status_ei,
    input  io_rocc_pptw_status_ps,
    input  io_rocc_pptw_status_s,
    input  io_rocc_pptw_invalidate,
    input  io_rocc_pptw_sret,
    input  io_rocc_exception,
    output[18:0] io_cacheWriteAddr,
    output[7:0] io_cacheWriteData,
    output io_cacheWriteEn,
    output[9:0] io_addrLenAddr,
    output[18:0] io_addrLenWriteData_addr,
    output[18:0] io_addrLenWriteData_len,
    output io_addrLenWriteEn_1,
    output io_addrLenWriteEn_0,
    input [18:0] io_addrLenReadData_addr,
    input [18:0] io_addrLenReadData_len,
    output io_addrLenReadEn,
    output[9:0] io_keyLenAddr,
    output[7:0] io_keyLenData,
    output io_keyLenWrite,
    output io_lock,
    input  io_halted,
    output io_writemode,
    output io_findAvailable,
    output io_resetCounts,
    input  io_keyInfo_ready,
    output io_keyInfo_valid,
    output[18:0] io_keyInfo_bits_len,
    output[3:0] io_keyInfo_bits_tag,
    input  io_keyData_ready,
    output io_keyData_valid,
    output[7:0] io_keyData_bits,
    output io_hashSel_ready,
    input  io_hashSel_valid,
    input [3:0] io_hashSel_bits_tag,
    input [9:0] io_hashSel_bits_hash,
    input  io_hashSel_bits_found,
    input  io_copyReq_ready,
    output io_copyReq_valid,
    output[9:0] io_copyReq_bits_hash,
    output[7:0] io_copyReq_bits_len
);

  reg [63:0] len;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg [3:0] state;
  wire[3:0] T123;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg [3:0] found_state;
  wire[3:0] T124;
  wire[3:0] T37;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  reg  delayCount;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[63:0] T125;
  wire[7:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire[63:0] T126;
  wire T67;
  reg [18:0] writestart;
  wire[18:0] T141;
  wire[18:0] T142;
  wire[18:0] T143;
  reg [63:0] readstart;
  wire[63:0] T144;
  wire[63:0] T145;
  wire[63:0] T146;
  reg  action;
  wire T147;
  wire T148;
  wire T149;
  wire memCmdValid;
  wire T150;
  wire T151;
  wire[7:0] T0;
  reg [9:0] hash;
  wire[9:0] T127;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire[63:0] T128;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[63:0] T129;
  wire[9:0] T76;
  wire[63:0] T130;
  wire T77;
  wire T78;
  reg [3:0] keytag;
  wire[3:0] T79;
  wire[3:0] T80;
  wire[18:0] T131;
  wire[7:0] T81;
  wire T82;
  reg  resetCounts;
  wire T132;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg  wantmode;
  wire T87;
  wire T88;
  wire T89;
  reg  findAvailable;
  wire T90;
  wire T91;
  wire T92;
  reg  writemode;
  wire T133;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  reg [2:0] setLen;
  wire[2:0] T97;
  wire[2:0] T134;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[7:0] T105;
  wire T106;
  wire T107;
  wire[1:0] T108;
  wire T109;
  reg [18:0] addrLenData_len;
  wire[18:0] T135;
  wire[63:0] T110;
  wire[63:0] T111;
  wire[63:0] T112;
  wire[63:0] T136;
  reg [18:0] addrLenData_addr;
  wire[18:0] T137;
  wire[63:0] T113;
  wire[63:0] T114;
  wire[63:0] T115;
  wire[63:0] T138;
  wire T116;
  reg [63:0] respData;
  wire[63:0] T117;
  wire[63:0] T118;
  wire[63:0] T119;
  wire[63:0] T139;
  wire[63:0] T140;
  reg [4:0] respDest;
  wire[4:0] T120;
  wire T121;
  wire T122;
  wire memhandler_io_mem_req_valid;
  wire memhandler_io_mem_req_bits_kill;
  wire[2:0] memhandler_io_mem_req_bits_typ;
  wire memhandler_io_mem_req_bits_phys;
  wire[42:0] memhandler_io_mem_req_bits_addr;
  wire[4:0] memhandler_io_mem_req_bits_cmd;
  wire memhandler_io_keyData_valid;
  wire[7:0] memhandler_io_keyData_bits;
  wire[18:0] memhandler_io_cacheWriteAddr;
  wire[7:0] memhandler_io_cacheWriteData;
  wire memhandler_io_cacheWriteEn;
  wire memhandler_io_cmd_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    len = {2{$random}};
    state = {1{$random}};
    found_state = {1{$random}};
    delayCount = {1{$random}};
    writestart = {1{$random}};
    readstart = {2{$random}};
    action = {1{$random}};
    hash = {1{$random}};
    keytag = {1{$random}};
    resetCounts = {1{$random}};
    wantmode = {1{$random}};
    findAvailable = {1{$random}};
    writemode = {1{$random}};
    setLen = {1{$random}};
    addrLenData_len = {1{$random}};
    addrLenData_addr = {1{$random}};
    respData = {2{$random}};
    respDest = {1{$random}};
  end
`endif

  assign T1 = T67 ? T126 : T2;
  assign T2 = T66 ? 64'h0 : T3;
  assign T3 = T64 ? T125 : T4;
  assign T4 = T5 ? io_rocc_cmd_bits_rs2 : len;
  assign T5 = T7 & T6;
  assign T6 = 7'h1 == io_rocc_cmd_bits_inst_funct;
  assign T7 = T8 & io_rocc_cmd_valid;
  assign T8 = 4'h0 == state;
  assign T123 = reset ? 4'h0 : T9;
  assign T9 = T61 ? 4'h0 : T10;
  assign T10 = T59 ? 4'hb : T11;
  assign T11 = T67 ? 4'ha : T12;
  assign T12 = T51 ? 4'h9 : T13;
  assign T13 = T49 ? 4'h0 : T14;
  assign T14 = T47 ? 4'hd : T15;
  assign T15 = T45 ? 4'h7 : T16;
  assign T16 = T44 ? 4'h6 : T17;
  assign T17 = T66 ? 4'hd : T18;
  assign T18 = T42 ? 4'hd : T19;
  assign T19 = T39 ? found_state : T20;
  assign T20 = T35 ? 4'h4 : T21;
  assign T21 = T33 ? 4'h3 : T22;
  assign T22 = T31 ? 4'h0 : T23;
  assign T23 = T29 ? 4'h8 : T24;
  assign T24 = T64 ? 4'h2 : T25;
  assign T25 = T5 ? 4'h2 : T26;
  assign T26 = T27 ? 4'h1 : state;
  assign T27 = T7 & T28;
  assign T28 = 7'h0 == io_rocc_cmd_bits_inst_funct;
  assign T29 = T7 & T30;
  assign T30 = 7'h5 == io_rocc_cmd_bits_inst_funct;
  assign T31 = T32 & io_halted;
  assign T32 = 4'h1 == state;
  assign T33 = T34 & io_keyInfo_ready;
  assign T34 = 4'h2 == state;
  assign T35 = T36 & memhandler_io_cmd_ready;
  assign T36 = 4'h3 == state;
  assign T124 = reset ? 4'h0 : T37;
  assign T37 = T64 ? 4'h5 : T38;
  assign T38 = T5 ? 4'hc : found_state;
  assign T39 = T40 & io_hashSel_bits_found;
  assign T40 = T41 & io_hashSel_valid;
  assign T41 = 4'h4 == state;
  assign T42 = T40 & T43;
  assign T43 = io_hashSel_bits_found ^ 1'h1;
  assign T44 = 4'h5 == state;
  assign T45 = T46 & io_copyReq_ready;
  assign T46 = 4'h6 == state;
  assign T47 = T48 & io_copyReq_ready;
  assign T48 = 4'h7 == state;
  assign T49 = T50 & io_rocc_resp_ready;
  assign T50 = 4'hd == state;
  assign T51 = T58 & T52;
  assign T52 = delayCount == 1'h0;
  assign T53 = T56 ? T55 : T54;
  assign T54 = T29 ? 1'h1 : delayCount;
  assign T55 = delayCount - 1'h1;
  assign T56 = T58 & T57;
  assign T57 = T52 ^ 1'h1;
  assign T58 = 4'h8 == state;
  assign T59 = T60 & memhandler_io_cmd_ready;
  assign T60 = 4'ha == state;
  assign T61 = T62 & memhandler_io_cmd_ready;
  assign T62 = 4'hb == state;
  assign T125 = {56'h0, T63};
  assign T63 = io_rocc_cmd_bits_rs2[3'h7:1'h0];
  assign T64 = T7 & T65;
  assign T65 = 7'h2 == io_rocc_cmd_bits_inst_funct;
  assign T66 = 4'hc == state;
  assign T126 = {45'h0, io_addrLenReadData_len};
  assign T67 = 4'h9 == state;
  assign T141 = T67 ? io_addrLenReadData_addr : T142;
  assign T142 = T64 ? 19'h0 : T143;
  assign T143 = T5 ? 19'h0 : writestart;
  assign T144 = T29 ? io_rocc_cmd_bits_rs2 : T145;
  assign T145 = T64 ? io_rocc_cmd_bits_rs1 : T146;
  assign T146 = T5 ? io_rocc_cmd_bits_rs1 : readstart;
  assign T147 = T29 ? 1'h1 : T148;
  assign T148 = T64 ? 1'h0 : T149;
  assign T149 = T5 ? 1'h0 : action;
  assign memCmdValid = T151 | T150;
  assign T150 = state == 4'ha;
  assign T151 = state == 4'h3;
  assign io_copyReq_bits_len = T0;
  assign T0 = len[3'h7:1'h0];
  assign io_copyReq_bits_hash = hash;
  assign T127 = T68[4'h9:1'h0];
  assign T68 = T39 ? T130 : T69;
  assign T69 = T29 ? T129 : T70;
  assign T70 = T74 ? io_rocc_cmd_bits_rs1 : T71;
  assign T71 = T72 ? io_rocc_cmd_bits_rs1 : T128;
  assign T128 = {54'h0, hash};
  assign T72 = T7 & T73;
  assign T73 = 7'h3 == io_rocc_cmd_bits_inst_funct;
  assign T74 = T7 & T75;
  assign T75 = 7'h4 == io_rocc_cmd_bits_inst_funct;
  assign T129 = {54'h0, T76};
  assign T76 = io_rocc_cmd_bits_rs1[4'h9:1'h0];
  assign T130 = {54'h0, io_hashSel_bits_hash};
  assign io_copyReq_valid = T77;
  assign T77 = state == 4'h6;
  assign io_hashSel_ready = T78;
  assign T78 = state == 4'h4;
  assign io_keyData_bits = memhandler_io_keyData_bits;
  assign io_keyData_valid = memhandler_io_keyData_valid;
  assign io_keyInfo_bits_tag = keytag;
  assign T79 = T64 ? T80 : keytag;
  assign T80 = io_rocc_cmd_bits_rs2[4'hb:4'h8];
  assign io_keyInfo_bits_len = T131;
  assign T131 = {11'h0, T81};
  assign T81 = len[3'h7:1'h0];
  assign io_keyInfo_valid = T82;
  assign T82 = state == 4'h2;
  assign io_resetCounts = resetCounts;
  assign T132 = reset ? 1'h0 : T83;
  assign T83 = T85 ? 1'h1 : T84;
  assign T84 = T8 ? 1'h0 : resetCounts;
  assign T85 = T31 & T86;
  assign T86 = wantmode == 1'h0;
  assign T87 = T27 ? T88 : wantmode;
  assign T88 = T89;
  assign T89 = io_rocc_cmd_bits_inst_rs1[1'h0:1'h0];
  assign io_findAvailable = findAvailable;
  assign T90 = T64 ? 1'h1 : T91;
  assign T91 = T5 ? 1'h0 : T92;
  assign T92 = T27 ? 1'h0 : findAvailable;
  assign io_writemode = writemode;
  assign T133 = reset ? 1'h1 : T93;
  assign T93 = T31 ? wantmode : writemode;
  assign io_lock = T94;
  assign T94 = state == 4'h1;
  assign io_keyLenWrite = T95;
  assign T95 = T96;
  assign T96 = setLen[1'h0:1'h0];
  assign T134 = reset ? T97 : T98;
  assign T98 = T50 ? 3'h0 : T99;
  assign T99 = T46 ? 3'h0 : T100;
  assign T100 = T44 ? 3'h1 : T101;
  assign T101 = T66 ? 3'h7 : T102;
  assign T102 = T74 ? 3'h4 : T103;
  assign T103 = T72 ? 3'h2 : T104;
  assign T104 = T8 ? 3'h0 : setLen;
  assign io_keyLenData = T105;
  assign T105 = len[3'h7:1'h0];
  assign io_keyLenAddr = hash;
  assign io_addrLenReadEn = T106;
  assign T106 = state == 4'h8;
  assign io_addrLenWriteEn_0 = T107;
  assign T107 = T108[1'h0:1'h0];
  assign T108 = setLen[2'h2:1'h1];
  assign io_addrLenWriteEn_1 = T109;
  assign T109 = T108[1'h1:1'h1];
  assign io_addrLenWriteData_len = addrLenData_len;
  assign T135 = T110[5'h12:1'h0];
  assign T110 = T44 ? 64'h0 : T111;
  assign T111 = T66 ? 64'h0 : T112;
  assign T112 = T74 ? io_rocc_cmd_bits_rs2 : T136;
  assign T136 = {45'h0, addrLenData_len};
  assign io_addrLenWriteData_addr = addrLenData_addr;
  assign T137 = T113[5'h12:1'h0];
  assign T113 = T44 ? 64'h0 : T114;
  assign T114 = T66 ? 64'h0 : T115;
  assign T115 = T72 ? io_rocc_cmd_bits_rs2 : T138;
  assign T138 = {45'h0, addrLenData_addr};
  assign io_addrLenAddr = hash;
  assign io_cacheWriteEn = memhandler_io_cacheWriteEn;
  assign io_cacheWriteData = memhandler_io_cacheWriteData;
  assign io_cacheWriteAddr = memhandler_io_cacheWriteAddr;
  assign io_rocc_pptw_req_valid = 1'h0;
  assign io_rocc_dptw_req_valid = 1'h0;
  assign io_rocc_iptw_req_valid = 1'h0;
  assign io_rocc_imem_finish_valid = 1'h0;
  assign io_rocc_imem_grant_ready = 1'h1;
  assign io_rocc_imem_acquire_valid = 1'h0;
  assign io_rocc_interrupt = 1'h0;
  assign io_rocc_busy = T116;
  assign T116 = state != 4'h0;
  assign io_rocc_mem_req_bits_cmd = memhandler_io_mem_req_bits_cmd;
  assign io_rocc_mem_req_bits_addr = memhandler_io_mem_req_bits_addr;
  assign io_rocc_mem_req_bits_phys = memhandler_io_mem_req_bits_phys;
  assign io_rocc_mem_req_bits_typ = memhandler_io_mem_req_bits_typ;
  assign io_rocc_mem_req_bits_kill = memhandler_io_mem_req_bits_kill;
  assign io_rocc_mem_req_valid = memhandler_io_mem_req_valid;
  assign io_rocc_resp_bits_data = respData;
  assign T117 = T44 ? T140 : T118;
  assign T118 = T66 ? T139 : T119;
  assign T119 = T42 ? 64'hffffff : respData;
  assign T139 = {54'h0, hash};
  assign T140 = {54'h0, hash};
  assign io_rocc_resp_bits_rd = respDest;
  assign T120 = T7 ? io_rocc_cmd_bits_inst_rd : respDest;
  assign io_rocc_resp_valid = T121;
  assign T121 = state == 4'hd;
  assign io_rocc_cmd_ready = T122;
  assign T122 = state == 4'h0;
  MemoryHandler memhandler(.clk(clk), .reset(reset),
       .io_mem_req_ready( io_rocc_mem_req_ready ),
       .io_mem_req_valid( memhandler_io_mem_req_valid ),
       .io_mem_req_bits_kill( memhandler_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( memhandler_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( memhandler_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( memhandler_io_mem_req_bits_addr ),
       //.io_mem_req_bits_data(  )
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( memhandler_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( io_rocc_mem_resp_valid ),
       .io_mem_resp_bits_nack( io_rocc_mem_resp_bits_nack ),
       .io_mem_resp_bits_replay( io_rocc_mem_resp_bits_replay ),
       .io_mem_resp_bits_typ( io_rocc_mem_resp_bits_typ ),
       .io_mem_resp_bits_has_data( io_rocc_mem_resp_bits_has_data ),
       .io_mem_resp_bits_data( io_rocc_mem_resp_bits_data ),
       .io_mem_resp_bits_data_subword( io_rocc_mem_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( io_rocc_mem_resp_bits_tag ),
       .io_mem_resp_bits_cmd( io_rocc_mem_resp_bits_cmd ),
       .io_mem_resp_bits_addr( io_rocc_mem_resp_bits_addr ),
       .io_mem_resp_bits_store_data( io_rocc_mem_resp_bits_store_data ),
       .io_mem_replay_next_valid( io_rocc_mem_replay_next_valid ),
       .io_mem_replay_next_bits( io_rocc_mem_replay_next_bits ),
       .io_mem_xcpt_ma_ld( io_rocc_mem_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( io_rocc_mem_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( io_rocc_mem_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( io_rocc_mem_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( io_rocc_mem_ptw_req_valid ),
       .io_mem_ptw_req_bits( io_rocc_mem_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( io_rocc_mem_ordered ),
       .io_keyData_ready( io_keyData_ready ),
       .io_keyData_valid( memhandler_io_keyData_valid ),
       .io_keyData_bits( memhandler_io_keyData_bits ),
       .io_cacheWriteAddr( memhandler_io_cacheWriteAddr ),
       .io_cacheWriteData( memhandler_io_cacheWriteData ),
       .io_cacheWriteEn( memhandler_io_cacheWriteEn ),
       .io_cmd_ready( memhandler_io_cmd_ready ),
       .io_cmd_valid( memCmdValid ),
       .io_cmd_bits_action( action ),
       .io_cmd_bits_readstart( readstart ),
       .io_cmd_bits_writestart( writestart ),
       .io_cmd_bits_len( len )
  );

  always @(posedge clk) begin
    if(T67) begin
      len <= T126;
    end else if(T66) begin
      len <= 64'h0;
    end else if(T64) begin
      len <= T125;
    end else if(T5) begin
      len <= io_rocc_cmd_bits_rs2;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T61) begin
      state <= 4'h0;
    end else if(T59) begin
      state <= 4'hb;
    end else if(T67) begin
      state <= 4'ha;
    end else if(T51) begin
      state <= 4'h9;
    end else if(T49) begin
      state <= 4'h0;
    end else if(T47) begin
      state <= 4'hd;
    end else if(T45) begin
      state <= 4'h7;
    end else if(T44) begin
      state <= 4'h6;
    end else if(T66) begin
      state <= 4'hd;
    end else if(T42) begin
      state <= 4'hd;
    end else if(T39) begin
      state <= found_state;
    end else if(T35) begin
      state <= 4'h4;
    end else if(T33) begin
      state <= 4'h3;
    end else if(T31) begin
      state <= 4'h0;
    end else if(T29) begin
      state <= 4'h8;
    end else if(T64) begin
      state <= 4'h2;
    end else if(T5) begin
      state <= 4'h2;
    end else if(T27) begin
      state <= 4'h1;
    end
    if(reset) begin
      found_state <= 4'h0;
    end else if(T64) begin
      found_state <= 4'h5;
    end else if(T5) begin
      found_state <= 4'hc;
    end
    if(T56) begin
      delayCount <= T55;
    end else if(T29) begin
      delayCount <= 1'h1;
    end
    if(T67) begin
      writestart <= io_addrLenReadData_addr;
    end else if(T64) begin
      writestart <= 19'h0;
    end else if(T5) begin
      writestart <= 19'h0;
    end
    if(T29) begin
      readstart <= io_rocc_cmd_bits_rs2;
    end else if(T64) begin
      readstart <= io_rocc_cmd_bits_rs1;
    end else if(T5) begin
      readstart <= io_rocc_cmd_bits_rs1;
    end
    if(T29) begin
      action <= 1'h1;
    end else if(T64) begin
      action <= 1'h0;
    end else if(T5) begin
      action <= 1'h0;
    end
    hash <= T127;
    if(T64) begin
      keytag <= T80;
    end
    if(reset) begin
      resetCounts <= 1'h0;
    end else if(T85) begin
      resetCounts <= 1'h1;
    end else if(T8) begin
      resetCounts <= 1'h0;
    end
    if(T27) begin
      wantmode <= T88;
    end
    if(T64) begin
      findAvailable <= 1'h1;
    end else if(T5) begin
      findAvailable <= 1'h0;
    end else if(T27) begin
      findAvailable <= 1'h0;
    end
    if(reset) begin
      writemode <= 1'h1;
    end else if(T31) begin
      writemode <= wantmode;
    end
    if(reset) begin
      setLen <= T97;
    end else if(T50) begin
      setLen <= 3'h0;
    end else if(T46) begin
      setLen <= 3'h0;
    end else if(T44) begin
      setLen <= 3'h1;
    end else if(T66) begin
      setLen <= 3'h7;
    end else if(T74) begin
      setLen <= 3'h4;
    end else if(T72) begin
      setLen <= 3'h2;
    end else if(T8) begin
      setLen <= 3'h0;
    end
    addrLenData_len <= T135;
    addrLenData_addr <= T137;
    if(T44) begin
      respData <= T140;
    end else if(T66) begin
      respData <= T139;
    end else if(T42) begin
      respData <= 64'hffffff;
    end
    if(T7) begin
      respDest <= io_rocc_cmd_bits_inst_rd;
    end
  end
endmodule

module KeyValueStore(input clk, input reset,
    output io_keyInfo_ready,
    input  io_keyInfo_valid,
    input [7:0] io_keyInfo_bits_len,
    input [3:0] io_keyInfo_bits_tag,
    output io_keyData_ready,
    input  io_keyData_valid,
    input [7:0] io_keyData_bits,
    input  io_resultInfo_ready,
    output io_resultInfo_valid,
    output[18:0] io_resultInfo_bits_len,
    output[3:0] io_resultInfo_bits_tag,
    input  io_resultData_ready,
    output io_resultData_valid,
    output[7:0] io_resultData_bits,
    output io_writeready,
    output io_readready,
    output io_rocc_cmd_ready,
    input  io_rocc_cmd_valid,
    input [6:0] io_rocc_cmd_bits_inst_funct,
    input [4:0] io_rocc_cmd_bits_inst_rs2,
    input [4:0] io_rocc_cmd_bits_inst_rs1,
    input  io_rocc_cmd_bits_inst_xd,
    input  io_rocc_cmd_bits_inst_xs1,
    input  io_rocc_cmd_bits_inst_xs2,
    input [4:0] io_rocc_cmd_bits_inst_rd,
    input [6:0] io_rocc_cmd_bits_inst_opcode,
    input [63:0] io_rocc_cmd_bits_rs1,
    input [63:0] io_rocc_cmd_bits_rs2,
    input  io_rocc_resp_ready,
    output io_rocc_resp_valid,
    output[4:0] io_rocc_resp_bits_rd,
    output[63:0] io_rocc_resp_bits_data,
    input  io_rocc_mem_req_ready,
    output io_rocc_mem_req_valid,
    output io_rocc_mem_req_bits_kill,
    output[2:0] io_rocc_mem_req_bits_typ,
    output io_rocc_mem_req_bits_phys,
    output[42:0] io_rocc_mem_req_bits_addr,
    //output[63:0] io_rocc_mem_req_bits_data
    //output[8:0] io_rocc_mem_req_bits_tag
    output[4:0] io_rocc_mem_req_bits_cmd,
    input  io_rocc_mem_resp_valid,
    input  io_rocc_mem_resp_bits_nack,
    input  io_rocc_mem_resp_bits_replay,
    input [2:0] io_rocc_mem_resp_bits_typ,
    input  io_rocc_mem_resp_bits_has_data,
    input [63:0] io_rocc_mem_resp_bits_data,
    input [63:0] io_rocc_mem_resp_bits_data_subword,
    input [8:0] io_rocc_mem_resp_bits_tag,
    input [3:0] io_rocc_mem_resp_bits_cmd,
    input [42:0] io_rocc_mem_resp_bits_addr,
    input [63:0] io_rocc_mem_resp_bits_store_data,
    input  io_rocc_mem_replay_next_valid,
    input [8:0] io_rocc_mem_replay_next_bits,
    input  io_rocc_mem_xcpt_ma_ld,
    input  io_rocc_mem_xcpt_ma_st,
    input  io_rocc_mem_xcpt_pf_ld,
    input  io_rocc_mem_xcpt_pf_st,
    //output io_rocc_mem_ptw_req_ready
    input  io_rocc_mem_ptw_req_valid,
    input [29:0] io_rocc_mem_ptw_req_bits,
    //output io_rocc_mem_ptw_resp_valid
    //output io_rocc_mem_ptw_resp_bits_error
    //output[18:0] io_rocc_mem_ptw_resp_bits_ppn
    //output[5:0] io_rocc_mem_ptw_resp_bits_perm
    //output[7:0] io_rocc_mem_ptw_status_ip
    //output[7:0] io_rocc_mem_ptw_status_im
    //output[6:0] io_rocc_mem_ptw_status_zero
    //output io_rocc_mem_ptw_status_er
    //output io_rocc_mem_ptw_status_vm
    //output io_rocc_mem_ptw_status_s64
    //output io_rocc_mem_ptw_status_u64
    //output io_rocc_mem_ptw_status_ef
    //output io_rocc_mem_ptw_status_pei
    //output io_rocc_mem_ptw_status_ei
    //output io_rocc_mem_ptw_status_ps
    //output io_rocc_mem_ptw_status_s
    //output io_rocc_mem_ptw_invalidate
    //output io_rocc_mem_ptw_sret
    input  io_rocc_mem_ordered,
    output io_rocc_busy,
    input  io_rocc_s,
    output io_rocc_interrupt,
    input  io_rocc_imem_acquire_ready,
    output io_rocc_imem_acquire_valid,
    //output[1:0] io_rocc_imem_acquire_bits_header_src
    //output[1:0] io_rocc_imem_acquire_bits_header_dst
    //output[25:0] io_rocc_imem_acquire_bits_payload_addr
    //output[2:0] io_rocc_imem_acquire_bits_payload_client_xact_id
    //output[511:0] io_rocc_imem_acquire_bits_payload_data
    //output[9:0] io_rocc_imem_acquire_bits_payload_a_type
    //output[5:0] io_rocc_imem_acquire_bits_payload_write_mask
    //output[2:0] io_rocc_imem_acquire_bits_payload_subword_addr
    //output[3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode
    output io_rocc_imem_grant_ready,
    input  io_rocc_imem_grant_valid,
    input [1:0] io_rocc_imem_grant_bits_header_src,
    input [1:0] io_rocc_imem_grant_bits_header_dst,
    input [511:0] io_rocc_imem_grant_bits_payload_data,
    input [2:0] io_rocc_imem_grant_bits_payload_client_xact_id,
    input [2:0] io_rocc_imem_grant_bits_payload_master_xact_id,
    input [4:0] io_rocc_imem_grant_bits_payload_g_type,
    input  io_rocc_imem_finish_ready,
    output io_rocc_imem_finish_valid,
    //output[1:0] io_rocc_imem_finish_bits_header_src
    //output[1:0] io_rocc_imem_finish_bits_header_dst
    //output[2:0] io_rocc_imem_finish_bits_payload_master_xact_id
    input  io_rocc_iptw_req_ready,
    output io_rocc_iptw_req_valid,
    //output[29:0] io_rocc_iptw_req_bits
    input  io_rocc_iptw_resp_valid,
    input  io_rocc_iptw_resp_bits_error,
    input [18:0] io_rocc_iptw_resp_bits_ppn,
    input [5:0] io_rocc_iptw_resp_bits_perm,
    input [7:0] io_rocc_iptw_status_ip,
    input [7:0] io_rocc_iptw_status_im,
    input [6:0] io_rocc_iptw_status_zero,
    input  io_rocc_iptw_status_er,
    input  io_rocc_iptw_status_vm,
    input  io_rocc_iptw_status_s64,
    input  io_rocc_iptw_status_u64,
    input  io_rocc_iptw_status_ef,
    input  io_rocc_iptw_status_pei,
    input  io_rocc_iptw_status_ei,
    input  io_rocc_iptw_status_ps,
    input  io_rocc_iptw_status_s,
    input  io_rocc_iptw_invalidate,
    input  io_rocc_iptw_sret,
    input  io_rocc_dptw_req_ready,
    output io_rocc_dptw_req_valid,
    //output[29:0] io_rocc_dptw_req_bits
    input  io_rocc_dptw_resp_valid,
    input  io_rocc_dptw_resp_bits_error,
    input [18:0] io_rocc_dptw_resp_bits_ppn,
    input [5:0] io_rocc_dptw_resp_bits_perm,
    input [7:0] io_rocc_dptw_status_ip,
    input [7:0] io_rocc_dptw_status_im,
    input [6:0] io_rocc_dptw_status_zero,
    input  io_rocc_dptw_status_er,
    input  io_rocc_dptw_status_vm,
    input  io_rocc_dptw_status_s64,
    input  io_rocc_dptw_status_u64,
    input  io_rocc_dptw_status_ef,
    input  io_rocc_dptw_status_pei,
    input  io_rocc_dptw_status_ei,
    input  io_rocc_dptw_status_ps,
    input  io_rocc_dptw_status_s,
    input  io_rocc_dptw_invalidate,
    input  io_rocc_dptw_sret,
    input  io_rocc_pptw_req_ready,
    output io_rocc_pptw_req_valid,
    //output[29:0] io_rocc_pptw_req_bits
    input  io_rocc_pptw_resp_valid,
    input  io_rocc_pptw_resp_bits_error,
    input [18:0] io_rocc_pptw_resp_bits_ppn,
    input [5:0] io_rocc_pptw_resp_bits_perm,
    input [7:0] io_rocc_pptw_status_ip,
    input [7:0] io_rocc_pptw_status_im,
    input [6:0] io_rocc_pptw_status_zero,
    input  io_rocc_pptw_status_er,
    input  io_rocc_pptw_status_vm,
    input  io_rocc_pptw_status_s64,
    input  io_rocc_pptw_status_u64,
    input  io_rocc_pptw_status_ef,
    input  io_rocc_pptw_status_pei,
    input  io_rocc_pptw_status_ei,
    input  io_rocc_pptw_status_ps,
    input  io_rocc_pptw_status_s,
    input  io_rocc_pptw_invalidate,
    input  io_rocc_pptw_sret,
    input  io_rocc_exception
);

  wire[7:0] T5;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire Queue_14_io_enq_ready;
  wire Queue_14_io_deq_valid;
  wire[7:0] Queue_14_io_deq_bits_len;
  wire[3:0] Queue_14_io_deq_bits_tag;
  wire Queue_15_io_enq_ready;
  wire Queue_15_io_deq_valid;
  wire[7:0] Queue_15_io_deq_bits;
  wire Queue_16_io_enq_ready;
  wire Queue_16_io_deq_valid;
  wire[18:0] Queue_16_io_deq_bits_len;
  wire[3:0] Queue_16_io_deq_bits_tag;
  wire Queue_17_io_enq_ready;
  wire Queue_17_io_deq_valid;
  wire[7:0] Queue_17_io_deq_bits;
  wire ctrl_io_rocc_cmd_ready;
  wire ctrl_io_rocc_resp_valid;
  wire[4:0] ctrl_io_rocc_resp_bits_rd;
  wire[63:0] ctrl_io_rocc_resp_bits_data;
  wire ctrl_io_rocc_mem_req_valid;
  wire ctrl_io_rocc_mem_req_bits_kill;
  wire[2:0] ctrl_io_rocc_mem_req_bits_typ;
  wire ctrl_io_rocc_mem_req_bits_phys;
  wire[42:0] ctrl_io_rocc_mem_req_bits_addr;
  wire[4:0] ctrl_io_rocc_mem_req_bits_cmd;
  wire ctrl_io_rocc_busy;
  wire ctrl_io_rocc_interrupt;
  wire ctrl_io_rocc_imem_acquire_valid;
  wire ctrl_io_rocc_imem_grant_ready;
  wire ctrl_io_rocc_imem_finish_valid;
  wire ctrl_io_rocc_iptw_req_valid;
  wire ctrl_io_rocc_dptw_req_valid;
  wire ctrl_io_rocc_pptw_req_valid;
  wire[18:0] ctrl_io_cacheWriteAddr;
  wire[7:0] ctrl_io_cacheWriteData;
  wire ctrl_io_cacheWriteEn;
  wire[9:0] ctrl_io_addrLenAddr;
  wire[18:0] ctrl_io_addrLenWriteData_addr;
  wire[18:0] ctrl_io_addrLenWriteData_len;
  wire ctrl_io_addrLenWriteEn_1;
  wire ctrl_io_addrLenWriteEn_0;
  wire ctrl_io_addrLenReadEn;
  wire[9:0] ctrl_io_keyLenAddr;
  wire[7:0] ctrl_io_keyLenData;
  wire ctrl_io_keyLenWrite;
  wire ctrl_io_lock;
  wire ctrl_io_writemode;
  wire ctrl_io_findAvailable;
  wire ctrl_io_resetCounts;
  wire ctrl_io_keyInfo_valid;
  wire[18:0] ctrl_io_keyInfo_bits_len;
  wire[3:0] ctrl_io_keyInfo_bits_tag;
  wire ctrl_io_keyData_valid;
  wire[7:0] ctrl_io_keyData_bits;
  wire ctrl_io_hashSel_ready;
  wire ctrl_io_copyReq_valid;
  wire[9:0] ctrl_io_copyReq_bits_hash;
  wire[7:0] ctrl_io_copyReq_bits_len;
  wire lookup_io_halted;
  wire lookup_io_readKeyInfo_ready;
  wire lookup_io_readKeyData_ready;
  wire lookup_io_writeKeyInfo_ready;
  wire lookup_io_writeKeyData_ready;
  wire lookup_io_hashSel_valid;
  wire[3:0] lookup_io_hashSel_bits_tag;
  wire[9:0] lookup_io_hashSel_bits_hash;
  wire lookup_io_hashSel_bits_found;
  wire lookup_io_copyReq_ready;
  wire lookup_io_resultInfo_valid;
  wire[18:0] lookup_io_resultInfo_bits_len;
  wire[3:0] lookup_io_resultInfo_bits_tag;
  wire lookup_io_resultData_valid;
  wire[7:0] lookup_io_resultData_bits;
  wire[18:0] lookup_io_addrLenReadData_addr;
  wire[18:0] lookup_io_addrLenReadData_len;


  assign T5 = ctrl_io_keyInfo_bits_len[3'h7:1'h0];
  assign io_rocc_pptw_req_valid = ctrl_io_rocc_pptw_req_valid;
  assign io_rocc_dptw_req_valid = ctrl_io_rocc_dptw_req_valid;
  assign io_rocc_iptw_req_valid = ctrl_io_rocc_iptw_req_valid;
  assign io_rocc_imem_finish_valid = ctrl_io_rocc_imem_finish_valid;
  assign io_rocc_imem_grant_ready = ctrl_io_rocc_imem_grant_ready;
  assign io_rocc_imem_acquire_valid = ctrl_io_rocc_imem_acquire_valid;
  assign io_rocc_interrupt = ctrl_io_rocc_interrupt;
  assign io_rocc_busy = ctrl_io_rocc_busy;
  assign io_rocc_mem_req_bits_cmd = ctrl_io_rocc_mem_req_bits_cmd;
  assign io_rocc_mem_req_bits_addr = ctrl_io_rocc_mem_req_bits_addr;
  assign io_rocc_mem_req_bits_phys = ctrl_io_rocc_mem_req_bits_phys;
  assign io_rocc_mem_req_bits_typ = ctrl_io_rocc_mem_req_bits_typ;
  assign io_rocc_mem_req_bits_kill = ctrl_io_rocc_mem_req_bits_kill;
  assign io_rocc_mem_req_valid = ctrl_io_rocc_mem_req_valid;
  assign io_rocc_resp_bits_data = ctrl_io_rocc_resp_bits_data;
  assign io_rocc_resp_bits_rd = ctrl_io_rocc_resp_bits_rd;
  assign io_rocc_resp_valid = ctrl_io_rocc_resp_valid;
  assign io_rocc_cmd_ready = ctrl_io_rocc_cmd_ready;
  assign io_readready = T0;
  assign T0 = T2 & T1;
  assign T1 = lookup_io_halted ^ 1'h1;
  assign T2 = ctrl_io_writemode ^ 1'h1;
  assign io_writeready = T3;
  assign T3 = ctrl_io_writemode & T4;
  assign T4 = lookup_io_halted ^ 1'h1;
  assign io_resultData_bits = Queue_17_io_deq_bits;
  assign io_resultData_valid = Queue_17_io_deq_valid;
  assign io_resultInfo_bits_tag = Queue_16_io_deq_bits_tag;
  assign io_resultInfo_bits_len = Queue_16_io_deq_bits_len;
  assign io_resultInfo_valid = Queue_16_io_deq_valid;
  assign io_keyData_ready = Queue_15_io_enq_ready;
  assign io_keyInfo_ready = Queue_14_io_enq_ready;
  LookupPipeline lookup(.clk(clk), .reset(reset),
       .io_lock( ctrl_io_lock ),
       .io_halted( lookup_io_halted ),
       .io_writemode( ctrl_io_writemode ),
       .io_findAvailable( ctrl_io_findAvailable ),
       .io_resetCounts( ctrl_io_resetCounts ),
       .io_readKeyInfo_ready( lookup_io_readKeyInfo_ready ),
       .io_readKeyInfo_valid( Queue_14_io_deq_valid ),
       .io_readKeyInfo_bits_len( Queue_14_io_deq_bits_len ),
       .io_readKeyInfo_bits_tag( Queue_14_io_deq_bits_tag ),
       .io_readKeyData_ready( lookup_io_readKeyData_ready ),
       .io_readKeyData_valid( Queue_15_io_deq_valid ),
       .io_readKeyData_bits( Queue_15_io_deq_bits ),
       .io_writeKeyInfo_ready( lookup_io_writeKeyInfo_ready ),
       .io_writeKeyInfo_valid( ctrl_io_keyInfo_valid ),
       .io_writeKeyInfo_bits_len( T5 ),
       .io_writeKeyInfo_bits_tag( ctrl_io_keyInfo_bits_tag ),
       .io_writeKeyData_ready( lookup_io_writeKeyData_ready ),
       .io_writeKeyData_valid( ctrl_io_keyData_valid ),
       .io_writeKeyData_bits( ctrl_io_keyData_bits ),
       .io_hashSel_ready( ctrl_io_hashSel_ready ),
       .io_hashSel_valid( lookup_io_hashSel_valid ),
       .io_hashSel_bits_tag( lookup_io_hashSel_bits_tag ),
       .io_hashSel_bits_hash( lookup_io_hashSel_bits_hash ),
       .io_hashSel_bits_found( lookup_io_hashSel_bits_found ),
       .io_copyReq_ready( lookup_io_copyReq_ready ),
       .io_copyReq_valid( ctrl_io_copyReq_valid ),
       .io_copyReq_bits_hash( ctrl_io_copyReq_bits_hash ),
       .io_copyReq_bits_len( ctrl_io_copyReq_bits_len ),
       .io_resultInfo_ready( Queue_16_io_enq_ready ),
       .io_resultInfo_valid( lookup_io_resultInfo_valid ),
       .io_resultInfo_bits_len( lookup_io_resultInfo_bits_len ),
       .io_resultInfo_bits_tag( lookup_io_resultInfo_bits_tag ),
       .io_resultData_ready( Queue_17_io_enq_ready ),
       .io_resultData_valid( lookup_io_resultData_valid ),
       .io_resultData_bits( lookup_io_resultData_bits ),
       .io_cacheWriteAddr( ctrl_io_cacheWriteAddr ),
       .io_cacheWriteData( ctrl_io_cacheWriteData ),
       .io_cacheWriteEn( ctrl_io_cacheWriteEn ),
       .io_addrLenAddr( ctrl_io_addrLenAddr ),
       .io_addrLenWriteData_addr( ctrl_io_addrLenWriteData_addr ),
       .io_addrLenWriteData_len( ctrl_io_addrLenWriteData_len ),
       .io_addrLenWriteEn_1( ctrl_io_addrLenWriteEn_1 ),
       .io_addrLenWriteEn_0( ctrl_io_addrLenWriteEn_0 ),
       .io_addrLenReadData_addr( lookup_io_addrLenReadData_addr ),
       .io_addrLenReadData_len( lookup_io_addrLenReadData_len ),
       .io_addrLenReadEn( ctrl_io_addrLenReadEn ),
       .io_keyLenAddr( ctrl_io_keyLenAddr ),
       .io_keyLenData( ctrl_io_keyLenData ),
       .io_keyLenWrite( ctrl_io_keyLenWrite )
  );
  Queue_8 Queue_14(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_14_io_enq_ready ),
       .io_enq_valid( io_keyInfo_valid ),
       .io_enq_bits_len( io_keyInfo_bits_len ),
       .io_enq_bits_tag( io_keyInfo_bits_tag ),
       .io_deq_ready( lookup_io_readKeyInfo_ready ),
       .io_deq_valid( Queue_14_io_deq_valid ),
       .io_deq_bits_len( Queue_14_io_deq_bits_len ),
       .io_deq_bits_tag( Queue_14_io_deq_bits_tag )
  );
  Queue_9 Queue_15(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_15_io_enq_ready ),
       .io_enq_valid( io_keyData_valid ),
       .io_enq_bits( io_keyData_bits ),
       .io_deq_ready( lookup_io_readKeyData_ready ),
       .io_deq_valid( Queue_15_io_deq_valid ),
       .io_deq_bits( Queue_15_io_deq_bits )
  );
  Queue_10 Queue_16(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_16_io_enq_ready ),
       .io_enq_valid( lookup_io_resultInfo_valid ),
       .io_enq_bits_len( lookup_io_resultInfo_bits_len ),
       .io_enq_bits_tag( lookup_io_resultInfo_bits_tag ),
       .io_deq_ready( io_resultInfo_ready ),
       .io_deq_valid( Queue_16_io_deq_valid ),
       .io_deq_bits_len( Queue_16_io_deq_bits_len ),
       .io_deq_bits_tag( Queue_16_io_deq_bits_tag )
  );
  Queue_9 Queue_17(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_17_io_enq_ready ),
       .io_enq_valid( lookup_io_resultData_valid ),
       .io_enq_bits( lookup_io_resultData_bits ),
       .io_deq_ready( io_resultData_ready ),
       .io_deq_valid( Queue_17_io_deq_valid ),
       .io_deq_bits( Queue_17_io_deq_bits )
  );
  CtrlModule ctrl(.clk(clk), .reset(reset),
       .io_rocc_cmd_ready( ctrl_io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( io_rocc_cmd_valid ),
       .io_rocc_cmd_bits_inst_funct( io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( io_rocc_cmd_bits_rs2 ),
       .io_rocc_resp_ready( io_rocc_resp_ready ),
       .io_rocc_resp_valid( ctrl_io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( ctrl_io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( ctrl_io_rocc_resp_bits_data ),
       .io_rocc_mem_req_ready( io_rocc_mem_req_ready ),
       .io_rocc_mem_req_valid( ctrl_io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( ctrl_io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( ctrl_io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( ctrl_io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( ctrl_io_rocc_mem_req_bits_addr ),
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_req_bits_tag(  )
       .io_rocc_mem_req_bits_cmd( ctrl_io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_resp_valid( io_rocc_mem_resp_valid ),
       .io_rocc_mem_resp_bits_nack( io_rocc_mem_resp_bits_nack ),
       .io_rocc_mem_resp_bits_replay( io_rocc_mem_resp_bits_replay ),
       .io_rocc_mem_resp_bits_typ( io_rocc_mem_resp_bits_typ ),
       .io_rocc_mem_resp_bits_has_data( io_rocc_mem_resp_bits_has_data ),
       .io_rocc_mem_resp_bits_data( io_rocc_mem_resp_bits_data ),
       .io_rocc_mem_resp_bits_data_subword( io_rocc_mem_resp_bits_data_subword ),
       .io_rocc_mem_resp_bits_tag( io_rocc_mem_resp_bits_tag ),
       .io_rocc_mem_resp_bits_cmd( io_rocc_mem_resp_bits_cmd ),
       .io_rocc_mem_resp_bits_addr( io_rocc_mem_resp_bits_addr ),
       .io_rocc_mem_resp_bits_store_data( io_rocc_mem_resp_bits_store_data ),
       .io_rocc_mem_replay_next_valid( io_rocc_mem_replay_next_valid ),
       .io_rocc_mem_replay_next_bits( io_rocc_mem_replay_next_bits ),
       .io_rocc_mem_xcpt_ma_ld( io_rocc_mem_xcpt_ma_ld ),
       .io_rocc_mem_xcpt_ma_st( io_rocc_mem_xcpt_ma_st ),
       .io_rocc_mem_xcpt_pf_ld( io_rocc_mem_xcpt_pf_ld ),
       .io_rocc_mem_xcpt_pf_st( io_rocc_mem_xcpt_pf_st ),
       //.io_rocc_mem_ptw_req_ready(  )
       .io_rocc_mem_ptw_req_valid( io_rocc_mem_ptw_req_valid ),
       .io_rocc_mem_ptw_req_bits( io_rocc_mem_ptw_req_bits ),
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       .io_rocc_mem_ordered( io_rocc_mem_ordered ),
       .io_rocc_busy( ctrl_io_rocc_busy ),
       .io_rocc_s( io_rocc_s ),
       .io_rocc_interrupt( ctrl_io_rocc_interrupt ),
       .io_rocc_imem_acquire_ready( io_rocc_imem_acquire_ready ),
       .io_rocc_imem_acquire_valid( ctrl_io_rocc_imem_acquire_valid ),
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_write_mask(  )
       //.io_rocc_imem_acquire_bits_payload_subword_addr(  )
       //.io_rocc_imem_acquire_bits_payload_atomic_opcode(  )
       .io_rocc_imem_grant_ready( ctrl_io_rocc_imem_grant_ready ),
       .io_rocc_imem_grant_valid( io_rocc_imem_grant_valid ),
       .io_rocc_imem_grant_bits_header_src( io_rocc_imem_grant_bits_header_src ),
       .io_rocc_imem_grant_bits_header_dst( io_rocc_imem_grant_bits_header_dst ),
       .io_rocc_imem_grant_bits_payload_data( io_rocc_imem_grant_bits_payload_data ),
       .io_rocc_imem_grant_bits_payload_client_xact_id( io_rocc_imem_grant_bits_payload_client_xact_id ),
       .io_rocc_imem_grant_bits_payload_master_xact_id( io_rocc_imem_grant_bits_payload_master_xact_id ),
       .io_rocc_imem_grant_bits_payload_g_type( io_rocc_imem_grant_bits_payload_g_type ),
       .io_rocc_imem_finish_ready( io_rocc_imem_finish_ready ),
       .io_rocc_imem_finish_valid( ctrl_io_rocc_imem_finish_valid ),
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       .io_rocc_iptw_req_ready( io_rocc_iptw_req_ready ),
       .io_rocc_iptw_req_valid( ctrl_io_rocc_iptw_req_valid ),
       //.io_rocc_iptw_req_bits(  )
       .io_rocc_iptw_resp_valid( io_rocc_iptw_resp_valid ),
       .io_rocc_iptw_resp_bits_error( io_rocc_iptw_resp_bits_error ),
       .io_rocc_iptw_resp_bits_ppn( io_rocc_iptw_resp_bits_ppn ),
       .io_rocc_iptw_resp_bits_perm( io_rocc_iptw_resp_bits_perm ),
       .io_rocc_iptw_status_ip( io_rocc_iptw_status_ip ),
       .io_rocc_iptw_status_im( io_rocc_iptw_status_im ),
       .io_rocc_iptw_status_zero( io_rocc_iptw_status_zero ),
       .io_rocc_iptw_status_er( io_rocc_iptw_status_er ),
       .io_rocc_iptw_status_vm( io_rocc_iptw_status_vm ),
       .io_rocc_iptw_status_s64( io_rocc_iptw_status_s64 ),
       .io_rocc_iptw_status_u64( io_rocc_iptw_status_u64 ),
       .io_rocc_iptw_status_ef( io_rocc_iptw_status_ef ),
       .io_rocc_iptw_status_pei( io_rocc_iptw_status_pei ),
       .io_rocc_iptw_status_ei( io_rocc_iptw_status_ei ),
       .io_rocc_iptw_status_ps( io_rocc_iptw_status_ps ),
       .io_rocc_iptw_status_s( io_rocc_iptw_status_s ),
       .io_rocc_iptw_invalidate( io_rocc_iptw_invalidate ),
       .io_rocc_iptw_sret( io_rocc_iptw_sret ),
       .io_rocc_dptw_req_ready( io_rocc_dptw_req_ready ),
       .io_rocc_dptw_req_valid( ctrl_io_rocc_dptw_req_valid ),
       //.io_rocc_dptw_req_bits(  )
       .io_rocc_dptw_resp_valid( io_rocc_dptw_resp_valid ),
       .io_rocc_dptw_resp_bits_error( io_rocc_dptw_resp_bits_error ),
       .io_rocc_dptw_resp_bits_ppn( io_rocc_dptw_resp_bits_ppn ),
       .io_rocc_dptw_resp_bits_perm( io_rocc_dptw_resp_bits_perm ),
       .io_rocc_dptw_status_ip( io_rocc_dptw_status_ip ),
       .io_rocc_dptw_status_im( io_rocc_dptw_status_im ),
       .io_rocc_dptw_status_zero( io_rocc_dptw_status_zero ),
       .io_rocc_dptw_status_er( io_rocc_dptw_status_er ),
       .io_rocc_dptw_status_vm( io_rocc_dptw_status_vm ),
       .io_rocc_dptw_status_s64( io_rocc_dptw_status_s64 ),
       .io_rocc_dptw_status_u64( io_rocc_dptw_status_u64 ),
       .io_rocc_dptw_status_ef( io_rocc_dptw_status_ef ),
       .io_rocc_dptw_status_pei( io_rocc_dptw_status_pei ),
       .io_rocc_dptw_status_ei( io_rocc_dptw_status_ei ),
       .io_rocc_dptw_status_ps( io_rocc_dptw_status_ps ),
       .io_rocc_dptw_status_s( io_rocc_dptw_status_s ),
       .io_rocc_dptw_invalidate( io_rocc_dptw_invalidate ),
       .io_rocc_dptw_sret( io_rocc_dptw_sret ),
       .io_rocc_pptw_req_ready( io_rocc_pptw_req_ready ),
       .io_rocc_pptw_req_valid( ctrl_io_rocc_pptw_req_valid ),
       //.io_rocc_pptw_req_bits(  )
       .io_rocc_pptw_resp_valid( io_rocc_pptw_resp_valid ),
       .io_rocc_pptw_resp_bits_error( io_rocc_pptw_resp_bits_error ),
       .io_rocc_pptw_resp_bits_ppn( io_rocc_pptw_resp_bits_ppn ),
       .io_rocc_pptw_resp_bits_perm( io_rocc_pptw_resp_bits_perm ),
       .io_rocc_pptw_status_ip( io_rocc_pptw_status_ip ),
       .io_rocc_pptw_status_im( io_rocc_pptw_status_im ),
       .io_rocc_pptw_status_zero( io_rocc_pptw_status_zero ),
       .io_rocc_pptw_status_er( io_rocc_pptw_status_er ),
       .io_rocc_pptw_status_vm( io_rocc_pptw_status_vm ),
       .io_rocc_pptw_status_s64( io_rocc_pptw_status_s64 ),
       .io_rocc_pptw_status_u64( io_rocc_pptw_status_u64 ),
       .io_rocc_pptw_status_ef( io_rocc_pptw_status_ef ),
       .io_rocc_pptw_status_pei( io_rocc_pptw_status_pei ),
       .io_rocc_pptw_status_ei( io_rocc_pptw_status_ei ),
       .io_rocc_pptw_status_ps( io_rocc_pptw_status_ps ),
       .io_rocc_pptw_status_s( io_rocc_pptw_status_s ),
       .io_rocc_pptw_invalidate( io_rocc_pptw_invalidate ),
       .io_rocc_pptw_sret( io_rocc_pptw_sret ),
       .io_rocc_exception( io_rocc_exception ),
       .io_cacheWriteAddr( ctrl_io_cacheWriteAddr ),
       .io_cacheWriteData( ctrl_io_cacheWriteData ),
       .io_cacheWriteEn( ctrl_io_cacheWriteEn ),
       .io_addrLenAddr( ctrl_io_addrLenAddr ),
       .io_addrLenWriteData_addr( ctrl_io_addrLenWriteData_addr ),
       .io_addrLenWriteData_len( ctrl_io_addrLenWriteData_len ),
       .io_addrLenWriteEn_1( ctrl_io_addrLenWriteEn_1 ),
       .io_addrLenWriteEn_0( ctrl_io_addrLenWriteEn_0 ),
       .io_addrLenReadData_addr( lookup_io_addrLenReadData_addr ),
       .io_addrLenReadData_len( lookup_io_addrLenReadData_len ),
       .io_addrLenReadEn( ctrl_io_addrLenReadEn ),
       .io_keyLenAddr( ctrl_io_keyLenAddr ),
       .io_keyLenData( ctrl_io_keyLenData ),
       .io_keyLenWrite( ctrl_io_keyLenWrite ),
       .io_lock( ctrl_io_lock ),
       .io_halted( lookup_io_halted ),
       .io_writemode( ctrl_io_writemode ),
       .io_findAvailable( ctrl_io_findAvailable ),
       .io_resetCounts( ctrl_io_resetCounts ),
       .io_keyInfo_ready( lookup_io_writeKeyInfo_ready ),
       .io_keyInfo_valid( ctrl_io_keyInfo_valid ),
       .io_keyInfo_bits_len( ctrl_io_keyInfo_bits_len ),
       .io_keyInfo_bits_tag( ctrl_io_keyInfo_bits_tag ),
       .io_keyData_ready( lookup_io_writeKeyData_ready ),
       .io_keyData_valid( ctrl_io_keyData_valid ),
       .io_keyData_bits( ctrl_io_keyData_bits ),
       .io_hashSel_ready( ctrl_io_hashSel_ready ),
       .io_hashSel_valid( lookup_io_hashSel_valid ),
       .io_hashSel_bits_tag( lookup_io_hashSel_bits_tag ),
       .io_hashSel_bits_hash( lookup_io_hashSel_bits_hash ),
       .io_hashSel_bits_found( lookup_io_hashSel_bits_found ),
       .io_copyReq_ready( lookup_io_copyReq_ready ),
       .io_copyReq_valid( ctrl_io_copyReq_valid ),
       .io_copyReq_bits_hash( ctrl_io_copyReq_bits_hash ),
       .io_copyReq_bits_len( ctrl_io_copyReq_bits_len )
  );
endmodule

module StreamWriter(input clk, input reset,
    output io_stream_ready,
    input  io_stream_valid,
    input [7:0] io_stream_data,
    input  io_stream_last,
    output[7:0] io_writeData,
    output io_writeEn,
    input  io_enable,
    input  io_ignore,
    output[15:0] io_count,
    output io_finished
);

  reg  finished;
  wire T13;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [15:0] count;
  wire[15:0] T14;
  wire[15:0] T7;
  wire[15:0] T8;
  wire[15:0] T9;
  reg  writeEn;
  wire T15;
  wire T10;
  wire T11;
  reg [7:0] writeData;
  wire[7:0] T12;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    finished = {1{$random}};
    count = {1{$random}};
    writeEn = {1{$random}};
    writeData = {1{$random}};
  end
`endif

  assign io_finished = finished;
  assign T13 = reset ? 1'h1 : T0;
  assign T0 = T4 ? 1'h1 : T1;
  assign T1 = T2 ? 1'h0 : finished;
  assign T2 = T3 & finished;
  assign T3 = io_stream_valid & io_enable;
  assign T4 = T5 & io_stream_last;
  assign T5 = T3 & T6;
  assign T6 = finished ^ 1'h1;
  assign io_count = count;
  assign T14 = reset ? 16'h0 : T7;
  assign T7 = T5 ? T9 : T8;
  assign T8 = T2 ? 16'h1 : count;
  assign T9 = count + 16'h1;
  assign io_writeEn = writeEn;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T3 ? T11 : 1'h0;
  assign T11 = io_ignore ^ 1'h1;
  assign io_writeData = writeData;
  assign T12 = T3 ? io_stream_data : writeData;
  assign io_stream_ready = io_enable;

  always @(posedge clk) begin
    if(reset) begin
      finished <= 1'h1;
    end else if(T4) begin
      finished <= 1'h1;
    end else if(T2) begin
      finished <= 1'h0;
    end
    if(reset) begin
      count <= 16'h0;
    end else if(T5) begin
      count <= T9;
    end else if(T2) begin
      count <= 16'h1;
    end
    if(reset) begin
      writeEn <= 1'h0;
    end else if(T3) begin
      writeEn <= T11;
    end else begin
      writeEn <= 1'h0;
    end
    if(T3) begin
      writeData <= io_stream_data;
    end
  end
endmodule

module PacketBuffer(input clk, input reset,
    input  io_readData_ready,
    output io_readData_valid,
    output[7:0] io_readData_data,
    output io_readData_last,
    output io_stream_ready,
    input  io_stream_valid,
    input [15:0] io_stream_bits,
    output io_skip_ready,
    input  io_skip_valid,
    input [15:0] io_skip_bits,
    input [7:0] io_writeData,
    input  io_writeEn,
    output io_empty,
    output io_full
);

  wire T0;
  reg [15:0] readHead;
  wire[15:0] T42;
  wire[15:0] T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire T4;
  wire T5;
  reg [1:0] state;
  wire[1:0] T43;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg [15:0] readCount;
  wire[15:0] T44;
  wire[15:0] T19;
  wire[15:0] T20;
  wire[15:0] T21;
  wire[15:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire readValid;
  reg [15:0] writeHead;
  wire[15:0] T45;
  wire[15:0] T26;
  wire[15:0] T27;
  reg  writeEn;
  wire T28;
  wire[15:0] T29;
  wire T30;
  reg  skipValid;
  wire T31;
  wire[15:0] T32;
  wire T33;
  wire[15:0] T34;
  wire T35;
  wire ctrlReady;
  reg  readLast;
  wire T36;
  wire T37;
  reg [7:0] readData;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  reg [7:0] writeData;
  wire T41;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    readHead = {1{$random}};
    state = {1{$random}};
    readCount = {1{$random}};
    writeHead = {1{$random}};
    writeEn = {1{$random}};
    skipValid = {1{$random}};
    readLast = {1{$random}};
    readData = {1{$random}};
    writeData = {1{$random}};
  end
`endif

  assign io_full = T0;
  assign T0 = T34 == readHead;
  assign T42 = reset ? 16'h0 : T1;
  assign T1 = T30 ? T29 : T2;
  assign T2 = T4 ? T3 : readHead;
  assign T3 = readHead + 16'h1;
  assign T4 = T5 & io_readData_ready;
  assign T5 = 2'h1 == state;
  assign T43 = reset ? 2'h0 : T6;
  assign T6 = T30 ? 2'h0 : T7;
  assign T7 = T25 ? 2'h1 : T8;
  assign T8 = T23 ? 2'h2 : T9;
  assign T9 = T17 ? 2'h0 : T10;
  assign T10 = T14 ? 2'h2 : T11;
  assign T11 = T12 ? 2'h3 : state;
  assign T12 = T13 & io_skip_valid;
  assign T13 = 2'h0 == state;
  assign T14 = T13 & T15;
  assign T15 = T16 & io_stream_valid;
  assign T16 = io_skip_valid ^ 1'h1;
  assign T17 = T4 & T18;
  assign T18 = readCount == 16'h0;
  assign T44 = reset ? 16'h0 : T19;
  assign T19 = T25 ? T22 : T20;
  assign T20 = T14 ? io_stream_bits : T21;
  assign T21 = T12 ? io_skip_bits : readCount;
  assign T22 = readCount - 16'h1;
  assign T23 = T4 & T24;
  assign T24 = T18 ^ 1'h1;
  assign T25 = T28 & readValid;
  assign readValid = readHead != writeHead;
  assign T45 = reset ? 16'h0 : T26;
  assign T26 = writeEn ? T27 : writeHead;
  assign T27 = writeHead + 16'h1;
  assign T28 = 2'h2 == state;
  assign T29 = readHead + readCount;
  assign T30 = T33 & skipValid;
  assign T31 = readCount <= T32;
  assign T32 = writeHead - readHead;
  assign T33 = 2'h3 == state;
  assign T34 = writeHead + 16'h1;
  assign io_empty = T35;
  assign T35 = writeHead == readHead;
  assign io_skip_ready = ctrlReady;
  assign ctrlReady = state == 2'h0;
  assign io_stream_ready = ctrlReady;
  assign io_readData_last = readLast;
  assign T36 = T25 ? T37 : readLast;
  assign T37 = readCount == 16'h1;
  assign io_readData_data = readData;
  assign T38 = T25 ? T39 : readData;
  PacketBuffer_mem mem (
    .CLK(clk),
    .W0A(writeHead),
    .W0E(writeEn),
    .W0I(writeData),
    .R1A(T42),
    .R1E(1'h1),
    .R1O(T39)
  );
  assign io_readData_valid = T41;
  assign T41 = state == 2'h1;

  always @(posedge clk) begin
    if(reset) begin
      readHead <= 16'h0;
    end else if(T30) begin
      readHead <= T29;
    end else if(T4) begin
      readHead <= T3;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T30) begin
      state <= 2'h0;
    end else if(T25) begin
      state <= 2'h1;
    end else if(T23) begin
      state <= 2'h2;
    end else if(T17) begin
      state <= 2'h0;
    end else if(T14) begin
      state <= 2'h2;
    end else if(T12) begin
      state <= 2'h3;
    end
    if(reset) begin
      readCount <= 16'h0;
    end else if(T25) begin
      readCount <= T22;
    end else if(T14) begin
      readCount <= io_stream_bits;
    end else if(T12) begin
      readCount <= io_skip_bits;
    end
    if(reset) begin
      writeHead <= 16'h0;
    end else if(writeEn) begin
      writeHead <= T27;
    end
    writeEn <= io_writeEn;
    skipValid <= T31;
    if(T25) begin
      readLast <= T37;
    end
    if(T25) begin
      readData <= T39;
    end
    writeData <= io_writeData;
  end
endmodule

module StreamSplit(
    output io_in_ready,
    input  io_in_valid,
    input [7:0] io_in_data,
    input  io_in_last,
    input  io_out_a_ready,
    output io_out_a_valid,
    output[7:0] io_out_a_data,
    output io_out_a_last,
    input  io_out_b_ready,
    output io_out_b_valid,
    output[7:0] io_out_b_data,
    output io_out_b_last,
    input  io_sel
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_out_b_last = T0;
  assign T0 = io_in_last & io_sel;
  assign io_out_b_data = io_in_data;
  assign io_out_b_valid = T1;
  assign T1 = io_in_valid & io_sel;
  assign io_out_a_last = T2;
  assign T2 = io_in_last & T3;
  assign T3 = io_sel ^ 1'h1;
  assign io_out_a_data = io_in_data;
  assign io_out_a_valid = T4;
  assign T4 = io_in_valid & T5;
  assign T5 = io_sel ^ 1'h1;
  assign io_in_ready = T6;
  assign T6 = io_sel ? io_out_b_ready : io_out_a_ready;
endmodule

module StreamArbiter(input clk, input reset,
    output io_ins_1_ready,
    input  io_ins_1_valid,
    input [7:0] io_ins_1_data,
    input  io_ins_1_last,
    output io_ins_0_ready,
    input  io_ins_0_valid,
    input [7:0] io_ins_0_data,
    input  io_ins_0_last,
    input  io_out_ready,
    output io_out_valid,
    output[7:0] io_out_data,
    output io_out_last
);

  wire T0;
  wire T1;
  reg  sel;
  wire T25;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg  running;
  wire T26;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sel = {1{$random}};
    running = {1{$random}};
  end
`endif

  assign io_out_last = T0;
  assign T0 = T1 ? io_ins_1_last : io_ins_0_last;
  assign T1 = sel;
  assign T25 = reset ? 1'h0 : T2;
  assign T2 = T13 ? T12 : T3;
  assign T3 = T5 ? T4 : sel;
  assign T4 = sel + 1'h1;
  assign T5 = T8 & T6;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T1 ? io_ins_1_valid : io_ins_0_valid;
  assign T8 = running ^ 1'h1;
  assign T26 = reset ? 1'h0 : T9;
  assign T9 = T13 ? 1'h0 : T10;
  assign T10 = T11 ? 1'h1 : running;
  assign T11 = T8 & T7;
  assign T12 = sel + 1'h1;
  assign T13 = T16 & T14;
  assign T14 = T15 & io_out_ready;
  assign T15 = io_out_valid & io_out_last;
  assign T16 = T8 ^ 1'h1;
  assign io_out_data = T17;
  assign T17 = T1 ? io_ins_1_data : io_ins_0_data;
  assign io_out_valid = T18;
  assign T18 = T7 & running;
  assign io_ins_0_ready = T19;
  assign T19 = T20 & running;
  assign T20 = io_out_ready & T21;
  assign T21 = sel == 1'h0;
  assign io_ins_1_ready = T22;
  assign T22 = T23 & running;
  assign T23 = io_out_ready & T24;
  assign T24 = sel == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      sel <= 1'h0;
    end else if(T13) begin
      sel <= T12;
    end else if(T5) begin
      sel <= T4;
    end
    if(reset) begin
      running <= 1'h0;
    end else if(T13) begin
      running <= 1'h0;
    end else if(T11) begin
      running <= 1'h1;
    end
  end
endmodule

module ChecksumCompute(input clk, input reset,
    output io_data_ready,
    input  io_data_valid,
    input [7:0] io_data_bits,
    output io_len_ready,
    input  io_len_valid,
    input [15:0] io_len_bits,
    input  io_result_ready,
    output io_result_valid,
    output[15:0] io_result_bits
);

  wire[15:0] T0;
  reg [31:0] cursum;
  wire[31:0] T1;
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[31:0] T5;
  wire T6;
  wire T7;
  reg [2:0] state;
  wire[2:0] T51;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire T16;
  wire T17;
  wire T18;
  reg [15:0] length;
  wire[15:0] T19;
  wire[15:0] T20;
  wire[15:0] T21;
  wire[15:0] T22;
  wire[15:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[31:0] T32;
  wire[31:0] T52;
  wire[15:0] T33;
  wire T34;
  wire[31:0] T35;
  wire[31:0] T53;
  wire[15:0] T36;
  reg [7:0] highbyte;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire[31:0] T54;
  wire[15:0] T40;
  wire[15:0] T41;
  wire[15:0] T42;
  wire T43;
  wire[31:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cursum = {1{$random}};
    state = {1{$random}};
    length = {1{$random}};
    highbyte = {1{$random}};
  end
`endif

  assign io_result_bits = T0;
  assign T0 = cursum[4'hf:1'h0];
  assign T1 = T45 ? T44 : T2;
  assign T2 = T43 ? T54 : T3;
  assign T3 = T38 ? T35 : T4;
  assign T4 = T34 ? T32 : T5;
  assign T5 = T6 ? 32'h0 : cursum;
  assign T6 = T7 & io_len_valid;
  assign T7 = 3'h0 == state;
  assign T51 = reset ? 3'h0 : T8;
  assign T8 = T30 ? 3'h0 : T9;
  assign T9 = T45 ? 3'h5 : T10;
  assign T10 = T43 ? 3'h4 : T11;
  assign T11 = T28 ? 3'h1 : T12;
  assign T12 = T26 ? 3'h3 : T13;
  assign T13 = T16 ? 3'h2 : T14;
  assign T14 = T34 ? 3'h3 : T15;
  assign T15 = T6 ? 3'h1 : state;
  assign T16 = T24 & T17;
  assign T17 = T18 ^ 1'h1;
  assign T18 = length == 16'h1;
  assign T19 = T38 ? T23 : T20;
  assign T20 = T24 ? T22 : T21;
  assign T21 = T6 ? io_len_bits : length;
  assign T22 = length - 16'h1;
  assign T23 = length - 16'h1;
  assign T24 = T25 & io_data_valid;
  assign T25 = 3'h1 == state;
  assign T26 = T38 & T27;
  assign T27 = length == 16'h1;
  assign T28 = T38 & T29;
  assign T29 = T27 ^ 1'h1;
  assign T30 = T31 & io_result_ready;
  assign T31 = 3'h5 == state;
  assign T32 = cursum + T52;
  assign T52 = {16'h0, T33};
  assign T33 = {io_data_bits, 8'h0};
  assign T34 = T24 & T18;
  assign T35 = cursum + T53;
  assign T53 = {16'h0, T36};
  assign T36 = {highbyte, io_data_bits};
  assign T37 = T24 ? io_data_bits : highbyte;
  assign T38 = T39 & io_data_valid;
  assign T39 = 3'h2 == state;
  assign T54 = {16'h0, T40};
  assign T40 = T42 + T41;
  assign T41 = cursum[4'hf:1'h0];
  assign T42 = cursum[5'h1f:5'h10];
  assign T43 = 3'h3 == state;
  assign T44 = ~ cursum;
  assign T45 = 3'h4 == state;
  assign io_result_valid = T46;
  assign T46 = state == 3'h5;
  assign io_len_ready = T47;
  assign T47 = state == 3'h0;
  assign io_data_ready = T48;
  assign T48 = T50 | T49;
  assign T49 = state == 3'h2;
  assign T50 = state == 3'h1;

  always @(posedge clk) begin
    if(T45) begin
      cursum <= T44;
    end else if(T43) begin
      cursum <= T54;
    end else if(T38) begin
      cursum <= T35;
    end else if(T34) begin
      cursum <= T32;
    end else if(T6) begin
      cursum <= 32'h0;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T30) begin
      state <= 3'h0;
    end else if(T45) begin
      state <= 3'h5;
    end else if(T43) begin
      state <= 3'h4;
    end else if(T28) begin
      state <= 3'h1;
    end else if(T26) begin
      state <= 3'h3;
    end else if(T16) begin
      state <= 3'h2;
    end else if(T34) begin
      state <= 3'h3;
    end else if(T6) begin
      state <= 3'h1;
    end
    if(T38) begin
      length <= T23;
    end else if(T24) begin
      length <= T22;
    end else if(T6) begin
      length <= io_len_bits;
    end
    if(T24) begin
      highbyte <= io_data_bits;
    end
  end
endmodule

module Responder(input clk, input reset,
    input  io_temac_tx_ready,
    output io_temac_tx_valid,
    output[7:0] io_temac_tx_data,
    output io_temac_tx_last,
    output io_resultData_ready,
    input  io_resultData_valid,
    input [7:0] io_resultData_bits,
    input [15:0] io_resLen,
    input [31:0] io_pktRoute_srcAddr,
    input [31:0] io_pktRoute_dstAddr,
    input [15:0] io_pktRoute_srcPort,
    input [15:0] io_pktRoute_dstPort,
    input [15:0] io_pktRoute_reqId,
    input [7:0] io_pktRoute_dstMac_5,
    input [7:0] io_pktRoute_dstMac_4,
    input [7:0] io_pktRoute_dstMac_3,
    input [7:0] io_pktRoute_dstMac_2,
    input [7:0] io_pktRoute_dstMac_1,
    input [7:0] io_pktRoute_dstMac_0,
    input [7:0] io_pktRoute_srcMac_5,
    input [7:0] io_pktRoute_srcMac_4,
    input [7:0] io_pktRoute_srcMac_3,
    input [7:0] io_pktRoute_srcMac_2,
    input [7:0] io_pktRoute_srcMac_1,
    input [7:0] io_pktRoute_srcMac_0,
    input  io_start,
    output io_ready
);

  wire T317;
  wire T318;
  reg [3:0] state;
  wire[3:0] T311;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [15:0] pktLen;
  wire[15:0] T20;
  wire[15:0] T21;
  wire[15:0] T22;
  wire[15:0] T23;
  wire[15:0] udpPktLen;
  wire[15:0] T312;
  reg [5:0] headerIndex;
  wire[5:0] T24;
  wire[5:0] T25;
  wire[5:0] T26;
  wire[5:0] T27;
  wire[5:0] T28;
  wire[5:0] T29;
  wire[5:0] T30;
  wire[5:0] T31;
  wire[5:0] T32;
  wire[5:0] T33;
  wire[5:0] T34;
  wire[5:0] T35;
  wire[5:0] T36;
  wire T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[15:0] T56;
  reg [15:0] bodyIndex;
  wire[15:0] T57;
  wire[15:0] T58;
  wire[15:0] T59;
  wire[15:0] T60;
  wire[15:0] T61;
  wire[15:0] T62;
  wire T63;
  wire T64;
  wire[15:0] T65;
  wire[15:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [3:0] ethHeaderIndex;
  wire[3:0] T79;
  wire[3:0] T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  reg [7:0] pktData;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] pseudoHeaderData;
  wire[7:0] T108;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T119;
  wire[7:0] T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire[7:0] T127;
  wire[7:0] T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire[7:0] T131;
  wire[7:0] T132;
  wire[7:0] T133;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire T137;
  wire[7:0] T138;
  wire T139;
  wire[7:0] T140;
  wire T141;
  wire[7:0] T142;
  wire T143;
  wire[7:0] T144;
  wire T145;
  wire[7:0] T146;
  wire T147;
  wire[7:0] T148;
  wire T149;
  wire[7:0] T150;
  wire T151;
  wire T152;
  wire[7:0] T153;
  wire T154;
  wire[7:0] T155;
  wire T156;
  wire[7:0] T157;
  wire T158;
  wire[7:0] T159;
  wire T160;
  wire[7:0] T161;
  wire T162;
  wire[7:0] T163;
  wire T164;
  wire[7:0] T165;
  wire T166;
  wire[7:0] T167;
  wire T168;
  wire[7:0] T169;
  wire T170;
  wire[7:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire[7:0] T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[7:0] ethHeaderData;
  wire[7:0] T185;
  wire[7:0] T186;
  wire[7:0] T187;
  wire[7:0] T188;
  wire[7:0] T189;
  wire[7:0] T190;
  wire[7:0] T191;
  wire[7:0] T192;
  wire[7:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[7:0] T196;
  wire[7:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire[7:0] headerData;
  wire[7:0] T211;
  wire[7:0] T212;
  wire[7:0] T213;
  wire[7:0] T214;
  wire[7:0] T215;
  wire[7:0] T216;
  wire[7:0] T217;
  wire[7:0] T218;
  wire[7:0] T219;
  wire[7:0] T220;
  wire[7:0] T221;
  wire[7:0] T222;
  wire[7:0] T223;
  wire[7:0] T224;
  wire[7:0] T225;
  wire[7:0] T226;
  wire[7:0] T227;
  wire[7:0] T228;
  wire[7:0] T229;
  wire[7:0] T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire[7:0] T240;
  wire[7:0] T241;
  wire[7:0] T242;
  wire[7:0] T243;
  wire[7:0] T314;
  wire[6:0] T244;
  wire T245;
  wire[7:0] T246;
  wire[15:0] ipPktLen;
  wire T247;
  wire[7:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire[7:0] T252;
  reg [15:0] ipChecksum;
  wire[15:0] T253;
  wire T254;
  wire[7:0] T255;
  wire T256;
  wire[7:0] T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire[7:0] T261;
  wire T262;
  wire[7:0] T263;
  wire T264;
  wire[7:0] T265;
  wire T266;
  wire[7:0] T267;
  wire T268;
  wire[7:0] T269;
  wire T270;
  wire[7:0] T271;
  wire T272;
  wire[7:0] T273;
  wire T274;
  wire[7:0] T275;
  wire T276;
  wire[7:0] T277;
  wire T278;
  wire[7:0] T279;
  wire T280;
  wire[7:0] T281;
  wire T282;
  wire[7:0] T283;
  wire T284;
  wire[7:0] T285;
  reg [15:0] udpChecksum;
  wire[15:0] T286;
  wire T287;
  wire[7:0] T288;
  wire T289;
  wire[7:0] T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[7:0] T297;
  wire T298;
  wire[7:0] T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire[7:0] bodyData;
  reg [7:0] buffer [4095:0];
  wire[7:0] T305;
  wire[11:0] T315;
  wire[11:0] T316;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T0;
  wire T90;
  wire T91;
  wire T92;
  reg  pktLast;
  wire T313;
  wire T93;
  wire T94;
  wire[15:0] T95;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire csCompute_io_len_ready;
  wire csCompute_io_result_valid;
  wire[15:0] csCompute_io_result_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    pktLen = {1{$random}};
    headerIndex = {1{$random}};
    bodyIndex = {1{$random}};
    ethHeaderIndex = {1{$random}};
    pktData = {1{$random}};
    ipChecksum = {1{$random}};
    udpChecksum = {1{$random}};
    for (initvar = 0; initvar < 4096; initvar = initvar+1)
      buffer[initvar] = {1{$random}};
    pktLast = {1{$random}};
  end
`endif

  assign T317 = T319 | T318;
  assign T318 = state == 4'h8;
  assign T311 = reset ? 4'h0 : T1;
  assign T1 = T89 ? 4'h0 : T2;
  assign T2 = T88 ? 4'hb : T3;
  assign T3 = T77 ? 4'ha : T4;
  assign T4 = T75 ? 4'h9 : T5;
  assign T5 = T73 ? 4'h6 : T6;
  assign T6 = T54 ? 4'h8 : T7;
  assign T7 = T52 ? 4'h7 : T8;
  assign T8 = T50 ? 4'h6 : T9;
  assign T9 = T48 ? 4'h5 : T10;
  assign T10 = T46 ? 4'h4 : T11;
  assign T11 = T18 ? 4'h3 : T12;
  assign T12 = T16 ? 4'h2 : T13;
  assign T13 = T14 ? 4'h1 : state;
  assign T14 = T15 & io_start;
  assign T15 = 4'h0 == state;
  assign T16 = T17 & csCompute_io_len_ready;
  assign T17 = 4'h1 == state;
  assign T18 = T45 & T19;
  assign T19 = T312 == pktLen;
  assign T20 = T75 ? io_resLen : T21;
  assign T21 = T46 ? T23 : T22;
  assign T22 = T14 ? 16'h14 : pktLen;
  assign T23 = udpPktLen + 16'hc;
  assign udpPktLen = io_resLen + 16'h2c;
  assign T312 = {10'h0, headerIndex};
  assign T24 = T40 ? T39 : T25;
  assign T25 = T77 ? T38 : T26;
  assign T26 = T54 ? 6'h0 : T27;
  assign T27 = T37 ? T36 : T28;
  assign T28 = T48 ? T35 : T29;
  assign T29 = T46 ? 6'h0 : T30;
  assign T30 = T45 ? T34 : T31;
  assign T31 = T16 ? T33 : T32;
  assign T32 = T14 ? 6'h0 : headerIndex;
  assign T33 = headerIndex + 6'h1;
  assign T34 = headerIndex + 6'h1;
  assign T35 = headerIndex + 6'h1;
  assign T36 = headerIndex + 6'h1;
  assign T37 = 4'h5 == state;
  assign T38 = headerIndex + 6'h1;
  assign T39 = headerIndex + 6'h1;
  assign T40 = T43 & T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = headerIndex == 6'h0;
  assign T43 = T44 & io_temac_tx_ready;
  assign T44 = 4'ha == state;
  assign T45 = 4'h2 == state;
  assign T46 = T47 & csCompute_io_result_valid;
  assign T47 = 4'h3 == state;
  assign T48 = T49 & csCompute_io_len_ready;
  assign T49 = 4'h4 == state;
  assign T50 = T37 & T51;
  assign T51 = headerIndex == 6'h38;
  assign T52 = T53 & io_resultData_valid;
  assign T53 = 4'h6 == state;
  assign T54 = T72 & T55;
  assign T55 = bodyIndex == T56;
  assign T56 = io_resLen - 16'h1;
  assign T57 = T67 ? T66 : T58;
  assign T58 = T88 ? T65 : T59;
  assign T59 = T75 ? 16'h0 : T60;
  assign T60 = T63 ? T62 : T61;
  assign T61 = T50 ? 16'h0 : bodyIndex;
  assign T62 = bodyIndex + 16'h1;
  assign T63 = T72 & T64;
  assign T64 = T55 ^ 1'h1;
  assign T65 = bodyIndex + 16'h1;
  assign T66 = bodyIndex + 16'h1;
  assign T67 = T70 & T68;
  assign T68 = T69 ^ 1'h1;
  assign T69 = bodyIndex == pktLen;
  assign T70 = T71 & io_temac_tx_ready;
  assign T71 = 4'hb == state;
  assign T72 = 4'h7 == state;
  assign T73 = T63 & T74;
  assign T74 = io_resultData_valid ^ 1'h1;
  assign T75 = T76 & csCompute_io_result_valid;
  assign T76 = 4'h8 == state;
  assign T77 = T86 & T78;
  assign T78 = ethHeaderIndex == 4'he;
  assign T79 = T84 ? T83 : T80;
  assign T80 = T75 ? T82 : T81;
  assign T81 = T14 ? 4'h0 : ethHeaderIndex;
  assign T82 = ethHeaderIndex + 4'h1;
  assign T83 = ethHeaderIndex + 4'h1;
  assign T84 = T86 & T85;
  assign T85 = T78 ^ 1'h1;
  assign T86 = T87 & io_temac_tx_ready;
  assign T87 = 4'h9 == state;
  assign T88 = T43 & T42;
  assign T89 = T70 & T69;
  assign T319 = state == 4'h3;
  assign T320 = T322 | T321;
  assign T321 = state == 4'h4;
  assign T322 = state == 4'h1;
  assign T96 = T67 ? bodyData : T97;
  assign T97 = T40 ? headerData : T98;
  assign T98 = T88 ? bodyData : T99;
  assign T99 = T84 ? ethHeaderData : T100;
  assign T100 = T77 ? headerData : T101;
  assign T101 = T75 ? ethHeaderData : T102;
  assign T102 = T184 ? io_resultData_bits : T103;
  assign T103 = T52 ? io_resultData_bits : T104;
  assign T104 = T37 ? pseudoHeaderData : T105;
  assign T105 = T48 ? pseudoHeaderData : T106;
  assign T106 = T45 ? headerData : T107;
  assign T107 = T16 ? headerData : pktData;
  assign pseudoHeaderData = T108;
  assign T108 = T183 ? 8'hef : T109;
  assign T109 = T182 ? 8'hbe : T110;
  assign T110 = T181 ? 8'had : T111;
  assign T111 = T180 ? 8'hde : T112;
  assign T112 = T179 ? T178 : T113;
  assign T113 = T177 ? T176 : T114;
  assign T114 = T175 ? 8'h4 : T115;
  assign T115 = T174 ? 8'h81 : T116;
  assign T116 = T173 ? 8'h1 : T117;
  assign T117 = T172 ? T171 : T118;
  assign T118 = T170 ? T169 : T119;
  assign T119 = T168 ? T167 : T120;
  assign T120 = T166 ? T165 : T121;
  assign T121 = T164 ? T163 : T122;
  assign T122 = T162 ? T161 : T123;
  assign T123 = T160 ? T159 : T124;
  assign T124 = T158 ? T157 : T125;
  assign T125 = T156 ? T155 : T126;
  assign T126 = T154 ? T153 : T127;
  assign T127 = T152 ? 8'h11 : T128;
  assign T128 = T151 ? T150 : T129;
  assign T129 = T149 ? T148 : T130;
  assign T130 = T147 ? T146 : T131;
  assign T131 = T145 ? T144 : T132;
  assign T132 = T143 ? T142 : T133;
  assign T133 = T141 ? T140 : T134;
  assign T134 = T139 ? T138 : T135;
  assign T135 = T137 ? T136 : 8'h0;
  assign T136 = io_pktRoute_dstAddr[5'h1f:5'h18];
  assign T137 = 6'h0 == headerIndex;
  assign T138 = io_pktRoute_dstAddr[5'h17:5'h10];
  assign T139 = 6'h1 == headerIndex;
  assign T140 = io_pktRoute_dstAddr[4'hf:4'h8];
  assign T141 = 6'h2 == headerIndex;
  assign T142 = io_pktRoute_dstAddr[3'h7:1'h0];
  assign T143 = 6'h3 == headerIndex;
  assign T144 = io_pktRoute_srcAddr[5'h1f:5'h18];
  assign T145 = 6'h4 == headerIndex;
  assign T146 = io_pktRoute_srcAddr[5'h17:5'h10];
  assign T147 = 6'h5 == headerIndex;
  assign T148 = io_pktRoute_srcAddr[4'hf:4'h8];
  assign T149 = 6'h6 == headerIndex;
  assign T150 = io_pktRoute_srcAddr[3'h7:1'h0];
  assign T151 = 6'h7 == headerIndex;
  assign T152 = 6'h9 == headerIndex;
  assign T153 = udpPktLen[4'hf:4'h8];
  assign T154 = 6'ha == headerIndex;
  assign T155 = udpPktLen[3'h7:1'h0];
  assign T156 = 6'hb == headerIndex;
  assign T157 = io_pktRoute_dstPort[4'hf:4'h8];
  assign T158 = 6'hc == headerIndex;
  assign T159 = io_pktRoute_dstPort[3'h7:1'h0];
  assign T160 = 6'hd == headerIndex;
  assign T161 = io_pktRoute_srcPort[4'hf:4'h8];
  assign T162 = 6'he == headerIndex;
  assign T163 = io_pktRoute_srcPort[3'h7:1'h0];
  assign T164 = 6'hf == headerIndex;
  assign T165 = udpPktLen[4'hf:4'h8];
  assign T166 = 6'h10 == headerIndex;
  assign T167 = udpPktLen[3'h7:1'h0];
  assign T168 = 6'h11 == headerIndex;
  assign T169 = io_pktRoute_reqId[4'hf:4'h8];
  assign T170 = 6'h14 == headerIndex;
  assign T171 = io_pktRoute_reqId[3'h7:1'h0];
  assign T172 = 6'h15 == headerIndex;
  assign T173 = 6'h19 == headerIndex;
  assign T174 = 6'h1c == headerIndex;
  assign T175 = 6'h20 == headerIndex;
  assign T176 = io_resLen[4'hf:4'h8];
  assign T177 = 6'h26 == headerIndex;
  assign T178 = io_resLen[3'h7:1'h0];
  assign T179 = 6'h27 == headerIndex;
  assign T180 = 6'h34 == headerIndex;
  assign T181 = 6'h35 == headerIndex;
  assign T182 = 6'h36 == headerIndex;
  assign T183 = 6'h37 == headerIndex;
  assign T184 = T63 & io_resultData_valid;
  assign ethHeaderData = T185;
  assign T185 = T210 ? 8'h8 : T186;
  assign T186 = T209 ? io_pktRoute_dstMac_5 : T187;
  assign T187 = T208 ? io_pktRoute_dstMac_4 : T188;
  assign T188 = T207 ? io_pktRoute_dstMac_3 : T189;
  assign T189 = T206 ? io_pktRoute_dstMac_2 : T190;
  assign T190 = T205 ? io_pktRoute_dstMac_1 : T191;
  assign T191 = T204 ? io_pktRoute_dstMac_0 : T192;
  assign T192 = T203 ? io_pktRoute_srcMac_5 : T193;
  assign T193 = T202 ? io_pktRoute_srcMac_4 : T194;
  assign T194 = T201 ? io_pktRoute_srcMac_3 : T195;
  assign T195 = T200 ? io_pktRoute_srcMac_2 : T196;
  assign T196 = T199 ? io_pktRoute_srcMac_1 : T197;
  assign T197 = T198 ? io_pktRoute_srcMac_0 : 8'h0;
  assign T198 = 4'h0 == ethHeaderIndex;
  assign T199 = 4'h1 == ethHeaderIndex;
  assign T200 = 4'h2 == ethHeaderIndex;
  assign T201 = 4'h3 == ethHeaderIndex;
  assign T202 = 4'h4 == ethHeaderIndex;
  assign T203 = 4'h5 == ethHeaderIndex;
  assign T204 = 4'h6 == ethHeaderIndex;
  assign T205 = 4'h7 == ethHeaderIndex;
  assign T206 = 4'h8 == ethHeaderIndex;
  assign T207 = 4'h9 == ethHeaderIndex;
  assign T208 = 4'ha == ethHeaderIndex;
  assign T209 = 4'hb == ethHeaderIndex;
  assign T210 = 4'hc == ethHeaderIndex;
  assign headerData = T211;
  assign T211 = T304 ? 8'hef : T212;
  assign T212 = T303 ? 8'hbe : T213;
  assign T213 = T302 ? 8'had : T214;
  assign T214 = T301 ? 8'hde : T215;
  assign T215 = T300 ? T299 : T216;
  assign T216 = T298 ? T297 : T217;
  assign T217 = T296 ? 8'h4 : T218;
  assign T218 = T295 ? 8'h81 : T219;
  assign T219 = T294 ? 8'h1 : T220;
  assign T220 = T293 ? T292 : T221;
  assign T221 = T291 ? T290 : T222;
  assign T222 = T289 ? T288 : T223;
  assign T223 = T287 ? T285 : T224;
  assign T224 = T284 ? T283 : T225;
  assign T225 = T282 ? T281 : T226;
  assign T226 = T280 ? T279 : T227;
  assign T227 = T278 ? T277 : T228;
  assign T228 = T276 ? T275 : T229;
  assign T229 = T274 ? T273 : T230;
  assign T230 = T272 ? T271 : T231;
  assign T231 = T270 ? T269 : T232;
  assign T232 = T268 ? T267 : T233;
  assign T233 = T266 ? T265 : T234;
  assign T234 = T264 ? T263 : T235;
  assign T235 = T262 ? T261 : T236;
  assign T236 = T260 ? T259 : T237;
  assign T237 = T258 ? T257 : T238;
  assign T238 = T256 ? T255 : T239;
  assign T239 = T254 ? T252 : T240;
  assign T240 = T251 ? 8'h11 : T241;
  assign T241 = T250 ? 8'h64 : T242;
  assign T242 = T249 ? T248 : T243;
  assign T243 = T247 ? T246 : T314;
  assign T314 = {1'h0, T244};
  assign T244 = T245 ? 7'h45 : 7'h0;
  assign T245 = 6'h0 == headerIndex;
  assign T246 = ipPktLen[4'hf:4'h8];
  assign ipPktLen = io_resLen + 16'h40;
  assign T247 = 6'h2 == headerIndex;
  assign T248 = ipPktLen[3'h7:1'h0];
  assign T249 = 6'h3 == headerIndex;
  assign T250 = 6'h8 == headerIndex;
  assign T251 = 6'h9 == headerIndex;
  assign T252 = ipChecksum[4'hf:4'h8];
  assign T253 = T46 ? csCompute_io_result_bits : ipChecksum;
  assign T254 = 6'ha == headerIndex;
  assign T255 = ipChecksum[3'h7:1'h0];
  assign T256 = 6'hb == headerIndex;
  assign T257 = io_pktRoute_dstAddr[5'h1f:5'h18];
  assign T258 = 6'hc == headerIndex;
  assign T259 = io_pktRoute_dstAddr[5'h17:5'h10];
  assign T260 = 6'hd == headerIndex;
  assign T261 = io_pktRoute_dstAddr[4'hf:4'h8];
  assign T262 = 6'he == headerIndex;
  assign T263 = io_pktRoute_dstAddr[3'h7:1'h0];
  assign T264 = 6'hf == headerIndex;
  assign T265 = io_pktRoute_srcAddr[5'h1f:5'h18];
  assign T266 = 6'h10 == headerIndex;
  assign T267 = io_pktRoute_srcAddr[5'h17:5'h10];
  assign T268 = 6'h11 == headerIndex;
  assign T269 = io_pktRoute_srcAddr[4'hf:4'h8];
  assign T270 = 6'h12 == headerIndex;
  assign T271 = io_pktRoute_srcAddr[3'h7:1'h0];
  assign T272 = 6'h13 == headerIndex;
  assign T273 = io_pktRoute_dstPort[4'hf:4'h8];
  assign T274 = 6'h14 == headerIndex;
  assign T275 = io_pktRoute_dstPort[3'h7:1'h0];
  assign T276 = 6'h15 == headerIndex;
  assign T277 = io_pktRoute_srcPort[4'hf:4'h8];
  assign T278 = 6'h16 == headerIndex;
  assign T279 = io_pktRoute_srcPort[3'h7:1'h0];
  assign T280 = 6'h17 == headerIndex;
  assign T281 = udpPktLen[4'hf:4'h8];
  assign T282 = 6'h18 == headerIndex;
  assign T283 = udpPktLen[3'h7:1'h0];
  assign T284 = 6'h19 == headerIndex;
  assign T285 = udpChecksum[4'hf:4'h8];
  assign T286 = T75 ? csCompute_io_result_bits : udpChecksum;
  assign T287 = 6'h1a == headerIndex;
  assign T288 = udpChecksum[3'h7:1'h0];
  assign T289 = 6'h1b == headerIndex;
  assign T290 = io_pktRoute_reqId[4'hf:4'h8];
  assign T291 = 6'h1c == headerIndex;
  assign T292 = io_pktRoute_reqId[3'h7:1'h0];
  assign T293 = 6'h1d == headerIndex;
  assign T294 = 6'h21 == headerIndex;
  assign T295 = 6'h24 == headerIndex;
  assign T296 = 6'h28 == headerIndex;
  assign T297 = io_resLen[4'hf:4'h8];
  assign T298 = 6'h2e == headerIndex;
  assign T299 = io_resLen[3'h7:1'h0];
  assign T300 = 6'h2f == headerIndex;
  assign T301 = 6'h3c == headerIndex;
  assign T302 = 6'h3d == headerIndex;
  assign T303 = 6'h3e == headerIndex;
  assign T304 = 6'h3f == headerIndex;
  assign bodyData = buffer[T316];
  assign T315 = bodyIndex[4'hb:1'h0];
  assign T316 = bodyIndex[4'hb:1'h0];
  assign T323 = T325 | T324;
  assign T324 = state == 4'h7;
  assign T325 = T327 | T326;
  assign T326 = state == 4'h5;
  assign T327 = state == 4'h2;
  assign io_ready = T0;
  assign T0 = state == 4'h0;
  assign io_resultData_ready = T90;
  assign T90 = T92 | T91;
  assign T91 = state == 4'h7;
  assign T92 = state == 4'h6;
  assign io_temac_tx_last = pktLast;
  assign T313 = reset ? 1'h0 : T93;
  assign T93 = T67 ? T94 : pktLast;
  assign T94 = bodyIndex == T95;
  assign T95 = io_resLen - 16'h1;
  assign io_temac_tx_data = pktData;
  assign io_temac_tx_valid = T306;
  assign T306 = T308 | T307;
  assign T307 = state == 4'hb;
  assign T308 = T310 | T309;
  assign T309 = state == 4'ha;
  assign T310 = state == 4'h9;
  ChecksumCompute csCompute(.clk(clk), .reset(reset),
       //.io_data_ready(  )
       .io_data_valid( T323 ),
       .io_data_bits( pktData ),
       .io_len_ready( csCompute_io_len_ready ),
       .io_len_valid( T320 ),
       .io_len_bits( pktLen ),
       .io_result_ready( T317 ),
       .io_result_valid( csCompute_io_result_valid ),
       .io_result_bits( csCompute_io_result_bits )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T89) begin
      state <= 4'h0;
    end else if(T88) begin
      state <= 4'hb;
    end else if(T77) begin
      state <= 4'ha;
    end else if(T75) begin
      state <= 4'h9;
    end else if(T73) begin
      state <= 4'h6;
    end else if(T54) begin
      state <= 4'h8;
    end else if(T52) begin
      state <= 4'h7;
    end else if(T50) begin
      state <= 4'h6;
    end else if(T48) begin
      state <= 4'h5;
    end else if(T46) begin
      state <= 4'h4;
    end else if(T18) begin
      state <= 4'h3;
    end else if(T16) begin
      state <= 4'h2;
    end else if(T14) begin
      state <= 4'h1;
    end
    if(T75) begin
      pktLen <= io_resLen;
    end else if(T46) begin
      pktLen <= T23;
    end else if(T14) begin
      pktLen <= 16'h14;
    end
    if(T40) begin
      headerIndex <= T39;
    end else if(T77) begin
      headerIndex <= T38;
    end else if(T54) begin
      headerIndex <= 6'h0;
    end else if(T37) begin
      headerIndex <= T36;
    end else if(T48) begin
      headerIndex <= T35;
    end else if(T46) begin
      headerIndex <= 6'h0;
    end else if(T45) begin
      headerIndex <= T34;
    end else if(T16) begin
      headerIndex <= T33;
    end else if(T14) begin
      headerIndex <= 6'h0;
    end
    if(T67) begin
      bodyIndex <= T66;
    end else if(T88) begin
      bodyIndex <= T65;
    end else if(T75) begin
      bodyIndex <= 16'h0;
    end else if(T63) begin
      bodyIndex <= T62;
    end else if(T50) begin
      bodyIndex <= 16'h0;
    end
    if(T84) begin
      ethHeaderIndex <= T83;
    end else if(T75) begin
      ethHeaderIndex <= T82;
    end else if(T14) begin
      ethHeaderIndex <= 4'h0;
    end
    if(T67) begin
      pktData <= bodyData;
    end else if(T40) begin
      pktData <= headerData;
    end else if(T88) begin
      pktData <= bodyData;
    end else if(T84) begin
      pktData <= ethHeaderData;
    end else if(T77) begin
      pktData <= headerData;
    end else if(T75) begin
      pktData <= ethHeaderData;
    end else if(T184) begin
      pktData <= io_resultData_bits;
    end else if(T52) begin
      pktData <= io_resultData_bits;
    end else if(T37) begin
      pktData <= pseudoHeaderData;
    end else if(T48) begin
      pktData <= pseudoHeaderData;
    end else if(T45) begin
      pktData <= headerData;
    end else if(T16) begin
      pktData <= headerData;
    end
    if(T46) begin
      ipChecksum <= csCompute_io_result_bits;
    end
    if(T75) begin
      udpChecksum <= csCompute_io_result_bits;
    end
    if (T72)
      buffer[T315] <= pktData;
    if(reset) begin
      pktLast <= 1'h0;
    end else if(T67) begin
      pktLast <= T94;
    end
  end
endmodule

module PacketFilter(input clk, input reset,
    output io_temac_rx_ready,
    input  io_temac_rx_valid,
    input [7:0] io_temac_rx_data,
    input  io_temac_rx_last,
    input  io_core_rx_ready,
    output io_core_rx_valid,
    output[7:0] io_core_rx_data,
    output io_core_rx_last,
    input  io_temac_tx_ready,
    output io_temac_tx_valid,
    output[7:0] io_temac_tx_data,
    output io_temac_tx_last,
    output io_core_tx_ready,
    input  io_core_tx_valid,
    input [7:0] io_core_tx_data,
    input  io_core_tx_last,
    input  io_keyInfo_ready,
    output io_keyInfo_valid,
    output[7:0] io_keyInfo_bits_len,
    output[3:0] io_keyInfo_bits_tag,
    input  io_keyData_ready,
    output io_keyData_valid,
    output[7:0] io_keyData_bits,
    output io_resultInfo_ready,
    input  io_resultInfo_valid,
    input [18:0] io_resultInfo_bits_len,
    input [3:0] io_resultInfo_bits_tag,
    output io_resultData_ready,
    input  io_resultData_valid,
    input [7:0] io_resultData_bits,
    input  io_readready
);

  wire T281;
  reg [2:0] d_state;
  wire[2:0] T265;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [7:0] resLen;
  wire[7:0] T266;
  wire[18:0] T11;
  wire[18:0] T267;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg [7:0] reqPktRoute_srcMac_0;
  wire[7:0] T282;
  wire[7:0] T283;
  wire[207:0] T284;
  wire[207:0] T285;
  wire[207:0] T286;
  wire[207:0] T287;
  wire[71:0] T288;
  wire[39:0] T289;
  wire[23:0] T290;
  wire[15:0] T291;
  wire[7:0] curRoute_srcMac_0;
  reg [7:0] srcMac_0;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire[7:0] T295;
  wire[2:0] T296;
  reg [2:0] macIndex;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T81;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg [5:0] m_state;
  wire[5:0] T268;
  wire[5:0] T23;
  wire[5:0] T24;
  wire[5:0] T25;
  wire[5:0] T26;
  wire[5:0] T27;
  wire[5:0] T28;
  wire[5:0] T29;
  wire[5:0] T30;
  wire[5:0] T31;
  wire[5:0] T32;
  wire[5:0] T33;
  wire[5:0] T34;
  wire[5:0] T35;
  wire[5:0] T36;
  wire[5:0] T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[5:0] T46;
  wire[5:0] T47;
  wire[5:0] T48;
  wire[5:0] T49;
  wire[5:0] T50;
  wire[5:0] T51;
  wire[5:0] T52;
  wire[5:0] T53;
  wire[5:0] T54;
  wire[5:0] T55;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire[5:0] T59;
  wire[5:0] T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] T65;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[5:0] T69;
  wire[5:0] T70;
  wire[5:0] T71;
  wire T93;
  wire T88;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[15:0] T99;
  reg [7:0] etherTypeHigh;
  wire[7:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[3:0] T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  reg [15:0] lenOffset;
  wire[15:0] T120;
  wire[15:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  reg  ipv6;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[15:0] T269;
  reg [7:0] headerLen;
  wire[7:0] T270;
  wire[7:0] T148;
  wire[7:0] T149;
  wire[7:0] T150;
  wire[7:0] T151;
  wire[7:0] T152;
  wire[7:0] T153;
  wire[7:0] T154;
  wire[7:0] T155;
  wire[7:0] T156;
  wire[7:0] T271;
  wire[5:0] T157;
  wire[3:0] T158;
  wire[7:0] T159;
  wire[7:0] T160;
  wire[7:0] T161;
  wire[7:0] T162;
  wire[7:0] T163;
  wire[7:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[15:0] T272;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[15:0] T273;
  wire T184;
  wire T185;
  wire T186;
  wire[15:0] T274;
  reg [15:0] pktLen;
  wire[15:0] T275;
  wire[15:0] T187;
  wire[15:0] T188;
  wire[15:0] T189;
  wire[15:0] T190;
  wire[15:0] T191;
  wire[15:0] T192;
  wire[15:0] T193;
  wire[7:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire[15:0] T276;
  wire T203;
  wire T204;
  wire T205;
  wire[15:0] T277;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire[15:0] T278;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T76;
  wire T77;
  wire T91;
  wire T92;
  wire[2:0] T82;
  wire T83;
  wire T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T89;
  wire T90;
  wire[7:0] curRoute_srcMac_1;
  reg [7:0] srcMac_1;
  wire[7:0] T297;
  wire T298;
  wire T299;
  wire[7:0] curRoute_srcMac_2;
  reg [7:0] srcMac_2;
  wire[7:0] T300;
  wire T301;
  wire T302;
  wire[15:0] T303;
  wire[7:0] curRoute_srcMac_3;
  reg [7:0] srcMac_3;
  wire[7:0] T304;
  wire T305;
  wire T306;
  wire[7:0] curRoute_srcMac_4;
  reg [7:0] srcMac_4;
  wire[7:0] T307;
  wire T308;
  wire T309;
  wire[31:0] T310;
  wire[15:0] T311;
  wire[7:0] curRoute_srcMac_5;
  reg [7:0] srcMac_5;
  wire[7:0] T312;
  wire T313;
  wire T314;
  wire[7:0] curRoute_dstMac_0;
  reg [7:0] dstMac_0;
  wire[7:0] T315;
  wire T316;
  wire T317;
  wire[7:0] T318;
  wire[2:0] T319;
  wire[15:0] T320;
  wire[7:0] curRoute_dstMac_1;
  reg [7:0] dstMac_1;
  wire[7:0] T321;
  wire T322;
  wire T323;
  wire[7:0] curRoute_dstMac_2;
  reg [7:0] dstMac_2;
  wire[7:0] T324;
  wire T325;
  wire T326;
  wire[135:0] T327;
  wire[39:0] T328;
  wire[15:0] T329;
  wire[7:0] curRoute_dstMac_3;
  reg [7:0] dstMac_3;
  wire[7:0] T330;
  wire T331;
  wire T332;
  wire[7:0] curRoute_dstMac_4;
  reg [7:0] dstMac_4;
  wire[7:0] T333;
  wire T334;
  wire T335;
  wire[23:0] T336;
  wire[7:0] curRoute_dstMac_5;
  reg [7:0] dstMac_5;
  wire[7:0] T337;
  wire T338;
  wire T339;
  wire[15:0] curRoute_reqId;
  reg [15:0] reqId;
  wire[15:0] T340;
  wire[15:0] T341;
  wire[15:0] T342;
  wire[15:0] T343;
  wire[7:0] T344;
  wire[95:0] T345;
  wire[31:0] T346;
  wire[15:0] curRoute_dstPort;
  reg [15:0] dstPort;
  wire[15:0] T347;
  wire[15:0] T348;
  wire[15:0] T349;
  wire[15:0] T350;
  wire[7:0] T351;
  wire[15:0] curRoute_srcPort;
  reg [15:0] srcPort;
  wire[15:0] T352;
  wire[15:0] T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[63:0] T357;
  wire[31:0] curRoute_dstAddr;
  reg [31:0] dstAddr;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[23:0] T361;
  wire[31:0] curRoute_srcAddr;
  reg [31:0] srcAddr;
  wire[31:0] T362;
  wire[31:0] T363;
  wire[31:0] T364;
  wire[23:0] T365;
  wire T224;
  wire T225;
  reg [3:0] curTag;
  wire[3:0] T279;
  wire[3:0] T256;
  wire[3:0] T257;
  reg [3:0] resTag;
  wire[3:0] T366;
  reg [7:0] reqPktRoute_srcMac_1;
  wire[7:0] T367;
  wire[7:0] T368;
  reg [7:0] reqPktRoute_srcMac_2;
  wire[7:0] T369;
  wire[7:0] T370;
  reg [7:0] reqPktRoute_srcMac_3;
  wire[7:0] T371;
  wire[7:0] T372;
  reg [7:0] reqPktRoute_srcMac_4;
  wire[7:0] T373;
  wire[7:0] T374;
  reg [7:0] reqPktRoute_srcMac_5;
  wire[7:0] T375;
  wire[7:0] T376;
  reg [7:0] reqPktRoute_dstMac_0;
  wire[7:0] T377;
  wire[7:0] T378;
  reg [7:0] reqPktRoute_dstMac_1;
  wire[7:0] T379;
  wire[7:0] T380;
  reg [7:0] reqPktRoute_dstMac_2;
  wire[7:0] T381;
  wire[7:0] T382;
  reg [7:0] reqPktRoute_dstMac_3;
  wire[7:0] T383;
  wire[7:0] T384;
  reg [7:0] reqPktRoute_dstMac_4;
  wire[7:0] T385;
  wire[7:0] T386;
  reg [7:0] reqPktRoute_dstMac_5;
  wire[7:0] T387;
  wire[7:0] T388;
  reg [15:0] reqPktRoute_reqId;
  wire[15:0] T389;
  wire[15:0] T390;
  reg [15:0] reqPktRoute_dstPort;
  wire[15:0] T391;
  wire[15:0] T392;
  reg [15:0] reqPktRoute_srcPort;
  wire[15:0] T393;
  wire[15:0] T394;
  reg [31:0] reqPktRoute_dstAddr;
  wire[31:0] T395;
  wire[31:0] T396;
  reg [31:0] reqPktRoute_srcAddr;
  wire[31:0] T397;
  wire[31:0] T398;
  wire[15:0] T399;
  reg  sendDefer;
  wire T400;
  wire T401;
  wire T402;
  reg [15:0] reqPktLen;
  wire[15:0] T403;
  wire[15:0] T404;
  wire[7:0] T405;
  wire[7:0] T406;
  wire[7:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg  ignore;
  wire T417;
  wire T418;
  wire T419;
  wire rx_ready;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T0;
  wire T21;
  wire T22;
  wire T255;
  wire[7:0] T258;
  reg [15:0] keyLen;
  wire[15:0] T280;
  wire[15:0] T259;
  wire[15:0] T260;
  wire[15:0] T261;
  wire[15:0] T262;
  wire[7:0] T263;
  wire T264;
  wire mainWriter_io_stream_ready;
  wire[7:0] mainWriter_io_writeData;
  wire mainWriter_io_writeEn;
  wire[15:0] mainWriter_io_count;
  wire mainWriter_io_finished;
  wire mainBuffer_io_readData_valid;
  wire[7:0] mainBuffer_io_readData_data;
  wire mainBuffer_io_readData_last;
  wire mainBuffer_io_stream_ready;
  wire mainBuffer_io_skip_ready;
  wire mainBuffer_io_full;
  wire deferWriter_io_stream_ready;
  wire[7:0] deferWriter_io_writeData;
  wire deferWriter_io_writeEn;
  wire deferBuffer_io_readData_valid;
  wire[7:0] deferBuffer_io_readData_data;
  wire deferBuffer_io_readData_last;
  wire deferBuffer_io_stream_ready;
  wire deferBuffer_io_skip_ready;
  wire deferBuffer_io_full;
  wire streamSplit_io_in_ready;
  wire streamSplit_io_out_a_valid;
  wire[7:0] streamSplit_io_out_a_data;
  wire streamSplit_io_out_a_last;
  wire streamSplit_io_out_b_valid;
  wire[7:0] streamSplit_io_out_b_data;
  wire streamSplit_io_out_b_last;
  wire StreamArbiter_0_io_ins_1_ready;
  wire StreamArbiter_0_io_ins_0_ready;
  wire StreamArbiter_0_io_out_valid;
  wire[7:0] StreamArbiter_0_io_out_data;
  wire StreamArbiter_0_io_out_last;
  wire StreamArbiter_1_io_ins_1_ready;
  wire StreamArbiter_1_io_ins_0_ready;
  wire StreamArbiter_1_io_out_valid;
  wire[7:0] StreamArbiter_1_io_out_data;
  wire StreamArbiter_1_io_out_last;
  wire responder_io_temac_tx_valid;
  wire[7:0] responder_io_temac_tx_data;
  wire responder_io_temac_tx_last;
  wire responder_io_resultData_ready;
  wire responder_io_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    d_state = {1{$random}};
    resLen = {1{$random}};
    reqPktRoute_srcMac_0 = {1{$random}};
    srcMac_0 = {1{$random}};
    macIndex = {1{$random}};
    m_state = {1{$random}};
    etherTypeHigh = {1{$random}};
    lenOffset = {1{$random}};
    ipv6 = {1{$random}};
    headerLen = {1{$random}};
    pktLen = {1{$random}};
    srcMac_1 = {1{$random}};
    srcMac_2 = {1{$random}};
    srcMac_3 = {1{$random}};
    srcMac_4 = {1{$random}};
    srcMac_5 = {1{$random}};
    dstMac_0 = {1{$random}};
    dstMac_1 = {1{$random}};
    dstMac_2 = {1{$random}};
    dstMac_3 = {1{$random}};
    dstMac_4 = {1{$random}};
    dstMac_5 = {1{$random}};
    reqId = {1{$random}};
    dstPort = {1{$random}};
    srcPort = {1{$random}};
    dstAddr = {1{$random}};
    srcAddr = {1{$random}};
    curTag = {1{$random}};
    resTag = {1{$random}};
    reqPktRoute_srcMac_1 = {1{$random}};
    reqPktRoute_srcMac_2 = {1{$random}};
    reqPktRoute_srcMac_3 = {1{$random}};
    reqPktRoute_srcMac_4 = {1{$random}};
    reqPktRoute_srcMac_5 = {1{$random}};
    reqPktRoute_dstMac_0 = {1{$random}};
    reqPktRoute_dstMac_1 = {1{$random}};
    reqPktRoute_dstMac_2 = {1{$random}};
    reqPktRoute_dstMac_3 = {1{$random}};
    reqPktRoute_dstMac_4 = {1{$random}};
    reqPktRoute_dstMac_5 = {1{$random}};
    reqPktRoute_reqId = {1{$random}};
    reqPktRoute_dstPort = {1{$random}};
    reqPktRoute_srcPort = {1{$random}};
    reqPktRoute_dstAddr = {1{$random}};
    reqPktRoute_srcAddr = {1{$random}};
    sendDefer = {1{$random}};
    reqPktLen = {1{$random}};
    ignore = {1{$random}};
    keyLen = {1{$random}};
  end
`endif

  assign T281 = d_state == 3'h4;
  assign T265 = reset ? 3'h0 : T1;
  assign T1 = T19 ? 3'h0 : T2;
  assign T2 = T17 ? 3'h4 : T3;
  assign T3 = T15 ? 3'h0 : T4;
  assign T4 = T13 ? 3'h3 : T5;
  assign T5 = T9 ? 3'h2 : T6;
  assign T6 = T7 ? 3'h1 : d_state;
  assign T7 = T8 & io_resultInfo_valid;
  assign T8 = 3'h0 == d_state;
  assign T9 = T12 & T10;
  assign T10 = resLen == 8'h0;
  assign T266 = T11[3'h7:1'h0];
  assign T11 = T7 ? io_resultInfo_bits_len : T267;
  assign T267 = {11'h0, resLen};
  assign T12 = 3'h1 == d_state;
  assign T13 = T12 & T14;
  assign T14 = T10 ^ 1'h1;
  assign T15 = T16 & deferBuffer_io_stream_ready;
  assign T16 = 3'h2 == d_state;
  assign T17 = T18 & deferBuffer_io_skip_ready;
  assign T18 = 3'h3 == d_state;
  assign T19 = T20 & responder_io_ready;
  assign T20 = 3'h4 == d_state;
  assign T282 = T12 ? T283 : reqPktRoute_srcMac_0;
  assign T283 = T284[3'h7:1'h0];
  PacketFilter_getReqRoutes getReqRoutes (
    .CLK(clk),
    .W0A(curTag),
    .W0E(T224),
    .W0I(T286),
    .R1A(io_resultInfo_bits_tag),
    .R1E(T7),
    .R1O(T284)
  );
  assign T286 = T287;
  assign T287 = {T327, T288};
  assign T288 = {T310, T289};
  assign T289 = {T303, T290};
  assign T290 = {curRoute_srcMac_2, T291};
  assign T291 = {curRoute_srcMac_1, curRoute_srcMac_0};
  assign curRoute_srcMac_0 = srcMac_0;
  assign T292 = T293 ? mainWriter_io_writeData : srcMac_0;
  assign T293 = T89 & T294;
  assign T294 = T295[1'h0:1'h0];
  assign T295 = 1'h1 << T296;
  assign T296 = macIndex;
  assign T78 = T86 ? T85 : T79;
  assign T79 = T83 ? T82 : T80;
  assign T80 = T76 ? 3'h0 : T81;
  assign T81 = T72 ? 3'h0 : macIndex;
  assign T72 = T75 & T73;
  assign T73 = io_temac_rx_valid & T74;
  assign T74 = mainBuffer_io_full ^ 1'h1;
  assign T75 = 6'h0 == m_state;
  assign T268 = reset ? 6'h0 : T23;
  assign T23 = T253 ? 6'h0 : T24;
  assign T24 = T251 ? 6'h25 : T25;
  assign T25 = T248 ? 6'h0 : T26;
  assign T26 = T246 ? 6'ha : T27;
  assign T27 = T244 ? 6'ha : T28;
  assign T28 = T242 ? 6'h0 : T29;
  assign T29 = T240 ? 6'h23 : T30;
  assign T30 = T238 ? 6'h20 : T31;
  assign T31 = T235 ? 6'h22 : T32;
  assign T32 = T233 ? 6'h21 : T33;
  assign T33 = T231 ? 6'h20 : T34;
  assign T34 = T228 ? 6'h1f : T35;
  assign T35 = T226 ? 6'h1e : T36;
  assign T36 = T224 ? 6'h1d : T37;
  assign T37 = T222 ? 6'h1c : T38;
  assign T38 = T220 ? 6'h1b : T39;
  assign T39 = T218 ? 6'h9 : T40;
  assign T40 = T214 ? 6'h1a : T41;
  assign T41 = T212 ? 6'h9 : T42;
  assign T42 = T207 ? 6'h19 : T43;
  assign T43 = T204 ? 6'h9 : T44;
  assign T44 = T201 ? 6'h18 : T45;
  assign T45 = T199 ? 6'h17 : T46;
  assign T46 = T196 ? 6'h16 : T47;
  assign T47 = T185 ? 6'h9 : T48;
  assign T48 = T182 ? 6'h15 : T49;
  assign T49 = T180 ? 6'h14 : T50;
  assign T50 = T178 ? 6'h13 : T51;
  assign T51 = T176 ? 6'h12 : T52;
  assign T52 = T174 ? 6'h11 : T53;
  assign T53 = T171 ? 6'h10 : T54;
  assign T54 = T167 ? 6'hf : T55;
  assign T55 = T146 ? 6'h10 : T56;
  assign T56 = T142 ? 6'he : T57;
  assign T57 = T139 ? 6'hd : T58;
  assign T58 = T137 ? 6'h9 : T59;
  assign T59 = T132 ? 6'hc : T60;
  assign T60 = T130 ? 6'h8 : T61;
  assign T61 = T123 ? 6'h9 : T62;
  assign T62 = T118 ? 6'h7 : T63;
  assign T63 = T115 ? 6'hb : T64;
  assign T64 = T111 ? 6'h6 : T65;
  assign T65 = T106 ? 6'h6 : T66;
  assign T66 = T104 ? 6'h24 : T67;
  assign T67 = T96 ? 6'h5 : T68;
  assign T68 = T94 ? 6'h4 : T69;
  assign T69 = T93 ? 6'h3 : T70;
  assign T70 = T76 ? 6'h2 : T71;
  assign T71 = T72 ? 6'h1 : m_state;
  assign T93 = T89 & T88;
  assign T88 = macIndex == 3'h5;
  assign T94 = T95 & mainWriter_io_writeEn;
  assign T95 = 6'h3 == m_state;
  assign T96 = T102 & T97;
  assign T97 = T101 | T98;
  assign T98 = T99 == 16'h86dd;
  assign T99 = {etherTypeHigh, mainWriter_io_writeData};
  assign T100 = T94 ? mainWriter_io_writeData : etherTypeHigh;
  assign T101 = T99 == 16'h800;
  assign T102 = T103 & mainWriter_io_writeEn;
  assign T103 = 6'h4 == m_state;
  assign T104 = T102 & T105;
  assign T105 = T97 ^ 1'h1;
  assign T106 = T109 & T107;
  assign T107 = T108 == 4'h4;
  assign T108 = mainWriter_io_writeData[3'h7:3'h4];
  assign T109 = T110 & mainWriter_io_writeEn;
  assign T110 = 6'h5 == m_state;
  assign T111 = T109 & T112;
  assign T112 = T114 & T113;
  assign T113 = T108 == 4'h6;
  assign T114 = T107 ^ 1'h1;
  assign T115 = T109 & T116;
  assign T116 = T117 ^ 1'h1;
  assign T117 = T107 | T113;
  assign T118 = T122 & T119;
  assign T119 = mainWriter_io_count == lenOffset;
  assign T120 = T111 ? 16'h13 : T121;
  assign T121 = T106 ? 16'h11 : lenOffset;
  assign T122 = 6'h6 == m_state;
  assign T123 = T128 & T124;
  assign T124 = ipv6 | T125;
  assign T125 = io_readready ^ 1'h1;
  assign T126 = T111 ? 1'h1 : T127;
  assign T127 = T106 ? 1'h0 : ipv6;
  assign T128 = T129 & mainWriter_io_writeEn;
  assign T129 = 6'h7 == m_state;
  assign T130 = T128 & T131;
  assign T131 = T124 ^ 1'h1;
  assign T132 = T134 & T133;
  assign T133 = mainWriter_io_writeData == 8'h11;
  assign T134 = T136 & T135;
  assign T135 = mainWriter_io_count == 16'h18;
  assign T136 = 6'h8 == m_state;
  assign T137 = T134 & T138;
  assign T138 = T133 ^ 1'h1;
  assign T139 = T141 & T140;
  assign T140 = mainWriter_io_count == 16'h1a;
  assign T141 = 6'hc == m_state;
  assign T142 = T144 & T143;
  assign T143 = mainWriter_io_count == 16'h1e;
  assign T144 = T145 & mainWriter_io_writeEn;
  assign T145 = 6'hd == m_state;
  assign T146 = T165 & T147;
  assign T147 = mainWriter_io_count == T269;
  assign T269 = {8'h0, headerLen};
  assign T270 = reset ? 8'h0 : T148;
  assign T148 = T224 ? T164 : T149;
  assign T149 = T201 ? T163 : T150;
  assign T150 = T182 ? T162 : T151;
  assign T151 = T171 ? T161 : T152;
  assign T152 = T146 ? T160 : T153;
  assign T153 = T111 ? T159 : T154;
  assign T154 = T106 ? T156 : T155;
  assign T155 = T72 ? 8'he : headerLen;
  assign T156 = headerLen + T271;
  assign T271 = {2'h0, T157};
  assign T157 = {T158, 2'h0};
  assign T158 = mainWriter_io_writeData[2'h3:1'h0];
  assign T159 = headerLen + 8'h28;
  assign T160 = headerLen + 8'h8;
  assign T161 = headerLen + 8'h8;
  assign T162 = headerLen + 8'h8;
  assign T163 = headerLen + 8'h18;
  assign T164 = headerLen + mainWriter_io_writeData;
  assign T165 = T166 & mainWriter_io_writeEn;
  assign T166 = 6'he == m_state;
  assign T167 = T165 & T168;
  assign T168 = T170 & T169;
  assign T169 = mainWriter_io_count == 16'h22;
  assign T170 = T147 ^ 1'h1;
  assign T171 = T173 & T172;
  assign T172 = mainWriter_io_count == T272;
  assign T272 = {8'h0, headerLen};
  assign T173 = 6'hf == m_state;
  assign T174 = T175 & mainWriter_io_writeEn;
  assign T175 = 6'h10 == m_state;
  assign T176 = T177 & mainWriter_io_writeEn;
  assign T177 = 6'h11 == m_state;
  assign T178 = T179 & mainWriter_io_writeEn;
  assign T179 = 6'h12 == m_state;
  assign T180 = T181 & mainWriter_io_writeEn;
  assign T181 = 6'h13 == m_state;
  assign T182 = T184 & T183;
  assign T183 = mainWriter_io_count == T273;
  assign T273 = {8'h0, headerLen};
  assign T184 = 6'h14 == m_state;
  assign T185 = T195 & T186;
  assign T186 = pktLen <= T274;
  assign T274 = {8'h0, headerLen};
  assign T275 = reset ? 16'h0 : T187;
  assign T187 = T251 ? mainWriter_io_count : T188;
  assign T188 = T128 ? T192 : T189;
  assign T189 = T118 ? T191 : T190;
  assign T190 = T115 ? 16'h10 : pktLen;
  assign T191 = {mainWriter_io_writeData, 8'h0};
  assign T192 = T193 + 16'he;
  assign T193 = {T194, mainWriter_io_writeData};
  assign T194 = pktLen[4'hf:4'h8];
  assign T195 = 6'h15 == m_state;
  assign T196 = T195 & T197;
  assign T197 = T198 & mainWriter_io_writeEn;
  assign T198 = T186 ^ 1'h1;
  assign T199 = T200 & mainWriter_io_writeEn;
  assign T200 = 6'h16 == m_state;
  assign T201 = T203 & T202;
  assign T202 = mainWriter_io_count == T276;
  assign T276 = {8'h0, headerLen};
  assign T203 = 6'h17 == m_state;
  assign T204 = T206 & T205;
  assign T205 = pktLen <= T277;
  assign T277 = {8'h0, headerLen};
  assign T206 = 6'h18 == m_state;
  assign T207 = T209 & T208;
  assign T208 = mainWriter_io_writeData == 8'h80;
  assign T209 = T206 & T210;
  assign T210 = T211 & mainWriter_io_writeEn;
  assign T211 = T205 ^ 1'h1;
  assign T212 = T209 & T213;
  assign T213 = T208 ^ 1'h1;
  assign T214 = T216 & T215;
  assign T215 = mainWriter_io_writeData == 8'h0;
  assign T216 = T217 & mainWriter_io_writeEn;
  assign T217 = 6'h19 == m_state;
  assign T218 = T216 & T219;
  assign T219 = T215 ^ 1'h1;
  assign T220 = T221 & mainWriter_io_writeEn;
  assign T221 = 6'h1a == m_state;
  assign T222 = T223 & mainWriter_io_writeEn;
  assign T223 = 6'h1b == m_state;
  assign T226 = T227 & io_keyInfo_ready;
  assign T227 = 6'h1d == m_state;
  assign T228 = T230 & T229;
  assign T229 = mainWriter_io_count == T278;
  assign T278 = {8'h0, headerLen};
  assign T230 = 6'h1e == m_state;
  assign T231 = T232 & mainBuffer_io_stream_ready;
  assign T232 = 6'h1f == m_state;
  assign T233 = T234 & io_keyData_ready;
  assign T234 = 6'h20 == m_state;
  assign T235 = T236 & io_temac_rx_last;
  assign T236 = T237 & io_temac_rx_valid;
  assign T237 = 6'h21 == m_state;
  assign T238 = T236 & T239;
  assign T239 = io_temac_rx_last ^ 1'h1;
  assign T240 = T241 & io_keyData_ready;
  assign T241 = 6'h22 == m_state;
  assign T242 = T243 & mainBuffer_io_stream_ready;
  assign T243 = 6'h23 == m_state;
  assign T244 = T245 & mainBuffer_io_stream_ready;
  assign T245 = 6'h9 == m_state;
  assign T246 = T247 & mainBuffer_io_skip_ready;
  assign T247 = 6'hb == m_state;
  assign T248 = T250 & T249;
  assign T249 = io_temac_rx_valid & io_temac_rx_last;
  assign T250 = 6'ha == m_state;
  assign T251 = T252 & mainWriter_io_finished;
  assign T252 = 6'h24 == m_state;
  assign T253 = T254 & mainBuffer_io_stream_ready;
  assign T254 = 6'h25 == m_state;
  assign T76 = T91 & T77;
  assign T77 = macIndex == 3'h5;
  assign T91 = T92 & mainWriter_io_writeEn;
  assign T92 = 6'h1 == m_state;
  assign T82 = macIndex + 3'h1;
  assign T83 = T91 & T84;
  assign T84 = T77 ^ 1'h1;
  assign T85 = macIndex + 3'h1;
  assign T86 = T89 & T87;
  assign T87 = T88 ^ 1'h1;
  assign T89 = T90 & mainWriter_io_writeEn;
  assign T90 = 6'h2 == m_state;
  assign curRoute_srcMac_1 = srcMac_1;
  assign T297 = T298 ? mainWriter_io_writeData : srcMac_1;
  assign T298 = T89 & T299;
  assign T299 = T295[1'h1:1'h1];
  assign curRoute_srcMac_2 = srcMac_2;
  assign T300 = T301 ? mainWriter_io_writeData : srcMac_2;
  assign T301 = T89 & T302;
  assign T302 = T295[2'h2:2'h2];
  assign T303 = {curRoute_srcMac_4, curRoute_srcMac_3};
  assign curRoute_srcMac_3 = srcMac_3;
  assign T304 = T305 ? mainWriter_io_writeData : srcMac_3;
  assign T305 = T89 & T306;
  assign T306 = T295[2'h3:2'h3];
  assign curRoute_srcMac_4 = srcMac_4;
  assign T307 = T308 ? mainWriter_io_writeData : srcMac_4;
  assign T308 = T89 & T309;
  assign T309 = T295[3'h4:3'h4];
  assign T310 = {T320, T311};
  assign T311 = {curRoute_dstMac_0, curRoute_srcMac_5};
  assign curRoute_srcMac_5 = srcMac_5;
  assign T312 = T313 ? mainWriter_io_writeData : srcMac_5;
  assign T313 = T89 & T314;
  assign T314 = T295[3'h5:3'h5];
  assign curRoute_dstMac_0 = dstMac_0;
  assign T315 = T316 ? mainWriter_io_writeData : dstMac_0;
  assign T316 = T91 & T317;
  assign T317 = T318[1'h0:1'h0];
  assign T318 = 1'h1 << T319;
  assign T319 = macIndex;
  assign T320 = {curRoute_dstMac_2, curRoute_dstMac_1};
  assign curRoute_dstMac_1 = dstMac_1;
  assign T321 = T322 ? mainWriter_io_writeData : dstMac_1;
  assign T322 = T91 & T323;
  assign T323 = T318[1'h1:1'h1];
  assign curRoute_dstMac_2 = dstMac_2;
  assign T324 = T325 ? mainWriter_io_writeData : dstMac_2;
  assign T325 = T91 & T326;
  assign T326 = T318[2'h2:2'h2];
  assign T327 = {T345, T328};
  assign T328 = {T336, T329};
  assign T329 = {curRoute_dstMac_4, curRoute_dstMac_3};
  assign curRoute_dstMac_3 = dstMac_3;
  assign T330 = T331 ? mainWriter_io_writeData : dstMac_3;
  assign T331 = T91 & T332;
  assign T332 = T318[2'h3:2'h3];
  assign curRoute_dstMac_4 = dstMac_4;
  assign T333 = T334 ? mainWriter_io_writeData : dstMac_4;
  assign T334 = T91 & T335;
  assign T335 = T318[3'h4:3'h4];
  assign T336 = {curRoute_reqId, curRoute_dstMac_5};
  assign curRoute_dstMac_5 = dstMac_5;
  assign T337 = T338 ? mainWriter_io_writeData : dstMac_5;
  assign T338 = T91 & T339;
  assign T339 = T318[3'h5:3'h5];
  assign curRoute_reqId = reqId;
  assign T340 = T199 ? T343 : T341;
  assign T341 = T196 ? T342 : reqId;
  assign T342 = {mainWriter_io_writeData, 8'h0};
  assign T343 = {T344, mainWriter_io_writeData};
  assign T344 = reqId[4'hf:4'h8];
  assign T345 = {T357, T346};
  assign T346 = {curRoute_srcPort, curRoute_dstPort};
  assign curRoute_dstPort = dstPort;
  assign T347 = T180 ? T350 : T348;
  assign T348 = T178 ? T349 : dstPort;
  assign T349 = {mainWriter_io_writeData, 8'h0};
  assign T350 = {T351, mainWriter_io_writeData};
  assign T351 = dstPort[4'hf:4'h8];
  assign curRoute_srcPort = srcPort;
  assign T352 = T176 ? T355 : T353;
  assign T353 = T174 ? T354 : srcPort;
  assign T354 = {mainWriter_io_writeData, 8'h0};
  assign T355 = {T356, mainWriter_io_writeData};
  assign T356 = srcPort[4'hf:4'h8];
  assign T357 = {curRoute_srcAddr, curRoute_dstAddr};
  assign curRoute_dstAddr = dstAddr;
  assign T358 = T165 ? T360 : T359;
  assign T359 = T142 ? 32'h0 : dstAddr;
  assign T360 = {T361, mainWriter_io_writeData};
  assign T361 = dstAddr[5'h17:1'h0];
  assign curRoute_srcAddr = srcAddr;
  assign T362 = T144 ? T364 : T363;
  assign T363 = T139 ? 32'h0 : srcAddr;
  assign T364 = {T365, mainWriter_io_writeData};
  assign T365 = srcAddr[5'h17:1'h0];
  assign T224 = T225 & mainWriter_io_writeEn;
  assign T225 = 6'h1c == m_state;
  assign T279 = reset ? 4'h0 : T256;
  assign T256 = T226 ? T257 : curTag;
  assign T257 = curTag + 4'h1;
  assign T366 = T7 ? io_resultInfo_bits_tag : resTag;
  assign T367 = T12 ? T368 : reqPktRoute_srcMac_1;
  assign T368 = T284[4'hf:4'h8];
  assign T369 = T12 ? T370 : reqPktRoute_srcMac_2;
  assign T370 = T284[5'h17:5'h10];
  assign T371 = T12 ? T372 : reqPktRoute_srcMac_3;
  assign T372 = T284[5'h1f:5'h18];
  assign T373 = T12 ? T374 : reqPktRoute_srcMac_4;
  assign T374 = T284[6'h27:6'h20];
  assign T375 = T12 ? T376 : reqPktRoute_srcMac_5;
  assign T376 = T284[6'h2f:6'h28];
  assign T377 = T12 ? T378 : reqPktRoute_dstMac_0;
  assign T378 = T284[6'h37:6'h30];
  assign T379 = T12 ? T380 : reqPktRoute_dstMac_1;
  assign T380 = T284[6'h3f:6'h38];
  assign T381 = T12 ? T382 : reqPktRoute_dstMac_2;
  assign T382 = T284[7'h47:7'h40];
  assign T383 = T12 ? T384 : reqPktRoute_dstMac_3;
  assign T384 = T284[7'h4f:7'h48];
  assign T385 = T12 ? T386 : reqPktRoute_dstMac_4;
  assign T386 = T284[7'h57:7'h50];
  assign T387 = T12 ? T388 : reqPktRoute_dstMac_5;
  assign T388 = T284[7'h5f:7'h58];
  assign T389 = T12 ? T390 : reqPktRoute_reqId;
  assign T390 = T284[7'h6f:7'h60];
  assign T391 = T12 ? T392 : reqPktRoute_dstPort;
  assign T392 = T284[7'h7f:7'h70];
  assign T393 = T12 ? T394 : reqPktRoute_srcPort;
  assign T394 = T284[8'h8f:8'h80];
  assign T395 = T12 ? T396 : reqPktRoute_dstAddr;
  assign T396 = T284[8'haf:8'h90];
  assign T397 = T12 ? T398 : reqPktRoute_srcAddr;
  assign T398 = T284[8'hcf:8'hb0];
  assign T399 = {8'h0, resLen};
  assign T400 = reset ? 1'h0 : T401;
  assign T401 = T242 ? 1'h0 : T402;
  assign T402 = T228 ? 1'h1 : sendDefer;
  assign T403 = T12 ? T404 : reqPktLen;
  assign T404 = {8'h0, T405};
  PacketFilter_getReqLens getReqLens (
    .CLK(clk),
    .W0A(curTag),
    .W0E(T226),
    .W0I(T407),
    .R1A(io_resultInfo_bits_tag),
    .R1E(T7),
    .R1O(T405)
  );
  assign T407 = pktLen[3'h7:1'h0];
  assign T408 = d_state == 3'h3;
  assign T409 = d_state == 3'h2;
  assign T410 = deferBuffer_io_full ^ 1'h1;
  assign T411 = m_state == 6'hb;
  assign T412 = T414 | T413;
  assign T413 = m_state == 6'h25;
  assign T414 = T416 | T415;
  assign T415 = m_state == 6'h1f;
  assign T416 = m_state == 6'h9;
  assign T417 = reset ? 1'h0 : T418;
  assign T418 = T248 ? 1'h0 : T419;
  assign T419 = T115 ? 1'h1 : ignore;
  assign rx_ready = T421 & T420;
  assign T420 = mainBuffer_io_full ^ 1'h1;
  assign T421 = T423 & T422;
  assign T422 = m_state != 6'h25;
  assign T423 = T425 & T424;
  assign T424 = m_state != 6'h23;
  assign T425 = T427 & T426;
  assign T426 = m_state != 6'h22;
  assign T427 = T429 & T428;
  assign T428 = m_state != 6'h20;
  assign T429 = T431 & T430;
  assign T430 = m_state != 6'h1f;
  assign T431 = T433 & T432;
  assign T432 = m_state != 6'h1d;
  assign T433 = T435 & T434;
  assign T434 = m_state != 6'hb;
  assign T435 = m_state != 6'h9;
  assign io_resultData_ready = responder_io_resultData_ready;
  assign io_resultInfo_ready = T0;
  assign T0 = d_state == 3'h0;
  assign io_keyData_bits = mainWriter_io_writeData;
  assign io_keyData_valid = T21;
  assign T21 = T255 | T22;
  assign T22 = m_state == 6'h22;
  assign T255 = m_state == 6'h20;
  assign io_keyInfo_bits_tag = curTag;
  assign io_keyInfo_bits_len = T258;
  assign T258 = keyLen[3'h7:1'h0];
  assign T280 = reset ? 16'h0 : T259;
  assign T259 = T222 ? T262 : T260;
  assign T260 = T220 ? T261 : keyLen;
  assign T261 = {mainWriter_io_writeData, 8'h0};
  assign T262 = {T263, mainWriter_io_writeData};
  assign T263 = keyLen[4'hf:4'h8];
  assign io_keyInfo_valid = T264;
  assign T264 = m_state == 6'h1d;
  assign io_core_tx_ready = StreamArbiter_1_io_ins_0_ready;
  assign io_temac_tx_last = StreamArbiter_1_io_out_last;
  assign io_temac_tx_data = StreamArbiter_1_io_out_data;
  assign io_temac_tx_valid = StreamArbiter_1_io_out_valid;
  assign io_core_rx_last = StreamArbiter_0_io_out_last;
  assign io_core_rx_data = StreamArbiter_0_io_out_data;
  assign io_core_rx_valid = StreamArbiter_0_io_out_valid;
  assign io_temac_rx_ready = mainWriter_io_stream_ready;
  StreamWriter mainWriter(.clk(clk), .reset(reset),
       .io_stream_ready( mainWriter_io_stream_ready ),
       .io_stream_valid( io_temac_rx_valid ),
       .io_stream_data( io_temac_rx_data ),
       .io_stream_last( io_temac_rx_last ),
       .io_writeData( mainWriter_io_writeData ),
       .io_writeEn( mainWriter_io_writeEn ),
       .io_enable( rx_ready ),
       .io_ignore( ignore ),
       .io_count( mainWriter_io_count ),
       .io_finished( mainWriter_io_finished )
  );
  PacketBuffer mainBuffer(.clk(clk), .reset(reset),
       .io_readData_ready( streamSplit_io_in_ready ),
       .io_readData_valid( mainBuffer_io_readData_valid ),
       .io_readData_data( mainBuffer_io_readData_data ),
       .io_readData_last( mainBuffer_io_readData_last ),
       .io_stream_ready( mainBuffer_io_stream_ready ),
       .io_stream_valid( T412 ),
       .io_stream_bits( pktLen ),
       .io_skip_ready( mainBuffer_io_skip_ready ),
       .io_skip_valid( T411 ),
       .io_skip_bits( pktLen ),
       .io_writeData( mainWriter_io_writeData ),
       .io_writeEn( mainWriter_io_writeEn ),
       //.io_empty(  )
       .io_full( mainBuffer_io_full )
  );
  StreamWriter deferWriter(.clk(clk), .reset(reset),
       .io_stream_ready( deferWriter_io_stream_ready ),
       .io_stream_valid( streamSplit_io_out_b_valid ),
       .io_stream_data( streamSplit_io_out_b_data ),
       .io_stream_last( streamSplit_io_out_b_last ),
       .io_writeData( deferWriter_io_writeData ),
       .io_writeEn( deferWriter_io_writeEn ),
       .io_enable( T410 ),
       .io_ignore( 1'h0 )
       //.io_count(  )
       //.io_finished(  )
  );
  PacketBuffer deferBuffer(.clk(clk), .reset(reset),
       .io_readData_ready( StreamArbiter_0_io_ins_1_ready ),
       .io_readData_valid( deferBuffer_io_readData_valid ),
       .io_readData_data( deferBuffer_io_readData_data ),
       .io_readData_last( deferBuffer_io_readData_last ),
       .io_stream_ready( deferBuffer_io_stream_ready ),
       .io_stream_valid( T409 ),
       .io_stream_bits( reqPktLen ),
       .io_skip_ready( deferBuffer_io_skip_ready ),
       .io_skip_valid( T408 ),
       .io_skip_bits( reqPktLen ),
       .io_writeData( deferWriter_io_writeData ),
       .io_writeEn( deferWriter_io_writeEn ),
       //.io_empty(  )
       .io_full( deferBuffer_io_full )
  );
  StreamSplit streamSplit(
       .io_in_ready( streamSplit_io_in_ready ),
       .io_in_valid( mainBuffer_io_readData_valid ),
       .io_in_data( mainBuffer_io_readData_data ),
       .io_in_last( mainBuffer_io_readData_last ),
       .io_out_a_ready( StreamArbiter_0_io_ins_0_ready ),
       .io_out_a_valid( streamSplit_io_out_a_valid ),
       .io_out_a_data( streamSplit_io_out_a_data ),
       .io_out_a_last( streamSplit_io_out_a_last ),
       .io_out_b_ready( deferWriter_io_stream_ready ),
       .io_out_b_valid( streamSplit_io_out_b_valid ),
       .io_out_b_data( streamSplit_io_out_b_data ),
       .io_out_b_last( streamSplit_io_out_b_last ),
       .io_sel( sendDefer )
  );
  StreamArbiter StreamArbiter_0(.clk(clk), .reset(reset),
       .io_ins_1_ready( StreamArbiter_0_io_ins_1_ready ),
       .io_ins_1_valid( deferBuffer_io_readData_valid ),
       .io_ins_1_data( deferBuffer_io_readData_data ),
       .io_ins_1_last( deferBuffer_io_readData_last ),
       .io_ins_0_ready( StreamArbiter_0_io_ins_0_ready ),
       .io_ins_0_valid( streamSplit_io_out_a_valid ),
       .io_ins_0_data( streamSplit_io_out_a_data ),
       .io_ins_0_last( streamSplit_io_out_a_last ),
       .io_out_ready( io_core_rx_ready ),
       .io_out_valid( StreamArbiter_0_io_out_valid ),
       .io_out_data( StreamArbiter_0_io_out_data ),
       .io_out_last( StreamArbiter_0_io_out_last )
  );
  Responder responder(.clk(clk), .reset(reset),
       .io_temac_tx_ready( StreamArbiter_1_io_ins_1_ready ),
       .io_temac_tx_valid( responder_io_temac_tx_valid ),
       .io_temac_tx_data( responder_io_temac_tx_data ),
       .io_temac_tx_last( responder_io_temac_tx_last ),
       .io_resultData_ready( responder_io_resultData_ready ),
       .io_resultData_valid( io_resultData_valid ),
       .io_resultData_bits( io_resultData_bits ),
       .io_resLen( T399 ),
       .io_pktRoute_srcAddr( reqPktRoute_srcAddr ),
       .io_pktRoute_dstAddr( reqPktRoute_dstAddr ),
       .io_pktRoute_srcPort( reqPktRoute_srcPort ),
       .io_pktRoute_dstPort( reqPktRoute_dstPort ),
       .io_pktRoute_reqId( reqPktRoute_reqId ),
       .io_pktRoute_dstMac_5( reqPktRoute_dstMac_5 ),
       .io_pktRoute_dstMac_4( reqPktRoute_dstMac_4 ),
       .io_pktRoute_dstMac_3( reqPktRoute_dstMac_3 ),
       .io_pktRoute_dstMac_2( reqPktRoute_dstMac_2 ),
       .io_pktRoute_dstMac_1( reqPktRoute_dstMac_1 ),
       .io_pktRoute_dstMac_0( reqPktRoute_dstMac_0 ),
       .io_pktRoute_srcMac_5( reqPktRoute_srcMac_5 ),
       .io_pktRoute_srcMac_4( reqPktRoute_srcMac_4 ),
       .io_pktRoute_srcMac_3( reqPktRoute_srcMac_3 ),
       .io_pktRoute_srcMac_2( reqPktRoute_srcMac_2 ),
       .io_pktRoute_srcMac_1( reqPktRoute_srcMac_1 ),
       .io_pktRoute_srcMac_0( reqPktRoute_srcMac_0 ),
       .io_start( T281 ),
       .io_ready( responder_io_ready )
  );
  StreamArbiter StreamArbiter_1(.clk(clk), .reset(reset),
       .io_ins_1_ready( StreamArbiter_1_io_ins_1_ready ),
       .io_ins_1_valid( responder_io_temac_tx_valid ),
       .io_ins_1_data( responder_io_temac_tx_data ),
       .io_ins_1_last( responder_io_temac_tx_last ),
       .io_ins_0_ready( StreamArbiter_1_io_ins_0_ready ),
       .io_ins_0_valid( io_core_tx_valid ),
       .io_ins_0_data( io_core_tx_data ),
       .io_ins_0_last( io_core_tx_last ),
       .io_out_ready( io_temac_tx_ready ),
       .io_out_valid( StreamArbiter_1_io_out_valid ),
       .io_out_data( StreamArbiter_1_io_out_data ),
       .io_out_last( StreamArbiter_1_io_out_last )
  );

  always @(posedge clk) begin
    if(reset) begin
      d_state <= 3'h0;
    end else if(T19) begin
      d_state <= 3'h0;
    end else if(T17) begin
      d_state <= 3'h4;
    end else if(T15) begin
      d_state <= 3'h0;
    end else if(T13) begin
      d_state <= 3'h3;
    end else if(T9) begin
      d_state <= 3'h2;
    end else if(T7) begin
      d_state <= 3'h1;
    end
    resLen <= T266;
    if(T12) begin
      reqPktRoute_srcMac_0 <= T283;
    end
    if(T293) begin
      srcMac_0 <= mainWriter_io_writeData;
    end
    if(T86) begin
      macIndex <= T85;
    end else if(T83) begin
      macIndex <= T82;
    end else if(T76) begin
      macIndex <= 3'h0;
    end else if(T72) begin
      macIndex <= 3'h0;
    end
    if(reset) begin
      m_state <= 6'h0;
    end else if(T253) begin
      m_state <= 6'h0;
    end else if(T251) begin
      m_state <= 6'h25;
    end else if(T248) begin
      m_state <= 6'h0;
    end else if(T246) begin
      m_state <= 6'ha;
    end else if(T244) begin
      m_state <= 6'ha;
    end else if(T242) begin
      m_state <= 6'h0;
    end else if(T240) begin
      m_state <= 6'h23;
    end else if(T238) begin
      m_state <= 6'h20;
    end else if(T235) begin
      m_state <= 6'h22;
    end else if(T233) begin
      m_state <= 6'h21;
    end else if(T231) begin
      m_state <= 6'h20;
    end else if(T228) begin
      m_state <= 6'h1f;
    end else if(T226) begin
      m_state <= 6'h1e;
    end else if(T224) begin
      m_state <= 6'h1d;
    end else if(T222) begin
      m_state <= 6'h1c;
    end else if(T220) begin
      m_state <= 6'h1b;
    end else if(T218) begin
      m_state <= 6'h9;
    end else if(T214) begin
      m_state <= 6'h1a;
    end else if(T212) begin
      m_state <= 6'h9;
    end else if(T207) begin
      m_state <= 6'h19;
    end else if(T204) begin
      m_state <= 6'h9;
    end else if(T201) begin
      m_state <= 6'h18;
    end else if(T199) begin
      m_state <= 6'h17;
    end else if(T196) begin
      m_state <= 6'h16;
    end else if(T185) begin
      m_state <= 6'h9;
    end else if(T182) begin
      m_state <= 6'h15;
    end else if(T180) begin
      m_state <= 6'h14;
    end else if(T178) begin
      m_state <= 6'h13;
    end else if(T176) begin
      m_state <= 6'h12;
    end else if(T174) begin
      m_state <= 6'h11;
    end else if(T171) begin
      m_state <= 6'h10;
    end else if(T167) begin
      m_state <= 6'hf;
    end else if(T146) begin
      m_state <= 6'h10;
    end else if(T142) begin
      m_state <= 6'he;
    end else if(T139) begin
      m_state <= 6'hd;
    end else if(T137) begin
      m_state <= 6'h9;
    end else if(T132) begin
      m_state <= 6'hc;
    end else if(T130) begin
      m_state <= 6'h8;
    end else if(T123) begin
      m_state <= 6'h9;
    end else if(T118) begin
      m_state <= 6'h7;
    end else if(T115) begin
      m_state <= 6'hb;
    end else if(T111) begin
      m_state <= 6'h6;
    end else if(T106) begin
      m_state <= 6'h6;
    end else if(T104) begin
      m_state <= 6'h24;
    end else if(T96) begin
      m_state <= 6'h5;
    end else if(T94) begin
      m_state <= 6'h4;
    end else if(T93) begin
      m_state <= 6'h3;
    end else if(T76) begin
      m_state <= 6'h2;
    end else if(T72) begin
      m_state <= 6'h1;
    end
    if(T94) begin
      etherTypeHigh <= mainWriter_io_writeData;
    end
    if(T111) begin
      lenOffset <= 16'h13;
    end else if(T106) begin
      lenOffset <= 16'h11;
    end
    if(T111) begin
      ipv6 <= 1'h1;
    end else if(T106) begin
      ipv6 <= 1'h0;
    end
    if(reset) begin
      headerLen <= 8'h0;
    end else if(T224) begin
      headerLen <= T164;
    end else if(T201) begin
      headerLen <= T163;
    end else if(T182) begin
      headerLen <= T162;
    end else if(T171) begin
      headerLen <= T161;
    end else if(T146) begin
      headerLen <= T160;
    end else if(T111) begin
      headerLen <= T159;
    end else if(T106) begin
      headerLen <= T156;
    end else if(T72) begin
      headerLen <= 8'he;
    end
    if(reset) begin
      pktLen <= 16'h0;
    end else if(T251) begin
      pktLen <= mainWriter_io_count;
    end else if(T128) begin
      pktLen <= T192;
    end else if(T118) begin
      pktLen <= T191;
    end else if(T115) begin
      pktLen <= 16'h10;
    end
    if(T298) begin
      srcMac_1 <= mainWriter_io_writeData;
    end
    if(T301) begin
      srcMac_2 <= mainWriter_io_writeData;
    end
    if(T305) begin
      srcMac_3 <= mainWriter_io_writeData;
    end
    if(T308) begin
      srcMac_4 <= mainWriter_io_writeData;
    end
    if(T313) begin
      srcMac_5 <= mainWriter_io_writeData;
    end
    if(T316) begin
      dstMac_0 <= mainWriter_io_writeData;
    end
    if(T322) begin
      dstMac_1 <= mainWriter_io_writeData;
    end
    if(T325) begin
      dstMac_2 <= mainWriter_io_writeData;
    end
    if(T331) begin
      dstMac_3 <= mainWriter_io_writeData;
    end
    if(T334) begin
      dstMac_4 <= mainWriter_io_writeData;
    end
    if(T338) begin
      dstMac_5 <= mainWriter_io_writeData;
    end
    if(T199) begin
      reqId <= T343;
    end else if(T196) begin
      reqId <= T342;
    end
    if(T180) begin
      dstPort <= T350;
    end else if(T178) begin
      dstPort <= T349;
    end
    if(T176) begin
      srcPort <= T355;
    end else if(T174) begin
      srcPort <= T354;
    end
    if(T165) begin
      dstAddr <= T360;
    end else if(T142) begin
      dstAddr <= 32'h0;
    end
    if(T144) begin
      srcAddr <= T364;
    end else if(T139) begin
      srcAddr <= 32'h0;
    end
    if(reset) begin
      curTag <= 4'h0;
    end else if(T226) begin
      curTag <= T257;
    end
    if(T7) begin
      resTag <= io_resultInfo_bits_tag;
    end
    if(T12) begin
      reqPktRoute_srcMac_1 <= T368;
    end
    if(T12) begin
      reqPktRoute_srcMac_2 <= T370;
    end
    if(T12) begin
      reqPktRoute_srcMac_3 <= T372;
    end
    if(T12) begin
      reqPktRoute_srcMac_4 <= T374;
    end
    if(T12) begin
      reqPktRoute_srcMac_5 <= T376;
    end
    if(T12) begin
      reqPktRoute_dstMac_0 <= T378;
    end
    if(T12) begin
      reqPktRoute_dstMac_1 <= T380;
    end
    if(T12) begin
      reqPktRoute_dstMac_2 <= T382;
    end
    if(T12) begin
      reqPktRoute_dstMac_3 <= T384;
    end
    if(T12) begin
      reqPktRoute_dstMac_4 <= T386;
    end
    if(T12) begin
      reqPktRoute_dstMac_5 <= T388;
    end
    if(T12) begin
      reqPktRoute_reqId <= T390;
    end
    if(T12) begin
      reqPktRoute_dstPort <= T392;
    end
    if(T12) begin
      reqPktRoute_srcPort <= T394;
    end
    if(T12) begin
      reqPktRoute_dstAddr <= T396;
    end
    if(T12) begin
      reqPktRoute_srcAddr <= T398;
    end
    if(reset) begin
      sendDefer <= 1'h0;
    end else if(T242) begin
      sendDefer <= 1'h0;
    end else if(T228) begin
      sendDefer <= 1'h1;
    end
    if(T12) begin
      reqPktLen <= T404;
    end
    if(reset) begin
      ignore <= 1'h0;
    end else if(T248) begin
      ignore <= 1'h0;
    end else if(T115) begin
      ignore <= 1'h1;
    end
    if(reset) begin
      keyLen <= 16'h0;
    end else if(T222) begin
      keyLen <= T262;
    end else if(T220) begin
      keyLen <= T261;
    end
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    input  io_mem_backup_en,
    output io_in_mem_ready,
    input  io_in_mem_valid,
    input  io_out_mem_ready,
    output io_out_mem_valid,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready,
    output io_temac_sfp_tx_disable,
    output io_debug_keyLen_valid,
    output[15:0] io_debug_keyLen_bits,
    output io_debug_keyData_valid,
    output[7:0] io_debug_keyData_bits,
    output io_debug_resultLen_valid,
    output[15:0] io_debug_resultLen_bits,
    output io_debug_resultData_valid,
    output[7:0] io_debug_resultData_bits,
    output io_debug_readready,
    output io_debug_rocc_inst_ready,
    output io_debug_rocc_inst_valid,
    output[6:0] io_debug_rocc_inst_bits_inst_funct,
    output[4:0] io_debug_rocc_inst_bits_inst_rs2,
    output[4:0] io_debug_rocc_inst_bits_inst_rs1,
    output io_debug_rocc_inst_bits_inst_xd,
    output io_debug_rocc_inst_bits_inst_xs1,
    output io_debug_rocc_inst_bits_inst_xs2,
    output[4:0] io_debug_rocc_inst_bits_inst_rd,
    output[6:0] io_debug_rocc_inst_bits_inst_opcode,
    output[63:0] io_debug_rocc_inst_bits_rs1,
    output[63:0] io_debug_rocc_inst_bits_rs2
);

  wire resetSigs_0;
  wire[4:0] T2;
  wire[42:0] T3;
  wire[43:0] T4;
  reg  R5;
  reg  R6;
  wire[15:0] T0;
  wire[15:0] T1;
  wire Queue_0_io_enq_ready;
  wire Queue_0_io_deq_valid;
  wire Queue_0_io_deq_bits_rw;
  wire[4:0] Queue_0_io_deq_bits_addr;
  wire[63:0] Queue_0_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire Queue_2_io_deq_bits;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire Queue_3_io_deq_bits;
  wire PacketFilter_io_temac_rx_ready;
  wire PacketFilter_io_core_rx_valid;
  wire[7:0] PacketFilter_io_core_rx_data;
  wire PacketFilter_io_core_rx_last;
  wire PacketFilter_io_temac_tx_valid;
  wire[7:0] PacketFilter_io_temac_tx_data;
  wire PacketFilter_io_temac_tx_last;
  wire PacketFilter_io_core_tx_ready;
  wire PacketFilter_io_keyInfo_valid;
  wire[7:0] PacketFilter_io_keyInfo_bits_len;
  wire[3:0] PacketFilter_io_keyInfo_bits_tag;
  wire PacketFilter_io_keyData_valid;
  wire[7:0] PacketFilter_io_keyData_bits;
  wire PacketFilter_io_resultInfo_ready;
  wire PacketFilter_io_resultData_ready;
  wire KeyValueStore_io_keyInfo_ready;
  wire KeyValueStore_io_keyData_ready;
  wire KeyValueStore_io_resultInfo_valid;
  wire[18:0] KeyValueStore_io_resultInfo_bits_len;
  wire[3:0] KeyValueStore_io_resultInfo_bits_tag;
  wire KeyValueStore_io_resultData_valid;
  wire[7:0] KeyValueStore_io_resultData_bits;
  wire KeyValueStore_io_readready;
  wire KeyValueStore_io_rocc_cmd_ready;
  wire KeyValueStore_io_rocc_resp_valid;
  wire[4:0] KeyValueStore_io_rocc_resp_bits_rd;
  wire[63:0] KeyValueStore_io_rocc_resp_bits_data;
  wire KeyValueStore_io_rocc_mem_req_valid;
  wire KeyValueStore_io_rocc_mem_req_bits_kill;
  wire[2:0] KeyValueStore_io_rocc_mem_req_bits_typ;
  wire KeyValueStore_io_rocc_mem_req_bits_phys;
  wire[42:0] KeyValueStore_io_rocc_mem_req_bits_addr;
  wire[4:0] KeyValueStore_io_rocc_mem_req_bits_cmd;
  wire KeyValueStore_io_rocc_busy;
  wire KeyValueStore_io_rocc_interrupt;
  wire KeyValueStore_io_rocc_imem_acquire_valid;
  wire KeyValueStore_io_rocc_imem_grant_ready;
  wire KeyValueStore_io_rocc_imem_finish_valid;
  wire KeyValueStore_io_rocc_iptw_req_valid;
  wire KeyValueStore_io_rocc_dptw_req_valid;
  wire KeyValueStore_io_rocc_pptw_req_valid;
  wire core_io_tilelink_acquire_valid;
  wire[1:0] core_io_tilelink_acquire_bits_header_src;
  wire[1:0] core_io_tilelink_acquire_bits_header_dst;
  wire[25:0] core_io_tilelink_acquire_bits_payload_addr;
  wire[2:0] core_io_tilelink_acquire_bits_payload_client_xact_id;
  wire[511:0] core_io_tilelink_acquire_bits_payload_data;
  wire core_io_tilelink_acquire_bits_payload_uncached;
  wire[1:0] core_io_tilelink_acquire_bits_payload_a_type;
  wire[511:0] core_io_tilelink_acquire_bits_payload_subblock;
  wire core_io_tilelink_grant_ready;
  wire core_io_tilelink_finish_valid;
  wire[1:0] core_io_tilelink_finish_bits_header_src;
  wire[1:0] core_io_tilelink_finish_bits_header_dst;
  wire[2:0] core_io_tilelink_finish_bits_payload_master_xact_id;
  wire core_io_tilelink_probe_ready;
  wire core_io_tilelink_release_valid;
  wire[1:0] core_io_tilelink_release_bits_header_src;
  wire[1:0] core_io_tilelink_release_bits_header_dst;
  wire[25:0] core_io_tilelink_release_bits_payload_addr;
  wire[2:0] core_io_tilelink_release_bits_payload_client_xact_id;
  wire[511:0] core_io_tilelink_release_bits_payload_data;
  wire[2:0] core_io_tilelink_release_bits_payload_r_type;
  wire core_io_host_pcr_req_ready;
  wire core_io_host_pcr_rep_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_pcr;
  wire core_io_temac_rx_axis_fifo_tready;
  wire[7:0] core_io_temac_tx_axis_fifo_tdata;
  wire core_io_temac_tx_axis_fifo_tvalid;
  wire core_io_temac_tx_axis_fifo_tlast;
  wire[11:0] core_io_temac_s_axi_awaddr;
  wire core_io_temac_s_axi_awvalid;
  wire[31:0] core_io_temac_s_axi_wdata;
  wire core_io_temac_s_axi_wvalid;
  wire core_io_temac_s_axi_bready;
  wire[11:0] core_io_temac_s_axi_araddr;
  wire core_io_temac_s_axi_arvalid;
  wire core_io_temac_s_axi_rready;
  wire core_io_temac_sfp_tx_disable;
  wire core_io_rocc_cmd_valid;
  wire[6:0] core_io_rocc_cmd_bits_inst_funct;
  wire[4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire core_io_rocc_cmd_bits_inst_xd;
  wire core_io_rocc_cmd_bits_inst_xs1;
  wire core_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] core_io_rocc_cmd_bits_inst_rd;
  wire[6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] core_io_rocc_cmd_bits_rs1;
  wire[63:0] core_io_rocc_cmd_bits_rs2;
  wire core_io_rocc_resp_ready;
  wire core_io_rocc_mem_req_ready;
  wire core_io_rocc_mem_resp_valid;
  wire[63:0] core_io_rocc_mem_resp_bits_data;
  wire core_io_rocc_mem_resp_bits_nack;
  wire core_io_rocc_mem_resp_bits_replay;
  wire[2:0] core_io_rocc_mem_resp_bits_typ;
  wire core_io_rocc_mem_resp_bits_has_data;
  wire[63:0] core_io_rocc_mem_resp_bits_data_subword;
  wire[8:0] core_io_rocc_mem_resp_bits_tag;
  wire[3:0] core_io_rocc_mem_resp_bits_cmd;
  wire[43:0] core_io_rocc_mem_resp_bits_addr;
  wire[63:0] core_io_rocc_mem_resp_bits_store_data;
  wire core_io_rocc_s;
  wire core_io_rocc_imem_acquire_ready;
  wire core_io_rocc_imem_grant_valid;
  wire[1:0] core_io_rocc_imem_grant_bits_header_src;
  wire[1:0] core_io_rocc_imem_grant_bits_header_dst;
  wire[511:0] core_io_rocc_imem_grant_bits_payload_data;
  wire[2:0] core_io_rocc_imem_grant_bits_payload_client_xact_id;
  wire[2:0] core_io_rocc_imem_grant_bits_payload_master_xact_id;
  wire[1:0] core_io_rocc_imem_grant_bits_payload_g_type;
  wire core_io_rocc_imem_finish_ready;
  wire core_io_rocc_iptw_req_ready;
  wire core_io_rocc_iptw_resp_valid;
  wire core_io_rocc_iptw_resp_bits_error;
  wire[18:0] core_io_rocc_iptw_resp_bits_ppn;
  wire[5:0] core_io_rocc_iptw_resp_bits_perm;
  wire[7:0] core_io_rocc_iptw_status_ip;
  wire[7:0] core_io_rocc_iptw_status_im;
  wire[6:0] core_io_rocc_iptw_status_zero;
  wire core_io_rocc_iptw_status_er;
  wire core_io_rocc_iptw_status_vm;
  wire core_io_rocc_iptw_status_s64;
  wire core_io_rocc_iptw_status_u64;
  wire core_io_rocc_iptw_status_ef;
  wire core_io_rocc_iptw_status_pei;
  wire core_io_rocc_iptw_status_ei;
  wire core_io_rocc_iptw_status_ps;
  wire core_io_rocc_iptw_status_s;
  wire core_io_rocc_iptw_invalidate;
  wire core_io_rocc_iptw_sret;
  wire core_io_rocc_dptw_req_ready;
  wire core_io_rocc_dptw_resp_valid;
  wire core_io_rocc_dptw_resp_bits_error;
  wire[18:0] core_io_rocc_dptw_resp_bits_ppn;
  wire[5:0] core_io_rocc_dptw_resp_bits_perm;
  wire[7:0] core_io_rocc_dptw_status_ip;
  wire[7:0] core_io_rocc_dptw_status_im;
  wire[6:0] core_io_rocc_dptw_status_zero;
  wire core_io_rocc_dptw_status_er;
  wire core_io_rocc_dptw_status_vm;
  wire core_io_rocc_dptw_status_s64;
  wire core_io_rocc_dptw_status_u64;
  wire core_io_rocc_dptw_status_ef;
  wire core_io_rocc_dptw_status_pei;
  wire core_io_rocc_dptw_status_ei;
  wire core_io_rocc_dptw_status_ps;
  wire core_io_rocc_dptw_status_s;
  wire core_io_rocc_dptw_invalidate;
  wire core_io_rocc_dptw_sret;
  wire core_io_rocc_pptw_req_ready;
  wire core_io_rocc_pptw_resp_valid;
  wire core_io_rocc_pptw_resp_bits_error;
  wire[18:0] core_io_rocc_pptw_resp_bits_ppn;
  wire[5:0] core_io_rocc_pptw_resp_bits_perm;
  wire[7:0] core_io_rocc_pptw_status_ip;
  wire[7:0] core_io_rocc_pptw_status_im;
  wire[6:0] core_io_rocc_pptw_status_zero;
  wire core_io_rocc_pptw_status_er;
  wire core_io_rocc_pptw_status_vm;
  wire core_io_rocc_pptw_status_s64;
  wire core_io_rocc_pptw_status_u64;
  wire core_io_rocc_pptw_status_ef;
  wire core_io_rocc_pptw_status_pei;
  wire core_io_rocc_pptw_status_ei;
  wire core_io_rocc_pptw_status_ps;
  wire core_io_rocc_pptw_status_s;
  wire core_io_rocc_pptw_invalidate;
  wire core_io_rocc_pptw_sret;
  wire core_io_rocc_exception;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_pcr;
  wire uncore_io_mem_req_cmd_valid;
  wire[25:0] uncore_io_mem_req_cmd_bits_addr;
  wire[4:0] uncore_io_mem_req_cmd_bits_tag;
  wire uncore_io_mem_req_cmd_bits_rw;
  wire uncore_io_mem_req_data_valid;
  wire[127:0] uncore_io_mem_req_data_bits_data;
  wire uncore_io_tiles_0_acquire_ready;
  wire uncore_io_tiles_0_grant_valid;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_src;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_dst;
  wire[511:0] uncore_io_tiles_0_grant_bits_payload_data;
  wire[2:0] uncore_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[2:0] uncore_io_tiles_0_grant_bits_payload_master_xact_id;
  wire uncore_io_tiles_0_grant_bits_payload_uncached;
  wire[1:0] uncore_io_tiles_0_grant_bits_payload_g_type;
  wire uncore_io_tiles_0_finish_ready;
  wire uncore_io_tiles_0_probe_valid;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_src;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_dst;
  wire[25:0] uncore_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] uncore_io_tiles_0_probe_bits_payload_p_type;
  wire uncore_io_tiles_0_release_ready;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_pcr_req_valid;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire[4:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire uncore_io_htif_0_ipi_req_ready;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_rep_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
    R6 = {1{$random}};
  end
`endif

  assign resetSigs_0 = uncore_io_htif_0_reset;
  assign T2 = {3'h0, core_io_rocc_imem_grant_bits_payload_g_type};
  assign T3 = core_io_rocc_mem_resp_bits_addr[6'h2a:1'h0];
  assign T4 = {1'h0, KeyValueStore_io_rocc_mem_req_bits_addr};
  assign io_debug_rocc_inst_bits_rs2 = core_io_rocc_cmd_bits_rs2;
  assign io_debug_rocc_inst_bits_rs1 = core_io_rocc_cmd_bits_rs1;
  assign io_debug_rocc_inst_bits_inst_opcode = core_io_rocc_cmd_bits_inst_opcode;
  assign io_debug_rocc_inst_bits_inst_rd = core_io_rocc_cmd_bits_inst_rd;
  assign io_debug_rocc_inst_bits_inst_xs2 = core_io_rocc_cmd_bits_inst_xs2;
  assign io_debug_rocc_inst_bits_inst_xs1 = core_io_rocc_cmd_bits_inst_xs1;
  assign io_debug_rocc_inst_bits_inst_xd = core_io_rocc_cmd_bits_inst_xd;
  assign io_debug_rocc_inst_bits_inst_rs1 = core_io_rocc_cmd_bits_inst_rs1;
  assign io_debug_rocc_inst_bits_inst_rs2 = core_io_rocc_cmd_bits_inst_rs2;
  assign io_debug_rocc_inst_bits_inst_funct = core_io_rocc_cmd_bits_inst_funct;
  assign io_debug_rocc_inst_valid = core_io_rocc_cmd_valid;
  assign io_debug_rocc_inst_ready = KeyValueStore_io_rocc_cmd_ready;
  assign io_debug_readready = KeyValueStore_io_readready;
  assign io_debug_resultData_bits = KeyValueStore_io_resultData_bits;
  assign io_debug_resultData_valid = KeyValueStore_io_resultData_valid;
  assign io_debug_resultLen_bits = T0;
  assign T0 = KeyValueStore_io_resultInfo_bits_len[4'hf:1'h0];
  assign io_debug_resultLen_valid = KeyValueStore_io_resultInfo_valid;
  assign io_debug_keyData_bits = PacketFilter_io_keyData_bits;
  assign io_debug_keyData_valid = PacketFilter_io_keyData_valid;
  assign io_debug_keyLen_bits = T1;
  assign T1 = {8'h0, PacketFilter_io_keyInfo_bits_len};
  assign io_debug_keyLen_valid = PacketFilter_io_keyInfo_valid;
  assign io_temac_sfp_tx_disable = core_io_temac_sfp_tx_disable;
  assign io_temac_s_axi_rready = core_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = core_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = core_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = core_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = core_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = core_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = core_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = core_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = PacketFilter_io_temac_tx_last;
  assign io_temac_tx_axis_fifo_tvalid = PacketFilter_io_temac_tx_valid;
  assign io_temac_tx_axis_fifo_tdata = PacketFilter_io_temac_tx_data;
  assign io_temac_rx_axis_fifo_tready = PacketFilter_io_temac_rx_ready;
  assign io_mem_req_data_bits_data = uncore_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = uncore_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = uncore_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = uncore_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = uncore_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = uncore_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = uncore_io_host_debug_stats_pcr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  RocketTile core(.clk(clk), .reset(resetSigs_0),
       .io_tilelink_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tilelink_acquire_valid( core_io_tilelink_acquire_valid ),
       .io_tilelink_acquire_bits_header_src( core_io_tilelink_acquire_bits_header_src ),
       .io_tilelink_acquire_bits_header_dst( core_io_tilelink_acquire_bits_header_dst ),
       .io_tilelink_acquire_bits_payload_addr( core_io_tilelink_acquire_bits_payload_addr ),
       .io_tilelink_acquire_bits_payload_client_xact_id( core_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tilelink_acquire_bits_payload_data( core_io_tilelink_acquire_bits_payload_data ),
       .io_tilelink_acquire_bits_payload_uncached( core_io_tilelink_acquire_bits_payload_uncached ),
       .io_tilelink_acquire_bits_payload_a_type( core_io_tilelink_acquire_bits_payload_a_type ),
       .io_tilelink_acquire_bits_payload_subblock( core_io_tilelink_acquire_bits_payload_subblock ),
       .io_tilelink_grant_ready( core_io_tilelink_grant_ready ),
       .io_tilelink_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tilelink_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tilelink_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tilelink_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tilelink_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tilelink_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tilelink_grant_bits_payload_uncached( uncore_io_tiles_0_grant_bits_payload_uncached ),
       .io_tilelink_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tilelink_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tilelink_finish_valid( core_io_tilelink_finish_valid ),
       .io_tilelink_finish_bits_header_src( core_io_tilelink_finish_bits_header_src ),
       .io_tilelink_finish_bits_header_dst( core_io_tilelink_finish_bits_header_dst ),
       .io_tilelink_finish_bits_payload_master_xact_id( core_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tilelink_probe_ready( core_io_tilelink_probe_ready ),
       .io_tilelink_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tilelink_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tilelink_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tilelink_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tilelink_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tilelink_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tilelink_release_valid( core_io_tilelink_release_valid ),
       .io_tilelink_release_bits_header_src( core_io_tilelink_release_bits_header_src ),
       .io_tilelink_release_bits_header_dst( core_io_tilelink_release_bits_header_dst ),
       .io_tilelink_release_bits_payload_addr( core_io_tilelink_release_bits_payload_addr ),
       .io_tilelink_release_bits_payload_client_xact_id( core_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tilelink_release_bits_payload_data( core_io_tilelink_release_bits_payload_data ),
       .io_tilelink_release_bits_payload_r_type( core_io_tilelink_release_bits_payload_r_type ),
       .io_host_reset( R5 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_0_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_0_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_temac_rx_axis_fifo_tdata( PacketFilter_io_core_rx_data ),
       .io_temac_rx_axis_fifo_tvalid( PacketFilter_io_core_rx_valid ),
       .io_temac_rx_axis_fifo_tready( core_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( PacketFilter_io_core_rx_last ),
       .io_temac_tx_axis_fifo_tdata( core_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( core_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( PacketFilter_io_core_tx_ready ),
       .io_temac_tx_axis_fifo_tlast( core_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( core_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( core_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( core_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( core_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( core_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( core_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( core_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( core_io_temac_s_axi_rready ),
       .io_temac_sfp_tx_disable( core_io_temac_sfp_tx_disable ),
       .io_rocc_cmd_ready( KeyValueStore_io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( core_io_rocc_cmd_valid ),
       .io_rocc_cmd_bits_inst_funct( core_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( core_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( core_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( core_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( core_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( core_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( core_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( core_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( core_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( core_io_rocc_cmd_bits_rs2 ),
       .io_rocc_resp_ready( core_io_rocc_resp_ready ),
       .io_rocc_resp_valid( KeyValueStore_io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( KeyValueStore_io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( KeyValueStore_io_rocc_resp_bits_data ),
       .io_rocc_mem_req_ready( core_io_rocc_mem_req_ready ),
       .io_rocc_mem_req_valid( KeyValueStore_io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( KeyValueStore_io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( KeyValueStore_io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( KeyValueStore_io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( T4 ),
       //.io_rocc_mem_req_bits_tag(  )
       .io_rocc_mem_req_bits_cmd( KeyValueStore_io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_req_bits_data(  )
       .io_rocc_mem_resp_valid( core_io_rocc_mem_resp_valid ),
       .io_rocc_mem_resp_bits_data( core_io_rocc_mem_resp_bits_data ),
       .io_rocc_mem_resp_bits_nack( core_io_rocc_mem_resp_bits_nack ),
       .io_rocc_mem_resp_bits_replay( core_io_rocc_mem_resp_bits_replay ),
       .io_rocc_mem_resp_bits_typ( core_io_rocc_mem_resp_bits_typ ),
       .io_rocc_mem_resp_bits_has_data( core_io_rocc_mem_resp_bits_has_data ),
       .io_rocc_mem_resp_bits_data_subword( core_io_rocc_mem_resp_bits_data_subword ),
       .io_rocc_mem_resp_bits_tag( core_io_rocc_mem_resp_bits_tag ),
       .io_rocc_mem_resp_bits_cmd( core_io_rocc_mem_resp_bits_cmd ),
       .io_rocc_mem_resp_bits_addr( core_io_rocc_mem_resp_bits_addr ),
       .io_rocc_mem_resp_bits_store_data( core_io_rocc_mem_resp_bits_store_data ),
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( KeyValueStore_io_rocc_busy ),
       .io_rocc_s( core_io_rocc_s ),
       .io_rocc_interrupt( KeyValueStore_io_rocc_interrupt ),
       .io_rocc_imem_acquire_ready( core_io_rocc_imem_acquire_ready ),
       .io_rocc_imem_acquire_valid( KeyValueStore_io_rocc_imem_acquire_valid ),
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_uncached(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_subblock(  )
       .io_rocc_imem_grant_ready( KeyValueStore_io_rocc_imem_grant_ready ),
       .io_rocc_imem_grant_valid( core_io_rocc_imem_grant_valid ),
       .io_rocc_imem_grant_bits_header_src( core_io_rocc_imem_grant_bits_header_src ),
       .io_rocc_imem_grant_bits_header_dst( core_io_rocc_imem_grant_bits_header_dst ),
       .io_rocc_imem_grant_bits_payload_data( core_io_rocc_imem_grant_bits_payload_data ),
       .io_rocc_imem_grant_bits_payload_client_xact_id( core_io_rocc_imem_grant_bits_payload_client_xact_id ),
       .io_rocc_imem_grant_bits_payload_master_xact_id( core_io_rocc_imem_grant_bits_payload_master_xact_id ),
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       .io_rocc_imem_grant_bits_payload_g_type( core_io_rocc_imem_grant_bits_payload_g_type ),
       .io_rocc_imem_finish_ready( core_io_rocc_imem_finish_ready ),
       .io_rocc_imem_finish_valid( KeyValueStore_io_rocc_imem_finish_valid ),
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       .io_rocc_iptw_req_ready( core_io_rocc_iptw_req_ready ),
       .io_rocc_iptw_req_valid( KeyValueStore_io_rocc_iptw_req_valid ),
       //.io_rocc_iptw_req_bits(  )
       .io_rocc_iptw_resp_valid( core_io_rocc_iptw_resp_valid ),
       .io_rocc_iptw_resp_bits_error( core_io_rocc_iptw_resp_bits_error ),
       .io_rocc_iptw_resp_bits_ppn( core_io_rocc_iptw_resp_bits_ppn ),
       .io_rocc_iptw_resp_bits_perm( core_io_rocc_iptw_resp_bits_perm ),
       .io_rocc_iptw_status_ip( core_io_rocc_iptw_status_ip ),
       .io_rocc_iptw_status_im( core_io_rocc_iptw_status_im ),
       .io_rocc_iptw_status_zero( core_io_rocc_iptw_status_zero ),
       .io_rocc_iptw_status_er( core_io_rocc_iptw_status_er ),
       .io_rocc_iptw_status_vm( core_io_rocc_iptw_status_vm ),
       .io_rocc_iptw_status_s64( core_io_rocc_iptw_status_s64 ),
       .io_rocc_iptw_status_u64( core_io_rocc_iptw_status_u64 ),
       .io_rocc_iptw_status_ef( core_io_rocc_iptw_status_ef ),
       .io_rocc_iptw_status_pei( core_io_rocc_iptw_status_pei ),
       .io_rocc_iptw_status_ei( core_io_rocc_iptw_status_ei ),
       .io_rocc_iptw_status_ps( core_io_rocc_iptw_status_ps ),
       .io_rocc_iptw_status_s( core_io_rocc_iptw_status_s ),
       .io_rocc_iptw_invalidate( core_io_rocc_iptw_invalidate ),
       .io_rocc_iptw_sret( core_io_rocc_iptw_sret ),
       .io_rocc_dptw_req_ready( core_io_rocc_dptw_req_ready ),
       .io_rocc_dptw_req_valid( KeyValueStore_io_rocc_dptw_req_valid ),
       //.io_rocc_dptw_req_bits(  )
       .io_rocc_dptw_resp_valid( core_io_rocc_dptw_resp_valid ),
       .io_rocc_dptw_resp_bits_error( core_io_rocc_dptw_resp_bits_error ),
       .io_rocc_dptw_resp_bits_ppn( core_io_rocc_dptw_resp_bits_ppn ),
       .io_rocc_dptw_resp_bits_perm( core_io_rocc_dptw_resp_bits_perm ),
       .io_rocc_dptw_status_ip( core_io_rocc_dptw_status_ip ),
       .io_rocc_dptw_status_im( core_io_rocc_dptw_status_im ),
       .io_rocc_dptw_status_zero( core_io_rocc_dptw_status_zero ),
       .io_rocc_dptw_status_er( core_io_rocc_dptw_status_er ),
       .io_rocc_dptw_status_vm( core_io_rocc_dptw_status_vm ),
       .io_rocc_dptw_status_s64( core_io_rocc_dptw_status_s64 ),
       .io_rocc_dptw_status_u64( core_io_rocc_dptw_status_u64 ),
       .io_rocc_dptw_status_ef( core_io_rocc_dptw_status_ef ),
       .io_rocc_dptw_status_pei( core_io_rocc_dptw_status_pei ),
       .io_rocc_dptw_status_ei( core_io_rocc_dptw_status_ei ),
       .io_rocc_dptw_status_ps( core_io_rocc_dptw_status_ps ),
       .io_rocc_dptw_status_s( core_io_rocc_dptw_status_s ),
       .io_rocc_dptw_invalidate( core_io_rocc_dptw_invalidate ),
       .io_rocc_dptw_sret( core_io_rocc_dptw_sret ),
       .io_rocc_pptw_req_ready( core_io_rocc_pptw_req_ready ),
       .io_rocc_pptw_req_valid( KeyValueStore_io_rocc_pptw_req_valid ),
       //.io_rocc_pptw_req_bits(  )
       .io_rocc_pptw_resp_valid( core_io_rocc_pptw_resp_valid ),
       .io_rocc_pptw_resp_bits_error( core_io_rocc_pptw_resp_bits_error ),
       .io_rocc_pptw_resp_bits_ppn( core_io_rocc_pptw_resp_bits_ppn ),
       .io_rocc_pptw_resp_bits_perm( core_io_rocc_pptw_resp_bits_perm ),
       .io_rocc_pptw_status_ip( core_io_rocc_pptw_status_ip ),
       .io_rocc_pptw_status_im( core_io_rocc_pptw_status_im ),
       .io_rocc_pptw_status_zero( core_io_rocc_pptw_status_zero ),
       .io_rocc_pptw_status_er( core_io_rocc_pptw_status_er ),
       .io_rocc_pptw_status_vm( core_io_rocc_pptw_status_vm ),
       .io_rocc_pptw_status_s64( core_io_rocc_pptw_status_s64 ),
       .io_rocc_pptw_status_u64( core_io_rocc_pptw_status_u64 ),
       .io_rocc_pptw_status_ef( core_io_rocc_pptw_status_ef ),
       .io_rocc_pptw_status_pei( core_io_rocc_pptw_status_pei ),
       .io_rocc_pptw_status_ei( core_io_rocc_pptw_status_ei ),
       .io_rocc_pptw_status_ps( core_io_rocc_pptw_status_ps ),
       .io_rocc_pptw_status_s( core_io_rocc_pptw_status_s ),
       .io_rocc_pptw_invalidate( core_io_rocc_pptw_invalidate ),
       .io_rocc_pptw_sret( core_io_rocc_pptw_sret ),
       .io_rocc_exception( core_io_rocc_exception )
  );
  `ifndef SYNTHESIS
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_ptw_req_ready = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_valid = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_error = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_ppn = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_perm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ip = {1{$random}};
    assign core.io_rocc_mem_ptw_status_im = {1{$random}};
    assign core.io_rocc_mem_ptw_status_zero = {1{$random}};
    assign core.io_rocc_mem_ptw_status_er = {1{$random}};
    assign core.io_rocc_mem_ptw_status_vm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_u64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ef = {1{$random}};
    assign core.io_rocc_mem_ptw_status_pei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ps = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s = {1{$random}};
    assign core.io_rocc_mem_ptw_invalidate = {1{$random}};
    assign core.io_rocc_mem_ptw_sret = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_data = {16{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_uncached = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_subblock = {16{$random}};
    assign core.io_rocc_imem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_finish_bits_payload_master_xact_id = {1{$random}};
    assign core.io_rocc_iptw_req_bits = {1{$random}};
    assign core.io_rocc_dptw_req_bits = {1{$random}};
    assign core.io_rocc_pptw_req_bits = {1{$random}};
  `endif
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_pcr( uncore_io_host_debug_stats_pcr ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( uncore_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( uncore_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( uncore_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( uncore_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( uncore_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( uncore_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_tiles_0_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( core_io_tilelink_acquire_valid ),
       .io_tiles_0_acquire_bits_header_src( core_io_tilelink_acquire_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( core_io_tilelink_acquire_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( core_io_tilelink_acquire_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( core_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( core_io_tilelink_acquire_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_uncached( core_io_tilelink_acquire_bits_payload_uncached ),
       .io_tiles_0_acquire_bits_payload_a_type( core_io_tilelink_acquire_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_subblock( core_io_tilelink_acquire_bits_payload_subblock ),
       .io_tiles_0_grant_ready( core_io_tilelink_grant_ready ),
       .io_tiles_0_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_uncached( uncore_io_tiles_0_grant_bits_payload_uncached ),
       .io_tiles_0_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( core_io_tilelink_finish_valid ),
       .io_tiles_0_finish_bits_header_src( core_io_tilelink_finish_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( core_io_tilelink_finish_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( core_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( core_io_tilelink_probe_ready ),
       .io_tiles_0_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( core_io_tilelink_release_valid ),
       .io_tiles_0_release_bits_header_src( core_io_tilelink_release_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( core_io_tilelink_release_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( core_io_tilelink_release_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( core_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_data( core_io_tilelink_release_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( core_io_tilelink_release_bits_payload_r_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_0_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_incoherent_0( uncore_io_htif_0_reset )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  `ifndef SYNTHESIS
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
  `endif
  Queue_0 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( core_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_0_io_deq_bits_data )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( core_io_host_pcr_rep_valid ),
       .io_enq_bits( core_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( core_io_host_ipi_req_valid ),
       .io_enq_bits( core_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( core_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
  );
  KeyValueStore KeyValueStore(.clk(clk), .reset(reset),
       .io_keyInfo_ready( KeyValueStore_io_keyInfo_ready ),
       .io_keyInfo_valid( PacketFilter_io_keyInfo_valid ),
       .io_keyInfo_bits_len( PacketFilter_io_keyInfo_bits_len ),
       .io_keyInfo_bits_tag( PacketFilter_io_keyInfo_bits_tag ),
       .io_keyData_ready( KeyValueStore_io_keyData_ready ),
       .io_keyData_valid( PacketFilter_io_keyData_valid ),
       .io_keyData_bits( PacketFilter_io_keyData_bits ),
       .io_resultInfo_ready( PacketFilter_io_resultInfo_ready ),
       .io_resultInfo_valid( KeyValueStore_io_resultInfo_valid ),
       .io_resultInfo_bits_len( KeyValueStore_io_resultInfo_bits_len ),
       .io_resultInfo_bits_tag( KeyValueStore_io_resultInfo_bits_tag ),
       .io_resultData_ready( PacketFilter_io_resultData_ready ),
       .io_resultData_valid( KeyValueStore_io_resultData_valid ),
       .io_resultData_bits( KeyValueStore_io_resultData_bits ),
       //.io_writeready(  )
       .io_readready( KeyValueStore_io_readready ),
       .io_rocc_cmd_ready( KeyValueStore_io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( core_io_rocc_cmd_valid ),
       .io_rocc_cmd_bits_inst_funct( core_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( core_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( core_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( core_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( core_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( core_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( core_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( core_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( core_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( core_io_rocc_cmd_bits_rs2 ),
       .io_rocc_resp_ready( core_io_rocc_resp_ready ),
       .io_rocc_resp_valid( KeyValueStore_io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( KeyValueStore_io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( KeyValueStore_io_rocc_resp_bits_data ),
       .io_rocc_mem_req_ready( core_io_rocc_mem_req_ready ),
       .io_rocc_mem_req_valid( KeyValueStore_io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( KeyValueStore_io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( KeyValueStore_io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( KeyValueStore_io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( KeyValueStore_io_rocc_mem_req_bits_addr ),
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_req_bits_tag(  )
       .io_rocc_mem_req_bits_cmd( KeyValueStore_io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_resp_valid( core_io_rocc_mem_resp_valid ),
       .io_rocc_mem_resp_bits_nack( core_io_rocc_mem_resp_bits_nack ),
       .io_rocc_mem_resp_bits_replay( core_io_rocc_mem_resp_bits_replay ),
       .io_rocc_mem_resp_bits_typ( core_io_rocc_mem_resp_bits_typ ),
       .io_rocc_mem_resp_bits_has_data( core_io_rocc_mem_resp_bits_has_data ),
       .io_rocc_mem_resp_bits_data( core_io_rocc_mem_resp_bits_data ),
       .io_rocc_mem_resp_bits_data_subword( core_io_rocc_mem_resp_bits_data_subword ),
       .io_rocc_mem_resp_bits_tag( core_io_rocc_mem_resp_bits_tag ),
       .io_rocc_mem_resp_bits_cmd( core_io_rocc_mem_resp_bits_cmd ),
       .io_rocc_mem_resp_bits_addr( T3 ),
       .io_rocc_mem_resp_bits_store_data( core_io_rocc_mem_resp_bits_store_data ),
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( KeyValueStore_io_rocc_busy ),
       .io_rocc_s( core_io_rocc_s ),
       .io_rocc_interrupt( KeyValueStore_io_rocc_interrupt ),
       .io_rocc_imem_acquire_ready( core_io_rocc_imem_acquire_ready ),
       .io_rocc_imem_acquire_valid( KeyValueStore_io_rocc_imem_acquire_valid ),
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_write_mask(  )
       //.io_rocc_imem_acquire_bits_payload_subword_addr(  )
       //.io_rocc_imem_acquire_bits_payload_atomic_opcode(  )
       .io_rocc_imem_grant_ready( KeyValueStore_io_rocc_imem_grant_ready ),
       .io_rocc_imem_grant_valid( core_io_rocc_imem_grant_valid ),
       .io_rocc_imem_grant_bits_header_src( core_io_rocc_imem_grant_bits_header_src ),
       .io_rocc_imem_grant_bits_header_dst( core_io_rocc_imem_grant_bits_header_dst ),
       .io_rocc_imem_grant_bits_payload_data( core_io_rocc_imem_grant_bits_payload_data ),
       .io_rocc_imem_grant_bits_payload_client_xact_id( core_io_rocc_imem_grant_bits_payload_client_xact_id ),
       .io_rocc_imem_grant_bits_payload_master_xact_id( core_io_rocc_imem_grant_bits_payload_master_xact_id ),
       .io_rocc_imem_grant_bits_payload_g_type( T2 ),
       .io_rocc_imem_finish_ready( core_io_rocc_imem_finish_ready ),
       .io_rocc_imem_finish_valid( KeyValueStore_io_rocc_imem_finish_valid ),
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       .io_rocc_iptw_req_ready( core_io_rocc_iptw_req_ready ),
       .io_rocc_iptw_req_valid( KeyValueStore_io_rocc_iptw_req_valid ),
       //.io_rocc_iptw_req_bits(  )
       .io_rocc_iptw_resp_valid( core_io_rocc_iptw_resp_valid ),
       .io_rocc_iptw_resp_bits_error( core_io_rocc_iptw_resp_bits_error ),
       .io_rocc_iptw_resp_bits_ppn( core_io_rocc_iptw_resp_bits_ppn ),
       .io_rocc_iptw_resp_bits_perm( core_io_rocc_iptw_resp_bits_perm ),
       .io_rocc_iptw_status_ip( core_io_rocc_iptw_status_ip ),
       .io_rocc_iptw_status_im( core_io_rocc_iptw_status_im ),
       .io_rocc_iptw_status_zero( core_io_rocc_iptw_status_zero ),
       .io_rocc_iptw_status_er( core_io_rocc_iptw_status_er ),
       .io_rocc_iptw_status_vm( core_io_rocc_iptw_status_vm ),
       .io_rocc_iptw_status_s64( core_io_rocc_iptw_status_s64 ),
       .io_rocc_iptw_status_u64( core_io_rocc_iptw_status_u64 ),
       .io_rocc_iptw_status_ef( core_io_rocc_iptw_status_ef ),
       .io_rocc_iptw_status_pei( core_io_rocc_iptw_status_pei ),
       .io_rocc_iptw_status_ei( core_io_rocc_iptw_status_ei ),
       .io_rocc_iptw_status_ps( core_io_rocc_iptw_status_ps ),
       .io_rocc_iptw_status_s( core_io_rocc_iptw_status_s ),
       .io_rocc_iptw_invalidate( core_io_rocc_iptw_invalidate ),
       .io_rocc_iptw_sret( core_io_rocc_iptw_sret ),
       .io_rocc_dptw_req_ready( core_io_rocc_dptw_req_ready ),
       .io_rocc_dptw_req_valid( KeyValueStore_io_rocc_dptw_req_valid ),
       //.io_rocc_dptw_req_bits(  )
       .io_rocc_dptw_resp_valid( core_io_rocc_dptw_resp_valid ),
       .io_rocc_dptw_resp_bits_error( core_io_rocc_dptw_resp_bits_error ),
       .io_rocc_dptw_resp_bits_ppn( core_io_rocc_dptw_resp_bits_ppn ),
       .io_rocc_dptw_resp_bits_perm( core_io_rocc_dptw_resp_bits_perm ),
       .io_rocc_dptw_status_ip( core_io_rocc_dptw_status_ip ),
       .io_rocc_dptw_status_im( core_io_rocc_dptw_status_im ),
       .io_rocc_dptw_status_zero( core_io_rocc_dptw_status_zero ),
       .io_rocc_dptw_status_er( core_io_rocc_dptw_status_er ),
       .io_rocc_dptw_status_vm( core_io_rocc_dptw_status_vm ),
       .io_rocc_dptw_status_s64( core_io_rocc_dptw_status_s64 ),
       .io_rocc_dptw_status_u64( core_io_rocc_dptw_status_u64 ),
       .io_rocc_dptw_status_ef( core_io_rocc_dptw_status_ef ),
       .io_rocc_dptw_status_pei( core_io_rocc_dptw_status_pei ),
       .io_rocc_dptw_status_ei( core_io_rocc_dptw_status_ei ),
       .io_rocc_dptw_status_ps( core_io_rocc_dptw_status_ps ),
       .io_rocc_dptw_status_s( core_io_rocc_dptw_status_s ),
       .io_rocc_dptw_invalidate( core_io_rocc_dptw_invalidate ),
       .io_rocc_dptw_sret( core_io_rocc_dptw_sret ),
       .io_rocc_pptw_req_ready( core_io_rocc_pptw_req_ready ),
       .io_rocc_pptw_req_valid( KeyValueStore_io_rocc_pptw_req_valid ),
       //.io_rocc_pptw_req_bits(  )
       .io_rocc_pptw_resp_valid( core_io_rocc_pptw_resp_valid ),
       .io_rocc_pptw_resp_bits_error( core_io_rocc_pptw_resp_bits_error ),
       .io_rocc_pptw_resp_bits_ppn( core_io_rocc_pptw_resp_bits_ppn ),
       .io_rocc_pptw_resp_bits_perm( core_io_rocc_pptw_resp_bits_perm ),
       .io_rocc_pptw_status_ip( core_io_rocc_pptw_status_ip ),
       .io_rocc_pptw_status_im( core_io_rocc_pptw_status_im ),
       .io_rocc_pptw_status_zero( core_io_rocc_pptw_status_zero ),
       .io_rocc_pptw_status_er( core_io_rocc_pptw_status_er ),
       .io_rocc_pptw_status_vm( core_io_rocc_pptw_status_vm ),
       .io_rocc_pptw_status_s64( core_io_rocc_pptw_status_s64 ),
       .io_rocc_pptw_status_u64( core_io_rocc_pptw_status_u64 ),
       .io_rocc_pptw_status_ef( core_io_rocc_pptw_status_ef ),
       .io_rocc_pptw_status_pei( core_io_rocc_pptw_status_pei ),
       .io_rocc_pptw_status_ei( core_io_rocc_pptw_status_ei ),
       .io_rocc_pptw_status_ps( core_io_rocc_pptw_status_ps ),
       .io_rocc_pptw_status_s( core_io_rocc_pptw_status_s ),
       .io_rocc_pptw_invalidate( core_io_rocc_pptw_invalidate ),
       .io_rocc_pptw_sret( core_io_rocc_pptw_sret ),
       .io_rocc_exception( core_io_rocc_exception )
  );
  `ifndef SYNTHESIS
    assign KeyValueStore.io_rocc_mem_replay_next_valid = {1{$random}};
    assign KeyValueStore.io_rocc_mem_replay_next_bits = {1{$random}};
    assign KeyValueStore.io_rocc_mem_xcpt_ma_ld = {1{$random}};
    assign KeyValueStore.io_rocc_mem_xcpt_ma_st = {1{$random}};
    assign KeyValueStore.io_rocc_mem_xcpt_pf_ld = {1{$random}};
    assign KeyValueStore.io_rocc_mem_xcpt_pf_st = {1{$random}};
    assign KeyValueStore.io_rocc_mem_ptw_req_valid = {1{$random}};
    assign KeyValueStore.io_rocc_mem_ptw_req_bits = {1{$random}};
    assign KeyValueStore.io_rocc_mem_ordered = {1{$random}};
  `endif
  PacketFilter PacketFilter(.clk(clk), .reset(reset),
       .io_temac_rx_ready( PacketFilter_io_temac_rx_ready ),
       .io_temac_rx_valid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_data( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_last( io_temac_rx_axis_fifo_tlast ),
       .io_core_rx_ready( core_io_temac_rx_axis_fifo_tready ),
       .io_core_rx_valid( PacketFilter_io_core_rx_valid ),
       .io_core_rx_data( PacketFilter_io_core_rx_data ),
       .io_core_rx_last( PacketFilter_io_core_rx_last ),
       .io_temac_tx_ready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_valid( PacketFilter_io_temac_tx_valid ),
       .io_temac_tx_data( PacketFilter_io_temac_tx_data ),
       .io_temac_tx_last( PacketFilter_io_temac_tx_last ),
       .io_core_tx_ready( PacketFilter_io_core_tx_ready ),
       .io_core_tx_valid( core_io_temac_tx_axis_fifo_tvalid ),
       .io_core_tx_data( core_io_temac_tx_axis_fifo_tdata ),
       .io_core_tx_last( core_io_temac_tx_axis_fifo_tlast ),
       .io_keyInfo_ready( KeyValueStore_io_keyInfo_ready ),
       .io_keyInfo_valid( PacketFilter_io_keyInfo_valid ),
       .io_keyInfo_bits_len( PacketFilter_io_keyInfo_bits_len ),
       .io_keyInfo_bits_tag( PacketFilter_io_keyInfo_bits_tag ),
       .io_keyData_ready( KeyValueStore_io_keyData_ready ),
       .io_keyData_valid( PacketFilter_io_keyData_valid ),
       .io_keyData_bits( PacketFilter_io_keyData_bits ),
       .io_resultInfo_ready( PacketFilter_io_resultInfo_ready ),
       .io_resultInfo_valid( KeyValueStore_io_resultInfo_valid ),
       .io_resultInfo_bits_len( KeyValueStore_io_resultInfo_bits_len ),
       .io_resultInfo_bits_tag( KeyValueStore_io_resultInfo_bits_tag ),
       .io_resultData_ready( PacketFilter_io_resultData_ready ),
       .io_resultData_valid( KeyValueStore_io_resultData_valid ),
       .io_resultData_bits( KeyValueStore_io_resultData_bits ),
       .io_readready( KeyValueStore_io_readready )
  );

  always @(posedge clk) begin
    R5 <= R6;
    R6 <= uncore_io_htif_0_reset;
  end
endmodule

module UnbankedMem_mem(
  input CLK,
  input RST,
  input init,
  input [6:0] W0A,
  input W0E,
  input [31:0] W0I,
  input [6:0] R1A,
  input R1E,
  output [31:0] R1O
);

reg [31:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [6:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module PacketFilter_getReqLens(
  input CLK,
  input RST,
  input init,
  input [3:0] W0A,
  input W0E,
  input [7:0] W0I,
  input [3:0] R1A,
  input R1E,
  output [7:0] R1O
);

reg [7:0] ram [15:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 16; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [3:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [6:0] W0A,
  input W0E,
  input [83:0] W0I,
  input [83:0] W0M,
  input [6:0] R1A,
  input R1E,
  output [83:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<4; i=i+21) begin
    for (j=1; j<21; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [83:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
    end
  `endif
  reg [6:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][20:0] <= W0I[20:0];
  if (W0E && W0M[21]) ram[W0A][41:21] <= W0I[41:21];
  if (W0E && W0M[42]) ram[W0A][62:42] <= W0I[62:42];
  if (W0E && W0M[63]) ram[W0A][83:63] <= W0I[83:63];
end
assign R1O = ram[reg_R1A];

endmodule


module PacketBuffer_mem(
  input CLK,
  input RST,
  input init,
  input [15:0] W0A,
  input W0E,
  input [7:0] W0I,
  input [15:0] R1A,
  input R1E,
  output [7:0] R1O
);

reg [7:0] ram [65535:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 65536; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [15:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module UnbankedMem_mem_3(
  input CLK,
  input RST,
  input init,
  input [9:0] W0A,
  input W0E,
  input [18:0] W0I,
  input [9:0] R1A,
  input R1E,
  output [18:0] R1O
);

reg [18:0] ram [1023:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 1024; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [9:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module HellaFlowQueue_ram(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [132:0] W0I,
  input [5:0] R1A,
  input R1E,
  output [132:0] R1O
);

reg [132:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {5 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [6:0] RW0A,
  input RW0E,
  input RW0W,
  input [37:0] RW0M,
  input [37:0] RW0I,
  output [37:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+19) begin
    for (j=1; j<19; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [37:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {2 {$random}};
    end
  `endif
  reg [6:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][18:0] <= RW0I[18:0];
  if (RW0E && RW0W && RW0M[19]) ram[RW0A][37:19] <= RW0I[37:19];
end
assign RW0O = ram[reg_RW0A];

endmodule


module DataArray_T6(
  input CLK,
  input RST,
  input init,
  input [8:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [8:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [511:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [8:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module PacketFilter_getReqRoutes(
  input CLK,
  input RST,
  input init,
  input [3:0] W0A,
  input W0E,
  input [207:0] W0I,
  input [3:0] R1A,
  input R1E,
  output [207:0] R1O
);

reg [207:0] ram [15:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 16; initvar = initvar+1)
        ram[initvar] = {7 {$random}};
    end
  `endif
  reg [3:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module UnbankedMem_mem_1(
  input CLK,
  input RST,
  input init,
  input [15:0] W0A,
  input W0E,
  input [31:0] W0I,
  input [15:0] R1A,
  input R1E,
  output [31:0] R1O
);

reg [31:0] ram [65535:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 65536; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [15:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module UnbankedMem_mem_2(
  input CLK,
  input RST,
  input init,
  input [18:0] W0A,
  input W0E,
  input [7:0] W0I,
  input [18:0] R1A,
  input R1E,
  output [7:0] R1O
);

reg [7:0] ram [524287:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 524288; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [18:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_T156(
  input CLK,
  input RST,
  input init,
  input [8:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [511:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [8:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


module LookupPipeline_lenMem(
  input CLK,
  input RST,
  input init,
  input [9:0] W0A,
  input W0E,
  input [7:0] W0I,
  input [9:0] R1A,
  input R1E,
  output [7:0] R1O
);

reg [7:0] ram [1023:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 1024; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [9:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


