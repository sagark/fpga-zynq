module BTB(input clk, input reset,
    input  io_req_valid,
    input [42:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output[42:0] io_resp_bits_target,
    output[5:0] io_resp_bits_entry,
    output[6:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_update_valid,
    input  io_update_bits_prediction_valid,
    input  io_update_bits_prediction_bits_taken,
    input [42:0] io_update_bits_prediction_bits_target,
    input [5:0] io_update_bits_prediction_bits_entry,
    input [6:0] io_update_bits_prediction_bits_bht_history,
    input [1:0] io_update_bits_prediction_bits_bht_value,
    input [42:0] io_update_bits_pc,
    input [42:0] io_update_bits_target,
    input [42:0] io_update_bits_returnAddr,
    input  io_update_bits_taken,
    input  io_update_bits_isJump,
    input  io_update_bits_isCall,
    input  io_update_bits_isReturn,
    input  io_update_bits_mispredict,
    input  io_invalidate
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg [42:0] R4;
  wire[42:0] T5;
  wire T6;
  wire T7;
  wire updateTarget;
  reg  R8;
  wire T9;
  wire T10;
  reg  R11;
  wire T12;
  wire updateValid;
  reg  updateHit;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  R18;
  wire T1590;
  wire[1:0] T19;
  wire[1:0] T20;
  reg [1:0] T21 [127:0];
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  reg [6:0] R38;
  wire[6:0] T39;
  wire[6:0] T40;
  wire[6:0] T41;
  wire[5:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[61:0] T47;
  reg [61:0] isJump;
  wire[61:0] T1591;
  wire[63:0] T48;
  wire[63:0] T1592;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T1593;
  wire[61:0] T52;
  wire[63:0] T53;
  wire[5:0] T54;
  reg [5:0] R55;
  wire[5:0] T1594;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg [5:0] R63;
  wire[5:0] T64;
  wire[63:0] T1595;
  wire T65;
  wire T66;
  reg  R67;
  wire T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T1596;
  wire[61:0] hits;
  wire[61:0] T71;
  wire[61:0] T72;
  wire[30:0] T73;
  wire[15:0] T74;
  wire[7:0] T75;
  wire[3:0] T76;
  wire[1:0] T77;
  wire T78;
  wire[5:0] T79;
  wire[5:0] pageHit;
  reg [5:0] pageValid;
  wire[5:0] T1597;
  wire[7:0] T1598;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T1599;
  wire[7:0] T82;
  wire[7:0] pageReplEn;
  wire[7:0] tgtPageReplEn;
  wire[7:0] tgtPageRepl;
  wire[7:0] T1600;
  wire[5:0] T83;
  wire[5:0] T1601;
  wire T84;
  wire[5:0] T85;
  wire[4:0] T86;
  wire[7:0] idxPageUpdateOH;
  wire[7:0] idxPageRepl;
  wire[7:0] T87;
  reg [2:0] R88;
  wire[2:0] T1602;
  wire[2:0] T89;
  wire[2:0] T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire T94;
  wire[7:0] T1603;
  wire[5:0] updatePageHit;
  wire[5:0] T95;
  wire[5:0] T96;
  wire[2:0] T97;
  wire[1:0] T98;
  wire T99;
  wire[29:0] T100;
  reg [42:0] R101;
  wire[42:0] T102;
  wire[29:0] T103;
  reg [29:0] pages [5:0];
  wire[29:0] T104;
  wire[29:0] T105;
  wire[29:0] T106;
  wire[29:0] T107;
  wire T108;
  wire[7:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire[29:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire[29:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[29:0] T122;
  wire[29:0] T123;
  wire[29:0] T124;
  wire[29:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire[29:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[29:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[29:0] T139;
  wire T140;
  wire[29:0] T141;
  wire[2:0] T142;
  wire[1:0] T143;
  wire T144;
  wire[29:0] T145;
  wire T146;
  wire[29:0] T147;
  wire T148;
  wire[29:0] T149;
  wire useUpdatePageHit;
  wire samePage;
  wire[29:0] T150;
  wire[29:0] T151;
  wire doTgtPageRepl;
  wire T152;
  wire usePageHit;
  wire[7:0] T153;
  wire[7:0] T154;
  wire[7:0] T1604;
  wire T155;
  wire T156;
  wire[7:0] idxPageReplEn;
  wire[7:0] T1605;
  wire T157;
  wire[5:0] T158;
  wire[5:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[29:0] T163;
  wire[29:0] T164;
  wire T165;
  wire[29:0] T166;
  wire T167;
  wire[29:0] T168;
  wire[2:0] T169;
  wire[1:0] T170;
  wire T171;
  wire[29:0] T172;
  wire T173;
  wire[29:0] T174;
  wire T175;
  wire[29:0] T176;
  wire[5:0] idxPagesOH_0;
  wire[7:0] T177;
  wire[2:0] T178;
  reg [2:0] idxPages [61:0];
  wire[2:0] T179;
  wire[2:0] T1606;
  wire[1:0] T1607;
  wire T1608;
  wire[1:0] T1609;
  wire[1:0] T1610;
  wire[3:0] T1611;
  wire[3:0] T1612;
  wire[3:0] T1613;
  wire[1:0] T1614;
  wire T1615;
  wire T1616;
  wire T180;
  wire T181;
  wire T182;
  wire[5:0] T183;
  wire[5:0] idxPagesOH_1;
  wire[7:0] T184;
  wire[2:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[5:0] T188;
  wire[5:0] idxPagesOH_2;
  wire[7:0] T189;
  wire[2:0] T190;
  wire T191;
  wire[5:0] T192;
  wire[5:0] idxPagesOH_3;
  wire[7:0] T193;
  wire[2:0] T194;
  wire[3:0] T195;
  wire[1:0] T196;
  wire T197;
  wire[5:0] T198;
  wire[5:0] idxPagesOH_4;
  wire[7:0] T199;
  wire[2:0] T200;
  wire T201;
  wire[5:0] T202;
  wire[5:0] idxPagesOH_5;
  wire[7:0] T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[5:0] T207;
  wire[5:0] idxPagesOH_6;
  wire[7:0] T208;
  wire[2:0] T209;
  wire T210;
  wire[5:0] T211;
  wire[5:0] idxPagesOH_7;
  wire[7:0] T212;
  wire[2:0] T213;
  wire[7:0] T214;
  wire[3:0] T215;
  wire[1:0] T216;
  wire T217;
  wire[5:0] T218;
  wire[5:0] idxPagesOH_8;
  wire[7:0] T219;
  wire[2:0] T220;
  wire T221;
  wire[5:0] T222;
  wire[5:0] idxPagesOH_9;
  wire[7:0] T223;
  wire[2:0] T224;
  wire[1:0] T225;
  wire T226;
  wire[5:0] T227;
  wire[5:0] idxPagesOH_10;
  wire[7:0] T228;
  wire[2:0] T229;
  wire T230;
  wire[5:0] T231;
  wire[5:0] idxPagesOH_11;
  wire[7:0] T232;
  wire[2:0] T233;
  wire[3:0] T234;
  wire[1:0] T235;
  wire T236;
  wire[5:0] T237;
  wire[5:0] idxPagesOH_12;
  wire[7:0] T238;
  wire[2:0] T239;
  wire T240;
  wire[5:0] T241;
  wire[5:0] idxPagesOH_13;
  wire[7:0] T242;
  wire[2:0] T243;
  wire[1:0] T244;
  wire T245;
  wire[5:0] T246;
  wire[5:0] idxPagesOH_14;
  wire[7:0] T247;
  wire[2:0] T248;
  wire T249;
  wire[5:0] T250;
  wire[5:0] idxPagesOH_15;
  wire[7:0] T251;
  wire[2:0] T252;
  wire[14:0] T253;
  wire[7:0] T254;
  wire[3:0] T255;
  wire[1:0] T256;
  wire T257;
  wire[5:0] T258;
  wire[5:0] idxPagesOH_16;
  wire[7:0] T259;
  wire[2:0] T260;
  wire T261;
  wire[5:0] T262;
  wire[5:0] idxPagesOH_17;
  wire[7:0] T263;
  wire[2:0] T264;
  wire[1:0] T265;
  wire T266;
  wire[5:0] T267;
  wire[5:0] idxPagesOH_18;
  wire[7:0] T268;
  wire[2:0] T269;
  wire T270;
  wire[5:0] T271;
  wire[5:0] idxPagesOH_19;
  wire[7:0] T272;
  wire[2:0] T273;
  wire[3:0] T274;
  wire[1:0] T275;
  wire T276;
  wire[5:0] T277;
  wire[5:0] idxPagesOH_20;
  wire[7:0] T278;
  wire[2:0] T279;
  wire T280;
  wire[5:0] T281;
  wire[5:0] idxPagesOH_21;
  wire[7:0] T282;
  wire[2:0] T283;
  wire[1:0] T284;
  wire T285;
  wire[5:0] T286;
  wire[5:0] idxPagesOH_22;
  wire[7:0] T287;
  wire[2:0] T288;
  wire T289;
  wire[5:0] T290;
  wire[5:0] idxPagesOH_23;
  wire[7:0] T291;
  wire[2:0] T292;
  wire[6:0] T293;
  wire[3:0] T294;
  wire[1:0] T295;
  wire T296;
  wire[5:0] T297;
  wire[5:0] idxPagesOH_24;
  wire[7:0] T298;
  wire[2:0] T299;
  wire T300;
  wire[5:0] T301;
  wire[5:0] idxPagesOH_25;
  wire[7:0] T302;
  wire[2:0] T303;
  wire[1:0] T304;
  wire T305;
  wire[5:0] T306;
  wire[5:0] idxPagesOH_26;
  wire[7:0] T307;
  wire[2:0] T308;
  wire T309;
  wire[5:0] T310;
  wire[5:0] idxPagesOH_27;
  wire[7:0] T311;
  wire[2:0] T312;
  wire[2:0] T313;
  wire[1:0] T314;
  wire T315;
  wire[5:0] T316;
  wire[5:0] idxPagesOH_28;
  wire[7:0] T317;
  wire[2:0] T318;
  wire T319;
  wire[5:0] T320;
  wire[5:0] idxPagesOH_29;
  wire[7:0] T321;
  wire[2:0] T322;
  wire T323;
  wire[5:0] T324;
  wire[5:0] idxPagesOH_30;
  wire[7:0] T325;
  wire[2:0] T326;
  wire[30:0] T327;
  wire[15:0] T328;
  wire[7:0] T329;
  wire[3:0] T330;
  wire[1:0] T331;
  wire T332;
  wire[5:0] T333;
  wire[5:0] idxPagesOH_31;
  wire[7:0] T334;
  wire[2:0] T335;
  wire T336;
  wire[5:0] T337;
  wire[5:0] idxPagesOH_32;
  wire[7:0] T338;
  wire[2:0] T339;
  wire[1:0] T340;
  wire T341;
  wire[5:0] T342;
  wire[5:0] idxPagesOH_33;
  wire[7:0] T343;
  wire[2:0] T344;
  wire T345;
  wire[5:0] T346;
  wire[5:0] idxPagesOH_34;
  wire[7:0] T347;
  wire[2:0] T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire T351;
  wire[5:0] T352;
  wire[5:0] idxPagesOH_35;
  wire[7:0] T353;
  wire[2:0] T354;
  wire T355;
  wire[5:0] T356;
  wire[5:0] idxPagesOH_36;
  wire[7:0] T357;
  wire[2:0] T358;
  wire[1:0] T359;
  wire T360;
  wire[5:0] T361;
  wire[5:0] idxPagesOH_37;
  wire[7:0] T362;
  wire[2:0] T363;
  wire T364;
  wire[5:0] T365;
  wire[5:0] idxPagesOH_38;
  wire[7:0] T366;
  wire[2:0] T367;
  wire[7:0] T368;
  wire[3:0] T369;
  wire[1:0] T370;
  wire T371;
  wire[5:0] T372;
  wire[5:0] idxPagesOH_39;
  wire[7:0] T373;
  wire[2:0] T374;
  wire T375;
  wire[5:0] T376;
  wire[5:0] idxPagesOH_40;
  wire[7:0] T377;
  wire[2:0] T378;
  wire[1:0] T379;
  wire T380;
  wire[5:0] T381;
  wire[5:0] idxPagesOH_41;
  wire[7:0] T382;
  wire[2:0] T383;
  wire T384;
  wire[5:0] T385;
  wire[5:0] idxPagesOH_42;
  wire[7:0] T386;
  wire[2:0] T387;
  wire[3:0] T388;
  wire[1:0] T389;
  wire T390;
  wire[5:0] T391;
  wire[5:0] idxPagesOH_43;
  wire[7:0] T392;
  wire[2:0] T393;
  wire T394;
  wire[5:0] T395;
  wire[5:0] idxPagesOH_44;
  wire[7:0] T396;
  wire[2:0] T397;
  wire[1:0] T398;
  wire T399;
  wire[5:0] T400;
  wire[5:0] idxPagesOH_45;
  wire[7:0] T401;
  wire[2:0] T402;
  wire T403;
  wire[5:0] T404;
  wire[5:0] idxPagesOH_46;
  wire[7:0] T405;
  wire[2:0] T406;
  wire[14:0] T407;
  wire[7:0] T408;
  wire[3:0] T409;
  wire[1:0] T410;
  wire T411;
  wire[5:0] T412;
  wire[5:0] idxPagesOH_47;
  wire[7:0] T413;
  wire[2:0] T414;
  wire T415;
  wire[5:0] T416;
  wire[5:0] idxPagesOH_48;
  wire[7:0] T417;
  wire[2:0] T418;
  wire[1:0] T419;
  wire T420;
  wire[5:0] T421;
  wire[5:0] idxPagesOH_49;
  wire[7:0] T422;
  wire[2:0] T423;
  wire T424;
  wire[5:0] T425;
  wire[5:0] idxPagesOH_50;
  wire[7:0] T426;
  wire[2:0] T427;
  wire[3:0] T428;
  wire[1:0] T429;
  wire T430;
  wire[5:0] T431;
  wire[5:0] idxPagesOH_51;
  wire[7:0] T432;
  wire[2:0] T433;
  wire T434;
  wire[5:0] T435;
  wire[5:0] idxPagesOH_52;
  wire[7:0] T436;
  wire[2:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[5:0] T440;
  wire[5:0] idxPagesOH_53;
  wire[7:0] T441;
  wire[2:0] T442;
  wire T443;
  wire[5:0] T444;
  wire[5:0] idxPagesOH_54;
  wire[7:0] T445;
  wire[2:0] T446;
  wire[6:0] T447;
  wire[3:0] T448;
  wire[1:0] T449;
  wire T450;
  wire[5:0] T451;
  wire[5:0] idxPagesOH_55;
  wire[7:0] T452;
  wire[2:0] T453;
  wire T454;
  wire[5:0] T455;
  wire[5:0] idxPagesOH_56;
  wire[7:0] T456;
  wire[2:0] T457;
  wire[1:0] T458;
  wire T459;
  wire[5:0] T460;
  wire[5:0] idxPagesOH_57;
  wire[7:0] T461;
  wire[2:0] T462;
  wire T463;
  wire[5:0] T464;
  wire[5:0] idxPagesOH_58;
  wire[7:0] T465;
  wire[2:0] T466;
  wire[2:0] T467;
  wire[1:0] T468;
  wire T469;
  wire[5:0] T470;
  wire[5:0] idxPagesOH_59;
  wire[7:0] T471;
  wire[2:0] T472;
  wire T473;
  wire[5:0] T474;
  wire[5:0] idxPagesOH_60;
  wire[7:0] T475;
  wire[2:0] T476;
  wire T477;
  wire[5:0] T478;
  wire[5:0] idxPagesOH_61;
  wire[7:0] T479;
  wire[2:0] T480;
  wire[61:0] T481;
  wire[61:0] T482;
  wire[61:0] T483;
  wire[30:0] T484;
  wire[15:0] T485;
  wire[7:0] T486;
  wire[3:0] T487;
  wire[1:0] T488;
  wire T489;
  wire[12:0] T490;
  wire[12:0] T491;
  reg [12:0] idxs [61:0];
  wire[12:0] T492;
  wire[12:0] T1617;
  wire T493;
  wire T494;
  wire T495;
  wire[12:0] T496;
  wire[1:0] T497;
  wire T498;
  wire[12:0] T499;
  wire T500;
  wire[12:0] T501;
  wire[3:0] T502;
  wire[1:0] T503;
  wire T504;
  wire[12:0] T505;
  wire T506;
  wire[12:0] T507;
  wire[1:0] T508;
  wire T509;
  wire[12:0] T510;
  wire T511;
  wire[12:0] T512;
  wire[7:0] T513;
  wire[3:0] T514;
  wire[1:0] T515;
  wire T516;
  wire[12:0] T517;
  wire T518;
  wire[12:0] T519;
  wire[1:0] T520;
  wire T521;
  wire[12:0] T522;
  wire T523;
  wire[12:0] T524;
  wire[3:0] T525;
  wire[1:0] T526;
  wire T527;
  wire[12:0] T528;
  wire T529;
  wire[12:0] T530;
  wire[1:0] T531;
  wire T532;
  wire[12:0] T533;
  wire T534;
  wire[12:0] T535;
  wire[14:0] T536;
  wire[7:0] T537;
  wire[3:0] T538;
  wire[1:0] T539;
  wire T540;
  wire[12:0] T541;
  wire T542;
  wire[12:0] T543;
  wire[1:0] T544;
  wire T545;
  wire[12:0] T546;
  wire T547;
  wire[12:0] T548;
  wire[3:0] T549;
  wire[1:0] T550;
  wire T551;
  wire[12:0] T552;
  wire T553;
  wire[12:0] T554;
  wire[1:0] T555;
  wire T556;
  wire[12:0] T557;
  wire T558;
  wire[12:0] T559;
  wire[6:0] T560;
  wire[3:0] T561;
  wire[1:0] T562;
  wire T563;
  wire[12:0] T564;
  wire T565;
  wire[12:0] T566;
  wire[1:0] T567;
  wire T568;
  wire[12:0] T569;
  wire T570;
  wire[12:0] T571;
  wire[2:0] T572;
  wire[1:0] T573;
  wire T574;
  wire[12:0] T575;
  wire T576;
  wire[12:0] T577;
  wire T578;
  wire[12:0] T579;
  wire[30:0] T580;
  wire[15:0] T581;
  wire[7:0] T582;
  wire[3:0] T583;
  wire[1:0] T584;
  wire T585;
  wire[12:0] T586;
  wire T587;
  wire[12:0] T588;
  wire[1:0] T589;
  wire T590;
  wire[12:0] T591;
  wire T592;
  wire[12:0] T593;
  wire[3:0] T594;
  wire[1:0] T595;
  wire T596;
  wire[12:0] T597;
  wire T598;
  wire[12:0] T599;
  wire[1:0] T600;
  wire T601;
  wire[12:0] T602;
  wire T603;
  wire[12:0] T604;
  wire[7:0] T605;
  wire[3:0] T606;
  wire[1:0] T607;
  wire T608;
  wire[12:0] T609;
  wire T610;
  wire[12:0] T611;
  wire[1:0] T612;
  wire T613;
  wire[12:0] T614;
  wire T615;
  wire[12:0] T616;
  wire[3:0] T617;
  wire[1:0] T618;
  wire T619;
  wire[12:0] T620;
  wire T621;
  wire[12:0] T622;
  wire[1:0] T623;
  wire T624;
  wire[12:0] T625;
  wire T626;
  wire[12:0] T627;
  wire[14:0] T628;
  wire[7:0] T629;
  wire[3:0] T630;
  wire[1:0] T631;
  wire T632;
  wire[12:0] T633;
  wire T634;
  wire[12:0] T635;
  wire[1:0] T636;
  wire T637;
  wire[12:0] T638;
  wire T639;
  wire[12:0] T640;
  wire[3:0] T641;
  wire[1:0] T642;
  wire T643;
  wire[12:0] T644;
  wire T645;
  wire[12:0] T646;
  wire[1:0] T647;
  wire T648;
  wire[12:0] T649;
  wire T650;
  wire[12:0] T651;
  wire[6:0] T652;
  wire[3:0] T653;
  wire[1:0] T654;
  wire T655;
  wire[12:0] T656;
  wire T657;
  wire[12:0] T658;
  wire[1:0] T659;
  wire T660;
  wire[12:0] T661;
  wire T662;
  wire[12:0] T663;
  wire[2:0] T664;
  wire[1:0] T665;
  wire T666;
  wire[12:0] T667;
  wire T668;
  wire[12:0] T669;
  wire T670;
  wire[12:0] T671;
  reg [61:0] idxValid;
  wire[61:0] T1618;
  wire[63:0] T1619;
  wire[63:0] T672;
  wire[63:0] T673;
  wire[63:0] T1620;
  wire[61:0] T674;
  wire[61:0] T675;
  wire[61:0] T676;
  wire[61:0] T677;
  wire[61:0] T678;
  wire[30:0] T679;
  wire[15:0] T680;
  wire[7:0] T681;
  wire[3:0] T682;
  wire[1:0] T683;
  wire T684;
  wire[7:0] T685;
  wire[7:0] T1621;
  wire[5:0] T686;
  wire[5:0] tgtPagesOH_0;
  wire[7:0] T687;
  wire[2:0] T688;
  reg [2:0] tgtPages [61:0];
  wire[2:0] T689;
  wire[2:0] T1622;
  wire[1:0] T1623;
  wire T1624;
  wire[1:0] T1625;
  wire[1:0] T1626;
  wire[3:0] T1627;
  wire[3:0] T1628;
  wire[7:0] T690;
  wire[7:0] T1629;
  wire[3:0] T1630;
  wire[1:0] T1631;
  wire T1632;
  wire T1633;
  wire T691;
  wire T692;
  wire T693;
  wire[7:0] T694;
  wire[7:0] T1634;
  wire[5:0] T695;
  wire[5:0] tgtPagesOH_1;
  wire[7:0] T696;
  wire[2:0] T697;
  wire[1:0] T698;
  wire T699;
  wire[7:0] T700;
  wire[7:0] T1635;
  wire[5:0] T701;
  wire[5:0] tgtPagesOH_2;
  wire[7:0] T702;
  wire[2:0] T703;
  wire T704;
  wire[7:0] T705;
  wire[7:0] T1636;
  wire[5:0] T706;
  wire[5:0] tgtPagesOH_3;
  wire[7:0] T707;
  wire[2:0] T708;
  wire[3:0] T709;
  wire[1:0] T710;
  wire T711;
  wire[7:0] T712;
  wire[7:0] T1637;
  wire[5:0] T713;
  wire[5:0] tgtPagesOH_4;
  wire[7:0] T714;
  wire[2:0] T715;
  wire T716;
  wire[7:0] T717;
  wire[7:0] T1638;
  wire[5:0] T718;
  wire[5:0] tgtPagesOH_5;
  wire[7:0] T719;
  wire[2:0] T720;
  wire[1:0] T721;
  wire T722;
  wire[7:0] T723;
  wire[7:0] T1639;
  wire[5:0] T724;
  wire[5:0] tgtPagesOH_6;
  wire[7:0] T725;
  wire[2:0] T726;
  wire T727;
  wire[7:0] T728;
  wire[7:0] T1640;
  wire[5:0] T729;
  wire[5:0] tgtPagesOH_7;
  wire[7:0] T730;
  wire[2:0] T731;
  wire[7:0] T732;
  wire[3:0] T733;
  wire[1:0] T734;
  wire T735;
  wire[7:0] T736;
  wire[7:0] T1641;
  wire[5:0] T737;
  wire[5:0] tgtPagesOH_8;
  wire[7:0] T738;
  wire[2:0] T739;
  wire T740;
  wire[7:0] T741;
  wire[7:0] T1642;
  wire[5:0] T742;
  wire[5:0] tgtPagesOH_9;
  wire[7:0] T743;
  wire[2:0] T744;
  wire[1:0] T745;
  wire T746;
  wire[7:0] T747;
  wire[7:0] T1643;
  wire[5:0] T748;
  wire[5:0] tgtPagesOH_10;
  wire[7:0] T749;
  wire[2:0] T750;
  wire T751;
  wire[7:0] T752;
  wire[7:0] T1644;
  wire[5:0] T753;
  wire[5:0] tgtPagesOH_11;
  wire[7:0] T754;
  wire[2:0] T755;
  wire[3:0] T756;
  wire[1:0] T757;
  wire T758;
  wire[7:0] T759;
  wire[7:0] T1645;
  wire[5:0] T760;
  wire[5:0] tgtPagesOH_12;
  wire[7:0] T761;
  wire[2:0] T762;
  wire T763;
  wire[7:0] T764;
  wire[7:0] T1646;
  wire[5:0] T765;
  wire[5:0] tgtPagesOH_13;
  wire[7:0] T766;
  wire[2:0] T767;
  wire[1:0] T768;
  wire T769;
  wire[7:0] T770;
  wire[7:0] T1647;
  wire[5:0] T771;
  wire[5:0] tgtPagesOH_14;
  wire[7:0] T772;
  wire[2:0] T773;
  wire T774;
  wire[7:0] T775;
  wire[7:0] T1648;
  wire[5:0] T776;
  wire[5:0] tgtPagesOH_15;
  wire[7:0] T777;
  wire[2:0] T778;
  wire[14:0] T779;
  wire[7:0] T780;
  wire[3:0] T781;
  wire[1:0] T782;
  wire T783;
  wire[7:0] T784;
  wire[7:0] T1649;
  wire[5:0] T785;
  wire[5:0] tgtPagesOH_16;
  wire[7:0] T786;
  wire[2:0] T787;
  wire T788;
  wire[7:0] T789;
  wire[7:0] T1650;
  wire[5:0] T790;
  wire[5:0] tgtPagesOH_17;
  wire[7:0] T791;
  wire[2:0] T792;
  wire[1:0] T793;
  wire T794;
  wire[7:0] T795;
  wire[7:0] T1651;
  wire[5:0] T796;
  wire[5:0] tgtPagesOH_18;
  wire[7:0] T797;
  wire[2:0] T798;
  wire T799;
  wire[7:0] T800;
  wire[7:0] T1652;
  wire[5:0] T801;
  wire[5:0] tgtPagesOH_19;
  wire[7:0] T802;
  wire[2:0] T803;
  wire[3:0] T804;
  wire[1:0] T805;
  wire T806;
  wire[7:0] T807;
  wire[7:0] T1653;
  wire[5:0] T808;
  wire[5:0] tgtPagesOH_20;
  wire[7:0] T809;
  wire[2:0] T810;
  wire T811;
  wire[7:0] T812;
  wire[7:0] T1654;
  wire[5:0] T813;
  wire[5:0] tgtPagesOH_21;
  wire[7:0] T814;
  wire[2:0] T815;
  wire[1:0] T816;
  wire T817;
  wire[7:0] T818;
  wire[7:0] T1655;
  wire[5:0] T819;
  wire[5:0] tgtPagesOH_22;
  wire[7:0] T820;
  wire[2:0] T821;
  wire T822;
  wire[7:0] T823;
  wire[7:0] T1656;
  wire[5:0] T824;
  wire[5:0] tgtPagesOH_23;
  wire[7:0] T825;
  wire[2:0] T826;
  wire[6:0] T827;
  wire[3:0] T828;
  wire[1:0] T829;
  wire T830;
  wire[7:0] T831;
  wire[7:0] T1657;
  wire[5:0] T832;
  wire[5:0] tgtPagesOH_24;
  wire[7:0] T833;
  wire[2:0] T834;
  wire T835;
  wire[7:0] T836;
  wire[7:0] T1658;
  wire[5:0] T837;
  wire[5:0] tgtPagesOH_25;
  wire[7:0] T838;
  wire[2:0] T839;
  wire[1:0] T840;
  wire T841;
  wire[7:0] T842;
  wire[7:0] T1659;
  wire[5:0] T843;
  wire[5:0] tgtPagesOH_26;
  wire[7:0] T844;
  wire[2:0] T845;
  wire T846;
  wire[7:0] T847;
  wire[7:0] T1660;
  wire[5:0] T848;
  wire[5:0] tgtPagesOH_27;
  wire[7:0] T849;
  wire[2:0] T850;
  wire[2:0] T851;
  wire[1:0] T852;
  wire T853;
  wire[7:0] T854;
  wire[7:0] T1661;
  wire[5:0] T855;
  wire[5:0] tgtPagesOH_28;
  wire[7:0] T856;
  wire[2:0] T857;
  wire T858;
  wire[7:0] T859;
  wire[7:0] T1662;
  wire[5:0] T860;
  wire[5:0] tgtPagesOH_29;
  wire[7:0] T861;
  wire[2:0] T862;
  wire T863;
  wire[7:0] T864;
  wire[7:0] T1663;
  wire[5:0] T865;
  wire[5:0] tgtPagesOH_30;
  wire[7:0] T866;
  wire[2:0] T867;
  wire[30:0] T868;
  wire[15:0] T869;
  wire[7:0] T870;
  wire[3:0] T871;
  wire[1:0] T872;
  wire T873;
  wire[7:0] T874;
  wire[7:0] T1664;
  wire[5:0] T875;
  wire[5:0] tgtPagesOH_31;
  wire[7:0] T876;
  wire[2:0] T877;
  wire T878;
  wire[7:0] T879;
  wire[7:0] T1665;
  wire[5:0] T880;
  wire[5:0] tgtPagesOH_32;
  wire[7:0] T881;
  wire[2:0] T882;
  wire[1:0] T883;
  wire T884;
  wire[7:0] T885;
  wire[7:0] T1666;
  wire[5:0] T886;
  wire[5:0] tgtPagesOH_33;
  wire[7:0] T887;
  wire[2:0] T888;
  wire T889;
  wire[7:0] T890;
  wire[7:0] T1667;
  wire[5:0] T891;
  wire[5:0] tgtPagesOH_34;
  wire[7:0] T892;
  wire[2:0] T893;
  wire[3:0] T894;
  wire[1:0] T895;
  wire T896;
  wire[7:0] T897;
  wire[7:0] T1668;
  wire[5:0] T898;
  wire[5:0] tgtPagesOH_35;
  wire[7:0] T899;
  wire[2:0] T900;
  wire T901;
  wire[7:0] T902;
  wire[7:0] T1669;
  wire[5:0] T903;
  wire[5:0] tgtPagesOH_36;
  wire[7:0] T904;
  wire[2:0] T905;
  wire[1:0] T906;
  wire T907;
  wire[7:0] T908;
  wire[7:0] T1670;
  wire[5:0] T909;
  wire[5:0] tgtPagesOH_37;
  wire[7:0] T910;
  wire[2:0] T911;
  wire T912;
  wire[7:0] T913;
  wire[7:0] T1671;
  wire[5:0] T914;
  wire[5:0] tgtPagesOH_38;
  wire[7:0] T915;
  wire[2:0] T916;
  wire[7:0] T917;
  wire[3:0] T918;
  wire[1:0] T919;
  wire T920;
  wire[7:0] T921;
  wire[7:0] T1672;
  wire[5:0] T922;
  wire[5:0] tgtPagesOH_39;
  wire[7:0] T923;
  wire[2:0] T924;
  wire T925;
  wire[7:0] T926;
  wire[7:0] T1673;
  wire[5:0] T927;
  wire[5:0] tgtPagesOH_40;
  wire[7:0] T928;
  wire[2:0] T929;
  wire[1:0] T930;
  wire T931;
  wire[7:0] T932;
  wire[7:0] T1674;
  wire[5:0] T933;
  wire[5:0] tgtPagesOH_41;
  wire[7:0] T934;
  wire[2:0] T935;
  wire T936;
  wire[7:0] T937;
  wire[7:0] T1675;
  wire[5:0] T938;
  wire[5:0] tgtPagesOH_42;
  wire[7:0] T939;
  wire[2:0] T940;
  wire[3:0] T941;
  wire[1:0] T942;
  wire T943;
  wire[7:0] T944;
  wire[7:0] T1676;
  wire[5:0] T945;
  wire[5:0] tgtPagesOH_43;
  wire[7:0] T946;
  wire[2:0] T947;
  wire T948;
  wire[7:0] T949;
  wire[7:0] T1677;
  wire[5:0] T950;
  wire[5:0] tgtPagesOH_44;
  wire[7:0] T951;
  wire[2:0] T952;
  wire[1:0] T953;
  wire T954;
  wire[7:0] T955;
  wire[7:0] T1678;
  wire[5:0] T956;
  wire[5:0] tgtPagesOH_45;
  wire[7:0] T957;
  wire[2:0] T958;
  wire T959;
  wire[7:0] T960;
  wire[7:0] T1679;
  wire[5:0] T961;
  wire[5:0] tgtPagesOH_46;
  wire[7:0] T962;
  wire[2:0] T963;
  wire[14:0] T964;
  wire[7:0] T965;
  wire[3:0] T966;
  wire[1:0] T967;
  wire T968;
  wire[7:0] T969;
  wire[7:0] T1680;
  wire[5:0] T970;
  wire[5:0] tgtPagesOH_47;
  wire[7:0] T971;
  wire[2:0] T972;
  wire T973;
  wire[7:0] T974;
  wire[7:0] T1681;
  wire[5:0] T975;
  wire[5:0] tgtPagesOH_48;
  wire[7:0] T976;
  wire[2:0] T977;
  wire[1:0] T978;
  wire T979;
  wire[7:0] T980;
  wire[7:0] T1682;
  wire[5:0] T981;
  wire[5:0] tgtPagesOH_49;
  wire[7:0] T982;
  wire[2:0] T983;
  wire T984;
  wire[7:0] T985;
  wire[7:0] T1683;
  wire[5:0] T986;
  wire[5:0] tgtPagesOH_50;
  wire[7:0] T987;
  wire[2:0] T988;
  wire[3:0] T989;
  wire[1:0] T990;
  wire T991;
  wire[7:0] T992;
  wire[7:0] T1684;
  wire[5:0] T993;
  wire[5:0] tgtPagesOH_51;
  wire[7:0] T994;
  wire[2:0] T995;
  wire T996;
  wire[7:0] T997;
  wire[7:0] T1685;
  wire[5:0] T998;
  wire[5:0] tgtPagesOH_52;
  wire[7:0] T999;
  wire[2:0] T1000;
  wire[1:0] T1001;
  wire T1002;
  wire[7:0] T1003;
  wire[7:0] T1686;
  wire[5:0] T1004;
  wire[5:0] tgtPagesOH_53;
  wire[7:0] T1005;
  wire[2:0] T1006;
  wire T1007;
  wire[7:0] T1008;
  wire[7:0] T1687;
  wire[5:0] T1009;
  wire[5:0] tgtPagesOH_54;
  wire[7:0] T1010;
  wire[2:0] T1011;
  wire[6:0] T1012;
  wire[3:0] T1013;
  wire[1:0] T1014;
  wire T1015;
  wire[7:0] T1016;
  wire[7:0] T1688;
  wire[5:0] T1017;
  wire[5:0] tgtPagesOH_55;
  wire[7:0] T1018;
  wire[2:0] T1019;
  wire T1020;
  wire[7:0] T1021;
  wire[7:0] T1689;
  wire[5:0] T1022;
  wire[5:0] tgtPagesOH_56;
  wire[7:0] T1023;
  wire[2:0] T1024;
  wire[1:0] T1025;
  wire T1026;
  wire[7:0] T1027;
  wire[7:0] T1690;
  wire[5:0] T1028;
  wire[5:0] tgtPagesOH_57;
  wire[7:0] T1029;
  wire[2:0] T1030;
  wire T1031;
  wire[7:0] T1032;
  wire[7:0] T1691;
  wire[5:0] T1033;
  wire[5:0] tgtPagesOH_58;
  wire[7:0] T1034;
  wire[2:0] T1035;
  wire[2:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire[7:0] T1039;
  wire[7:0] T1692;
  wire[5:0] T1040;
  wire[5:0] tgtPagesOH_59;
  wire[7:0] T1041;
  wire[2:0] T1042;
  wire T1043;
  wire[7:0] T1044;
  wire[7:0] T1693;
  wire[5:0] T1045;
  wire[5:0] tgtPagesOH_60;
  wire[7:0] T1046;
  wire[2:0] T1047;
  wire T1048;
  wire[7:0] T1049;
  wire[7:0] T1694;
  wire[5:0] T1050;
  wire[5:0] tgtPagesOH_61;
  wire[7:0] T1051;
  wire[2:0] T1052;
  wire[63:0] T1053;
  wire[63:0] T1054;
  wire[63:0] T1055;
  wire[63:0] T1695;
  wire[61:0] T1056;
  wire[63:0] T1057;
  wire[63:0] T1696;
  wire T1058;
  wire T1059;
  wire[63:0] T1060;
  wire[63:0] T1061;
  wire[63:0] T1697;
  wire T1062;
  wire T1063;
  wire[6:0] T1064;
  wire[5:0] T1065;
  wire T1066;
  wire[6:0] T1067;
  wire[6:0] T1068;
  wire[5:0] T1698;
  wire[4:0] T1699;
  wire[3:0] T1700;
  wire[2:0] T1701;
  wire[1:0] T1702;
  wire T1703;
  wire[1:0] T1704;
  wire[1:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[7:0] T1708;
  wire[7:0] T1709;
  wire[15:0] T1710;
  wire[15:0] T1711;
  wire[31:0] T1712;
  wire[31:0] T1713;
  wire[29:0] T1714;
  wire[15:0] T1715;
  wire[7:0] T1716;
  wire[3:0] T1717;
  wire[1:0] T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire T1723;
  wire[42:0] T1070;
  wire[42:0] T1071;
  wire[42:0] T1072;
  wire[12:0] T1073;
  wire[12:0] T1074;
  wire[12:0] T1075;
  reg [12:0] tgts [61:0];
  wire[12:0] T1076;
  wire[12:0] T1724;
  wire T1077;
  wire T1078;
  wire T1079;
  wire[12:0] T1080;
  wire[12:0] T1081;
  wire[12:0] T1082;
  wire T1083;
  wire[12:0] T1084;
  wire[12:0] T1085;
  wire[12:0] T1086;
  wire T1087;
  wire[12:0] T1088;
  wire[12:0] T1089;
  wire[12:0] T1090;
  wire T1091;
  wire[12:0] T1092;
  wire[12:0] T1093;
  wire[12:0] T1094;
  wire T1095;
  wire[12:0] T1096;
  wire[12:0] T1097;
  wire[12:0] T1098;
  wire T1099;
  wire[12:0] T1100;
  wire[12:0] T1101;
  wire[12:0] T1102;
  wire T1103;
  wire[12:0] T1104;
  wire[12:0] T1105;
  wire[12:0] T1106;
  wire T1107;
  wire[12:0] T1108;
  wire[12:0] T1109;
  wire[12:0] T1110;
  wire T1111;
  wire[12:0] T1112;
  wire[12:0] T1113;
  wire[12:0] T1114;
  wire T1115;
  wire[12:0] T1116;
  wire[12:0] T1117;
  wire[12:0] T1118;
  wire T1119;
  wire[12:0] T1120;
  wire[12:0] T1121;
  wire[12:0] T1122;
  wire T1123;
  wire[12:0] T1124;
  wire[12:0] T1125;
  wire[12:0] T1126;
  wire T1127;
  wire[12:0] T1128;
  wire[12:0] T1129;
  wire[12:0] T1130;
  wire T1131;
  wire[12:0] T1132;
  wire[12:0] T1133;
  wire[12:0] T1134;
  wire T1135;
  wire[12:0] T1136;
  wire[12:0] T1137;
  wire[12:0] T1138;
  wire T1139;
  wire[12:0] T1140;
  wire[12:0] T1141;
  wire[12:0] T1142;
  wire T1143;
  wire[12:0] T1144;
  wire[12:0] T1145;
  wire[12:0] T1146;
  wire T1147;
  wire[12:0] T1148;
  wire[12:0] T1149;
  wire[12:0] T1150;
  wire T1151;
  wire[12:0] T1152;
  wire[12:0] T1153;
  wire[12:0] T1154;
  wire T1155;
  wire[12:0] T1156;
  wire[12:0] T1157;
  wire[12:0] T1158;
  wire T1159;
  wire[12:0] T1160;
  wire[12:0] T1161;
  wire[12:0] T1162;
  wire T1163;
  wire[12:0] T1164;
  wire[12:0] T1165;
  wire[12:0] T1166;
  wire T1167;
  wire[12:0] T1168;
  wire[12:0] T1169;
  wire[12:0] T1170;
  wire T1171;
  wire[12:0] T1172;
  wire[12:0] T1173;
  wire[12:0] T1174;
  wire T1175;
  wire[12:0] T1176;
  wire[12:0] T1177;
  wire[12:0] T1178;
  wire T1179;
  wire[12:0] T1180;
  wire[12:0] T1181;
  wire[12:0] T1182;
  wire T1183;
  wire[12:0] T1184;
  wire[12:0] T1185;
  wire[12:0] T1186;
  wire T1187;
  wire[12:0] T1188;
  wire[12:0] T1189;
  wire[12:0] T1190;
  wire T1191;
  wire[12:0] T1192;
  wire[12:0] T1193;
  wire[12:0] T1194;
  wire T1195;
  wire[12:0] T1196;
  wire[12:0] T1197;
  wire[12:0] T1198;
  wire T1199;
  wire[12:0] T1200;
  wire[12:0] T1201;
  wire[12:0] T1202;
  wire T1203;
  wire[12:0] T1204;
  wire[12:0] T1205;
  wire[12:0] T1206;
  wire T1207;
  wire[12:0] T1208;
  wire[12:0] T1209;
  wire[12:0] T1210;
  wire T1211;
  wire[12:0] T1212;
  wire[12:0] T1213;
  wire[12:0] T1214;
  wire T1215;
  wire[12:0] T1216;
  wire[12:0] T1217;
  wire[12:0] T1218;
  wire T1219;
  wire[12:0] T1220;
  wire[12:0] T1221;
  wire[12:0] T1222;
  wire T1223;
  wire[12:0] T1224;
  wire[12:0] T1225;
  wire[12:0] T1226;
  wire T1227;
  wire[12:0] T1228;
  wire[12:0] T1229;
  wire[12:0] T1230;
  wire T1231;
  wire[12:0] T1232;
  wire[12:0] T1233;
  wire[12:0] T1234;
  wire T1235;
  wire[12:0] T1236;
  wire[12:0] T1237;
  wire[12:0] T1238;
  wire T1239;
  wire[12:0] T1240;
  wire[12:0] T1241;
  wire[12:0] T1242;
  wire T1243;
  wire[12:0] T1244;
  wire[12:0] T1245;
  wire[12:0] T1246;
  wire T1247;
  wire[12:0] T1248;
  wire[12:0] T1249;
  wire[12:0] T1250;
  wire T1251;
  wire[12:0] T1252;
  wire[12:0] T1253;
  wire[12:0] T1254;
  wire T1255;
  wire[12:0] T1256;
  wire[12:0] T1257;
  wire[12:0] T1258;
  wire T1259;
  wire[12:0] T1260;
  wire[12:0] T1261;
  wire[12:0] T1262;
  wire T1263;
  wire[12:0] T1264;
  wire[12:0] T1265;
  wire[12:0] T1266;
  wire T1267;
  wire[12:0] T1268;
  wire[12:0] T1269;
  wire[12:0] T1270;
  wire T1271;
  wire[12:0] T1272;
  wire[12:0] T1273;
  wire[12:0] T1274;
  wire T1275;
  wire[12:0] T1276;
  wire[12:0] T1277;
  wire[12:0] T1278;
  wire T1279;
  wire[12:0] T1280;
  wire[12:0] T1281;
  wire[12:0] T1282;
  wire T1283;
  wire[12:0] T1284;
  wire[12:0] T1285;
  wire[12:0] T1286;
  wire T1287;
  wire[12:0] T1288;
  wire[12:0] T1289;
  wire[12:0] T1290;
  wire T1291;
  wire[12:0] T1292;
  wire[12:0] T1293;
  wire[12:0] T1294;
  wire T1295;
  wire[12:0] T1296;
  wire[12:0] T1297;
  wire[12:0] T1298;
  wire T1299;
  wire[12:0] T1300;
  wire[12:0] T1301;
  wire[12:0] T1302;
  wire T1303;
  wire[12:0] T1304;
  wire[12:0] T1305;
  wire[12:0] T1306;
  wire T1307;
  wire[12:0] T1308;
  wire[12:0] T1309;
  wire[12:0] T1310;
  wire T1311;
  wire[12:0] T1312;
  wire[12:0] T1313;
  wire[12:0] T1314;
  wire T1315;
  wire[12:0] T1316;
  wire[12:0] T1317;
  wire[12:0] T1318;
  wire T1319;
  wire[12:0] T1320;
  wire[12:0] T1321;
  wire T1322;
  wire[29:0] T1323;
  wire[29:0] T1324;
  wire[29:0] T1325;
  wire T1326;
  wire[5:0] T1327;
  wire[5:0] T1328;
  wire T1329;
  wire[5:0] T1330;
  wire[5:0] T1331;
  wire T1332;
  wire[5:0] T1333;
  wire[5:0] T1334;
  wire T1335;
  wire[5:0] T1336;
  wire[5:0] T1337;
  wire T1338;
  wire[5:0] T1339;
  wire[5:0] T1340;
  wire T1341;
  wire[5:0] T1342;
  wire[5:0] T1343;
  wire T1344;
  wire[5:0] T1345;
  wire[5:0] T1346;
  wire T1347;
  wire[5:0] T1348;
  wire[5:0] T1349;
  wire T1350;
  wire[5:0] T1351;
  wire[5:0] T1352;
  wire T1353;
  wire[5:0] T1354;
  wire[5:0] T1355;
  wire T1356;
  wire[5:0] T1357;
  wire[5:0] T1358;
  wire T1359;
  wire[5:0] T1360;
  wire[5:0] T1361;
  wire T1362;
  wire[5:0] T1363;
  wire[5:0] T1364;
  wire T1365;
  wire[5:0] T1366;
  wire[5:0] T1367;
  wire T1368;
  wire[5:0] T1369;
  wire[5:0] T1370;
  wire T1371;
  wire[5:0] T1372;
  wire[5:0] T1373;
  wire T1374;
  wire[5:0] T1375;
  wire[5:0] T1376;
  wire T1377;
  wire[5:0] T1378;
  wire[5:0] T1379;
  wire T1380;
  wire[5:0] T1381;
  wire[5:0] T1382;
  wire T1383;
  wire[5:0] T1384;
  wire[5:0] T1385;
  wire T1386;
  wire[5:0] T1387;
  wire[5:0] T1388;
  wire T1389;
  wire[5:0] T1390;
  wire[5:0] T1391;
  wire T1392;
  wire[5:0] T1393;
  wire[5:0] T1394;
  wire T1395;
  wire[5:0] T1396;
  wire[5:0] T1397;
  wire T1398;
  wire[5:0] T1399;
  wire[5:0] T1400;
  wire T1401;
  wire[5:0] T1402;
  wire[5:0] T1403;
  wire T1404;
  wire[5:0] T1405;
  wire[5:0] T1406;
  wire T1407;
  wire[5:0] T1408;
  wire[5:0] T1409;
  wire T1410;
  wire[5:0] T1411;
  wire[5:0] T1412;
  wire T1413;
  wire[5:0] T1414;
  wire[5:0] T1415;
  wire T1416;
  wire[5:0] T1417;
  wire[5:0] T1418;
  wire T1419;
  wire[5:0] T1420;
  wire[5:0] T1421;
  wire T1422;
  wire[5:0] T1423;
  wire[5:0] T1424;
  wire T1425;
  wire[5:0] T1426;
  wire[5:0] T1427;
  wire T1428;
  wire[5:0] T1429;
  wire[5:0] T1430;
  wire T1431;
  wire[5:0] T1432;
  wire[5:0] T1433;
  wire T1434;
  wire[5:0] T1435;
  wire[5:0] T1436;
  wire T1437;
  wire[5:0] T1438;
  wire[5:0] T1439;
  wire T1440;
  wire[5:0] T1441;
  wire[5:0] T1442;
  wire T1443;
  wire[5:0] T1444;
  wire[5:0] T1445;
  wire T1446;
  wire[5:0] T1447;
  wire[5:0] T1448;
  wire T1449;
  wire[5:0] T1450;
  wire[5:0] T1451;
  wire T1452;
  wire[5:0] T1453;
  wire[5:0] T1454;
  wire T1455;
  wire[5:0] T1456;
  wire[5:0] T1457;
  wire T1458;
  wire[5:0] T1459;
  wire[5:0] T1460;
  wire T1461;
  wire[5:0] T1462;
  wire[5:0] T1463;
  wire T1464;
  wire[5:0] T1465;
  wire[5:0] T1466;
  wire T1467;
  wire[5:0] T1468;
  wire[5:0] T1469;
  wire T1470;
  wire[5:0] T1471;
  wire[5:0] T1472;
  wire T1473;
  wire[5:0] T1474;
  wire[5:0] T1475;
  wire T1476;
  wire[5:0] T1477;
  wire[5:0] T1478;
  wire T1479;
  wire[5:0] T1480;
  wire[5:0] T1481;
  wire T1482;
  wire[5:0] T1483;
  wire[5:0] T1484;
  wire T1485;
  wire[5:0] T1486;
  wire[5:0] T1487;
  wire T1488;
  wire[5:0] T1489;
  wire[5:0] T1490;
  wire T1491;
  wire[5:0] T1492;
  wire[5:0] T1493;
  wire T1494;
  wire[5:0] T1495;
  wire[5:0] T1496;
  wire T1497;
  wire[5:0] T1498;
  wire[5:0] T1499;
  wire T1500;
  wire[5:0] T1501;
  wire[5:0] T1502;
  wire T1503;
  wire[5:0] T1504;
  wire[5:0] T1505;
  wire T1506;
  wire[5:0] T1507;
  wire[5:0] T1508;
  wire T1509;
  wire[5:0] T1510;
  wire T1511;
  wire[29:0] T1512;
  wire[29:0] T1513;
  wire[29:0] T1514;
  wire T1515;
  wire[29:0] T1516;
  wire[29:0] T1517;
  wire[29:0] T1518;
  wire T1519;
  wire[29:0] T1520;
  wire[29:0] T1521;
  wire[29:0] T1522;
  wire T1523;
  wire[29:0] T1524;
  wire[29:0] T1525;
  wire[29:0] T1526;
  wire T1527;
  wire[29:0] T1528;
  wire[29:0] T1529;
  wire T1530;
  wire[42:0] T1531;
  reg [42:0] R1532;
  wire[42:0] T1533;
  wire T1534;
  wire T1535;
  wire[1:0] T1536;
  wire T1537;
  wire T1538;
  reg  R1539;
  wire T1725;
  wire T1540;
  wire T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire T1545;
  reg [1:0] R1546;
  wire[1:0] T1726;
  wire[1:0] T1547;
  wire[1:0] T1548;
  wire[1:0] T1549;
  wire[1:0] T1550;
  wire T1551;
  wire T1552;
  wire[1:0] T1553;
  wire T1554;
  wire T1555;
  wire T1556;
  wire T1557;
  wire T1558;
  reg [42:0] R1559;
  wire[42:0] T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire T1564;
  wire T1565;
  wire[61:0] T1566;
  reg [61:0] useRAS;
  wire[61:0] T1727;
  wire[63:0] T1567;
  wire[63:0] T1728;
  wire[63:0] T1568;
  wire[63:0] T1569;
  wire[63:0] T1570;
  wire[63:0] T1729;
  wire[61:0] T1571;
  wire[63:0] T1572;
  wire[63:0] T1730;
  wire T1573;
  wire T1574;
  reg  R1575;
  wire T1576;
  wire[63:0] T1577;
  wire[63:0] T1578;
  wire[63:0] T1731;
  wire T1579;
  wire T1580;
  wire T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire T1585;
  wire[61:0] T1586;
  wire T1587;
  wire T1588;
  wire T1589;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R8 = {1{$random}};
    R11 = {1{$random}};
    updateHit = {1{$random}};
    R18 = {1{$random}};
    for (initvar = 0; initvar < 128; initvar = initvar+1)
      T21[initvar] = {1{$random}};
    R38 = {1{$random}};
    isJump = {2{$random}};
    R55 = {1{$random}};
    R63 = {1{$random}};
    R67 = {1{$random}};
    pageValid = {1{$random}};
    R88 = {1{$random}};
    R101 = {2{$random}};
    for (initvar = 0; initvar < 6; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {2{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R1532 = {2{$random}};
    R1539 = {1{$random}};
    R1546 = {1{$random}};
    R1559 = {2{$random}};
    useRAS = {2{$random}};
    R1575 = {1{$random}};
  end
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_update_valid ? io_update_bits_target : R4;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T14 & updateTarget;
  assign updateTarget = T10 & R8;
  assign T9 = io_update_valid ? io_update_bits_taken : R8;
  assign T10 = updateValid & R11;
  assign T12 = io_update_valid ? io_update_bits_mispredict : R11;
  assign updateValid = R11 | updateHit;
  assign T13 = io_update_valid ? io_update_bits_prediction_valid : updateHit;
  assign T14 = R18 & T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = updateValid & T17;
  assign T17 = updateTarget ^ 1'h1;
  assign T1590 = reset ? 1'h0 : io_update_valid;
  assign io_resp_bits_bht_value = T19;
  assign T19 = T20;
  assign T20 = T21[T37];
  assign T23 = {io_update_bits_taken, T24};
  assign T24 = T29 | T25;
  assign T25 = T26 & io_update_bits_taken;
  assign T26 = T28 | T27;
  assign T27 = io_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T28 = io_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T29 = T31 & T30;
  assign T30 = io_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T31 = io_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T32 = T34 & T33;
  assign T33 = io_update_bits_isJump ^ 1'h1;
  assign T34 = io_update_valid & io_update_bits_prediction_valid;
  assign T35 = T36 ^ io_update_bits_prediction_bits_bht_history;
  assign T36 = io_update_bits_pc[4'h8:2'h2];
  assign T37 = T1067 ^ R38;
  assign T39 = T1066 ? T1064 : T40;
  assign T40 = T44 ? T41 : R38;
  assign T41 = {T43, T42};
  assign T42 = R38[3'h6:1'h1];
  assign T43 = T19[1'h0:1'h0];
  assign T44 = T1062 & T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 != 62'h0;
  assign T47 = hits & isJump;
  assign T1591 = T48[6'h3d:1'h0];
  assign T48 = T7 ? T49 : T1592;
  assign T1592 = {2'h0, isJump};
  assign T49 = T69 | T50;
  assign T50 = T1595 & T51;
  assign T51 = T53 | T1593;
  assign T1593 = {2'h0, T52};
  assign T52 = isJump ^ isJump;
  assign T53 = 1'h1 << T54;
  assign T54 = updateHit ? R63 : R55;
  assign T1594 = reset ? 6'h0 : T56;
  assign T56 = T60 ? T57 : R55;
  assign T57 = T59 ? 6'h0 : T58;
  assign T58 = R55 + 6'h1;
  assign T59 = R55 == 6'h3d;
  assign T60 = T14 & T61;
  assign T61 = T62 & updateValid;
  assign T62 = updateHit ^ 1'h1;
  assign T64 = io_update_valid ? io_update_bits_prediction_bits_entry : R63;
  assign T1595 = T65 ? 64'hffffffffffffffff : 64'h0;
  assign T65 = T66;
  assign T66 = R67;
  assign T68 = io_update_valid ? io_update_bits_isJump : R67;
  assign T69 = T1596 & T70;
  assign T70 = ~ T51;
  assign T1596 = {2'h0, isJump};
  assign hits = T481 & T71;
  assign T71 = T72;
  assign T72 = {T327, T73};
  assign T73 = {T253, T74};
  assign T74 = {T214, T75};
  assign T75 = {T195, T76};
  assign T76 = {T186, T77};
  assign T77 = {T182, T78};
  assign T78 = T79 != 6'h0;
  assign T79 = idxPagesOH_0 & pageHit;
  assign pageHit = T158 & pageValid;
  assign T1597 = T1598[3'h5:1'h0];
  assign T1598 = reset ? 8'h0 : T80;
  assign T80 = io_invalidate ? 8'h0 : T81;
  assign T81 = T157 ? T82 : T1599;
  assign T1599 = {2'h0, pageValid};
  assign T82 = T1605 | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T1600;
  assign T1600 = {2'h0, T83};
  assign T83 = T85 | T1601;
  assign T1601 = {5'h0, T84};
  assign T84 = idxPageUpdateOH[3'h5:3'h5];
  assign T85 = T86 << 1'h1;
  assign T86 = idxPageUpdateOH[3'h4:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? T1603 : idxPageRepl;
  assign idxPageRepl = T87;
  assign T87 = 1'h1 << R88;
  assign T1602 = reset ? 3'h0 : T89;
  assign T89 = T93 ? T90 : R88;
  assign T90 = T92 ? 3'h0 : T91;
  assign T91 = R88 + 3'h1;
  assign T92 = R88 == 3'h5;
  assign T93 = R18 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = updateTarget & T94;
  assign T94 = useUpdatePageHit ^ 1'h1;
  assign T1603 = {2'h0, updatePageHit};
  assign updatePageHit = T95 & pageValid;
  assign T95 = T96;
  assign T96 = {T142, T97};
  assign T97 = {T140, T98};
  assign T98 = {T138, T99};
  assign T99 = T103 == T100;
  assign T100 = R101 >> 4'hd;
  assign T102 = io_update_valid ? io_update_bits_pc : R101;
  assign T103 = pages[3'h0];
  assign T105 = T108 ? T107 : T106;
  assign T106 = R101 >> 4'hd;
  assign T107 = io_req_bits_addr >> 4'hd;
  assign T108 = T109 != 8'h0;
  assign T109 = idxPageUpdateOH & 8'h15;
  assign T110 = T14 & T111;
  assign T111 = T113 & T112;
  assign T112 = pageReplEn[3'h5:3'h5];
  assign T113 = T108 ? doTgtPageRepl : doIdxPageRepl;
  assign T115 = T14 & T116;
  assign T116 = T113 & T117;
  assign T117 = pageReplEn[2'h3:2'h3];
  assign T119 = T14 & T120;
  assign T120 = T113 & T121;
  assign T121 = pageReplEn[1'h1:1'h1];
  assign T123 = T108 ? T125 : T124;
  assign T124 = io_req_bits_addr >> 4'hd;
  assign T125 = R101 >> 4'hd;
  assign T126 = T14 & T127;
  assign T127 = T129 & T128;
  assign T128 = pageReplEn[3'h4:3'h4];
  assign T129 = T108 ? doIdxPageRepl : doTgtPageRepl;
  assign T131 = T14 & T132;
  assign T132 = T129 & T133;
  assign T133 = pageReplEn[2'h2:2'h2];
  assign T135 = T14 & T136;
  assign T136 = T129 & T137;
  assign T137 = pageReplEn[1'h0:1'h0];
  assign T138 = T139 == T100;
  assign T139 = pages[3'h1];
  assign T140 = T141 == T100;
  assign T141 = pages[3'h2];
  assign T142 = {T148, T143};
  assign T143 = {T146, T144};
  assign T144 = T145 == T100;
  assign T145 = pages[3'h3];
  assign T146 = T147 == T100;
  assign T147 = pages[3'h4];
  assign T148 = T149 == T100;
  assign T149 = pages[3'h5];
  assign useUpdatePageHit = updatePageHit != 6'h0;
  assign samePage = T151 == T150;
  assign T150 = io_req_bits_addr >> 4'hd;
  assign T151 = R101 >> 4'hd;
  assign doTgtPageRepl = T155 & T152;
  assign T152 = usePageHit ^ 1'h1;
  assign usePageHit = T153 != 8'h0;
  assign T153 = T1604 & T154;
  assign T154 = ~ idxPageReplEn;
  assign T1604 = {2'h0, pageHit};
  assign T155 = updateTarget & T156;
  assign T156 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0;
  assign T1605 = {2'h0, pageValid};
  assign T157 = T14 & doPageRepl;
  assign T158 = T159;
  assign T159 = {T169, T160};
  assign T160 = {T167, T161};
  assign T161 = {T165, T162};
  assign T162 = T164 == T163;
  assign T163 = io_req_bits_addr >> 4'hd;
  assign T164 = pages[3'h0];
  assign T165 = T166 == T163;
  assign T166 = pages[3'h1];
  assign T167 = T168 == T163;
  assign T168 = pages[3'h2];
  assign T169 = {T175, T170};
  assign T170 = {T173, T171};
  assign T171 = T172 == T163;
  assign T172 = pages[3'h3];
  assign T173 = T174 == T163;
  assign T174 = pages[3'h4];
  assign T175 = T176 == T163;
  assign T176 = pages[3'h5];
  assign idxPagesOH_0 = T177[3'h5:1'h0];
  assign T177 = 1'h1 << T178;
  assign T178 = idxPages[6'h0];
  assign T1606 = {T1616, T1607};
  assign T1607 = {T1615, T1608};
  assign T1608 = T1609[1'h1:1'h1];
  assign T1609 = T1614 | T1610;
  assign T1610 = T1611[1'h1:1'h0];
  assign T1611 = T1613 | T1612;
  assign T1612 = idxPageUpdateOH[2'h3:1'h0];
  assign T1613 = idxPageUpdateOH[3'h7:3'h4];
  assign T1614 = T1611[2'h3:2'h2];
  assign T1615 = T1614 != 2'h0;
  assign T1616 = T1613 != 4'h0;
  assign T180 = T7 & T181;
  assign T181 = T54 < 6'h3e;
  assign T182 = T183 != 6'h0;
  assign T183 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T184[3'h5:1'h0];
  assign T184 = 1'h1 << T185;
  assign T185 = idxPages[6'h1];
  assign T186 = {T191, T187};
  assign T187 = T188 != 6'h0;
  assign T188 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T189[3'h5:1'h0];
  assign T189 = 1'h1 << T190;
  assign T190 = idxPages[6'h2];
  assign T191 = T192 != 6'h0;
  assign T192 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T193[3'h5:1'h0];
  assign T193 = 1'h1 << T194;
  assign T194 = idxPages[6'h3];
  assign T195 = {T205, T196};
  assign T196 = {T201, T197};
  assign T197 = T198 != 6'h0;
  assign T198 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T199[3'h5:1'h0];
  assign T199 = 1'h1 << T200;
  assign T200 = idxPages[6'h4];
  assign T201 = T202 != 6'h0;
  assign T202 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T203[3'h5:1'h0];
  assign T203 = 1'h1 << T204;
  assign T204 = idxPages[6'h5];
  assign T205 = {T210, T206};
  assign T206 = T207 != 6'h0;
  assign T207 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T208[3'h5:1'h0];
  assign T208 = 1'h1 << T209;
  assign T209 = idxPages[6'h6];
  assign T210 = T211 != 6'h0;
  assign T211 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T212[3'h5:1'h0];
  assign T212 = 1'h1 << T213;
  assign T213 = idxPages[6'h7];
  assign T214 = {T234, T215};
  assign T215 = {T225, T216};
  assign T216 = {T221, T217};
  assign T217 = T218 != 6'h0;
  assign T218 = idxPagesOH_8 & pageHit;
  assign idxPagesOH_8 = T219[3'h5:1'h0];
  assign T219 = 1'h1 << T220;
  assign T220 = idxPages[6'h8];
  assign T221 = T222 != 6'h0;
  assign T222 = idxPagesOH_9 & pageHit;
  assign idxPagesOH_9 = T223[3'h5:1'h0];
  assign T223 = 1'h1 << T224;
  assign T224 = idxPages[6'h9];
  assign T225 = {T230, T226};
  assign T226 = T227 != 6'h0;
  assign T227 = idxPagesOH_10 & pageHit;
  assign idxPagesOH_10 = T228[3'h5:1'h0];
  assign T228 = 1'h1 << T229;
  assign T229 = idxPages[6'ha];
  assign T230 = T231 != 6'h0;
  assign T231 = idxPagesOH_11 & pageHit;
  assign idxPagesOH_11 = T232[3'h5:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = idxPages[6'hb];
  assign T234 = {T244, T235};
  assign T235 = {T240, T236};
  assign T236 = T237 != 6'h0;
  assign T237 = idxPagesOH_12 & pageHit;
  assign idxPagesOH_12 = T238[3'h5:1'h0];
  assign T238 = 1'h1 << T239;
  assign T239 = idxPages[6'hc];
  assign T240 = T241 != 6'h0;
  assign T241 = idxPagesOH_13 & pageHit;
  assign idxPagesOH_13 = T242[3'h5:1'h0];
  assign T242 = 1'h1 << T243;
  assign T243 = idxPages[6'hd];
  assign T244 = {T249, T245};
  assign T245 = T246 != 6'h0;
  assign T246 = idxPagesOH_14 & pageHit;
  assign idxPagesOH_14 = T247[3'h5:1'h0];
  assign T247 = 1'h1 << T248;
  assign T248 = idxPages[6'he];
  assign T249 = T250 != 6'h0;
  assign T250 = idxPagesOH_15 & pageHit;
  assign idxPagesOH_15 = T251[3'h5:1'h0];
  assign T251 = 1'h1 << T252;
  assign T252 = idxPages[6'hf];
  assign T253 = {T293, T254};
  assign T254 = {T274, T255};
  assign T255 = {T265, T256};
  assign T256 = {T261, T257};
  assign T257 = T258 != 6'h0;
  assign T258 = idxPagesOH_16 & pageHit;
  assign idxPagesOH_16 = T259[3'h5:1'h0];
  assign T259 = 1'h1 << T260;
  assign T260 = idxPages[6'h10];
  assign T261 = T262 != 6'h0;
  assign T262 = idxPagesOH_17 & pageHit;
  assign idxPagesOH_17 = T263[3'h5:1'h0];
  assign T263 = 1'h1 << T264;
  assign T264 = idxPages[6'h11];
  assign T265 = {T270, T266};
  assign T266 = T267 != 6'h0;
  assign T267 = idxPagesOH_18 & pageHit;
  assign idxPagesOH_18 = T268[3'h5:1'h0];
  assign T268 = 1'h1 << T269;
  assign T269 = idxPages[6'h12];
  assign T270 = T271 != 6'h0;
  assign T271 = idxPagesOH_19 & pageHit;
  assign idxPagesOH_19 = T272[3'h5:1'h0];
  assign T272 = 1'h1 << T273;
  assign T273 = idxPages[6'h13];
  assign T274 = {T284, T275};
  assign T275 = {T280, T276};
  assign T276 = T277 != 6'h0;
  assign T277 = idxPagesOH_20 & pageHit;
  assign idxPagesOH_20 = T278[3'h5:1'h0];
  assign T278 = 1'h1 << T279;
  assign T279 = idxPages[6'h14];
  assign T280 = T281 != 6'h0;
  assign T281 = idxPagesOH_21 & pageHit;
  assign idxPagesOH_21 = T282[3'h5:1'h0];
  assign T282 = 1'h1 << T283;
  assign T283 = idxPages[6'h15];
  assign T284 = {T289, T285};
  assign T285 = T286 != 6'h0;
  assign T286 = idxPagesOH_22 & pageHit;
  assign idxPagesOH_22 = T287[3'h5:1'h0];
  assign T287 = 1'h1 << T288;
  assign T288 = idxPages[6'h16];
  assign T289 = T290 != 6'h0;
  assign T290 = idxPagesOH_23 & pageHit;
  assign idxPagesOH_23 = T291[3'h5:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = idxPages[6'h17];
  assign T293 = {T313, T294};
  assign T294 = {T304, T295};
  assign T295 = {T300, T296};
  assign T296 = T297 != 6'h0;
  assign T297 = idxPagesOH_24 & pageHit;
  assign idxPagesOH_24 = T298[3'h5:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = idxPages[6'h18];
  assign T300 = T301 != 6'h0;
  assign T301 = idxPagesOH_25 & pageHit;
  assign idxPagesOH_25 = T302[3'h5:1'h0];
  assign T302 = 1'h1 << T303;
  assign T303 = idxPages[6'h19];
  assign T304 = {T309, T305};
  assign T305 = T306 != 6'h0;
  assign T306 = idxPagesOH_26 & pageHit;
  assign idxPagesOH_26 = T307[3'h5:1'h0];
  assign T307 = 1'h1 << T308;
  assign T308 = idxPages[6'h1a];
  assign T309 = T310 != 6'h0;
  assign T310 = idxPagesOH_27 & pageHit;
  assign idxPagesOH_27 = T311[3'h5:1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = idxPages[6'h1b];
  assign T313 = {T323, T314};
  assign T314 = {T319, T315};
  assign T315 = T316 != 6'h0;
  assign T316 = idxPagesOH_28 & pageHit;
  assign idxPagesOH_28 = T317[3'h5:1'h0];
  assign T317 = 1'h1 << T318;
  assign T318 = idxPages[6'h1c];
  assign T319 = T320 != 6'h0;
  assign T320 = idxPagesOH_29 & pageHit;
  assign idxPagesOH_29 = T321[3'h5:1'h0];
  assign T321 = 1'h1 << T322;
  assign T322 = idxPages[6'h1d];
  assign T323 = T324 != 6'h0;
  assign T324 = idxPagesOH_30 & pageHit;
  assign idxPagesOH_30 = T325[3'h5:1'h0];
  assign T325 = 1'h1 << T326;
  assign T326 = idxPages[6'h1e];
  assign T327 = {T407, T328};
  assign T328 = {T368, T329};
  assign T329 = {T349, T330};
  assign T330 = {T340, T331};
  assign T331 = {T336, T332};
  assign T332 = T333 != 6'h0;
  assign T333 = idxPagesOH_31 & pageHit;
  assign idxPagesOH_31 = T334[3'h5:1'h0];
  assign T334 = 1'h1 << T335;
  assign T335 = idxPages[6'h1f];
  assign T336 = T337 != 6'h0;
  assign T337 = idxPagesOH_32 & pageHit;
  assign idxPagesOH_32 = T338[3'h5:1'h0];
  assign T338 = 1'h1 << T339;
  assign T339 = idxPages[6'h20];
  assign T340 = {T345, T341};
  assign T341 = T342 != 6'h0;
  assign T342 = idxPagesOH_33 & pageHit;
  assign idxPagesOH_33 = T343[3'h5:1'h0];
  assign T343 = 1'h1 << T344;
  assign T344 = idxPages[6'h21];
  assign T345 = T346 != 6'h0;
  assign T346 = idxPagesOH_34 & pageHit;
  assign idxPagesOH_34 = T347[3'h5:1'h0];
  assign T347 = 1'h1 << T348;
  assign T348 = idxPages[6'h22];
  assign T349 = {T359, T350};
  assign T350 = {T355, T351};
  assign T351 = T352 != 6'h0;
  assign T352 = idxPagesOH_35 & pageHit;
  assign idxPagesOH_35 = T353[3'h5:1'h0];
  assign T353 = 1'h1 << T354;
  assign T354 = idxPages[6'h23];
  assign T355 = T356 != 6'h0;
  assign T356 = idxPagesOH_36 & pageHit;
  assign idxPagesOH_36 = T357[3'h5:1'h0];
  assign T357 = 1'h1 << T358;
  assign T358 = idxPages[6'h24];
  assign T359 = {T364, T360};
  assign T360 = T361 != 6'h0;
  assign T361 = idxPagesOH_37 & pageHit;
  assign idxPagesOH_37 = T362[3'h5:1'h0];
  assign T362 = 1'h1 << T363;
  assign T363 = idxPages[6'h25];
  assign T364 = T365 != 6'h0;
  assign T365 = idxPagesOH_38 & pageHit;
  assign idxPagesOH_38 = T366[3'h5:1'h0];
  assign T366 = 1'h1 << T367;
  assign T367 = idxPages[6'h26];
  assign T368 = {T388, T369};
  assign T369 = {T379, T370};
  assign T370 = {T375, T371};
  assign T371 = T372 != 6'h0;
  assign T372 = idxPagesOH_39 & pageHit;
  assign idxPagesOH_39 = T373[3'h5:1'h0];
  assign T373 = 1'h1 << T374;
  assign T374 = idxPages[6'h27];
  assign T375 = T376 != 6'h0;
  assign T376 = idxPagesOH_40 & pageHit;
  assign idxPagesOH_40 = T377[3'h5:1'h0];
  assign T377 = 1'h1 << T378;
  assign T378 = idxPages[6'h28];
  assign T379 = {T384, T380};
  assign T380 = T381 != 6'h0;
  assign T381 = idxPagesOH_41 & pageHit;
  assign idxPagesOH_41 = T382[3'h5:1'h0];
  assign T382 = 1'h1 << T383;
  assign T383 = idxPages[6'h29];
  assign T384 = T385 != 6'h0;
  assign T385 = idxPagesOH_42 & pageHit;
  assign idxPagesOH_42 = T386[3'h5:1'h0];
  assign T386 = 1'h1 << T387;
  assign T387 = idxPages[6'h2a];
  assign T388 = {T398, T389};
  assign T389 = {T394, T390};
  assign T390 = T391 != 6'h0;
  assign T391 = idxPagesOH_43 & pageHit;
  assign idxPagesOH_43 = T392[3'h5:1'h0];
  assign T392 = 1'h1 << T393;
  assign T393 = idxPages[6'h2b];
  assign T394 = T395 != 6'h0;
  assign T395 = idxPagesOH_44 & pageHit;
  assign idxPagesOH_44 = T396[3'h5:1'h0];
  assign T396 = 1'h1 << T397;
  assign T397 = idxPages[6'h2c];
  assign T398 = {T403, T399};
  assign T399 = T400 != 6'h0;
  assign T400 = idxPagesOH_45 & pageHit;
  assign idxPagesOH_45 = T401[3'h5:1'h0];
  assign T401 = 1'h1 << T402;
  assign T402 = idxPages[6'h2d];
  assign T403 = T404 != 6'h0;
  assign T404 = idxPagesOH_46 & pageHit;
  assign idxPagesOH_46 = T405[3'h5:1'h0];
  assign T405 = 1'h1 << T406;
  assign T406 = idxPages[6'h2e];
  assign T407 = {T447, T408};
  assign T408 = {T428, T409};
  assign T409 = {T419, T410};
  assign T410 = {T415, T411};
  assign T411 = T412 != 6'h0;
  assign T412 = idxPagesOH_47 & pageHit;
  assign idxPagesOH_47 = T413[3'h5:1'h0];
  assign T413 = 1'h1 << T414;
  assign T414 = idxPages[6'h2f];
  assign T415 = T416 != 6'h0;
  assign T416 = idxPagesOH_48 & pageHit;
  assign idxPagesOH_48 = T417[3'h5:1'h0];
  assign T417 = 1'h1 << T418;
  assign T418 = idxPages[6'h30];
  assign T419 = {T424, T420};
  assign T420 = T421 != 6'h0;
  assign T421 = idxPagesOH_49 & pageHit;
  assign idxPagesOH_49 = T422[3'h5:1'h0];
  assign T422 = 1'h1 << T423;
  assign T423 = idxPages[6'h31];
  assign T424 = T425 != 6'h0;
  assign T425 = idxPagesOH_50 & pageHit;
  assign idxPagesOH_50 = T426[3'h5:1'h0];
  assign T426 = 1'h1 << T427;
  assign T427 = idxPages[6'h32];
  assign T428 = {T438, T429};
  assign T429 = {T434, T430};
  assign T430 = T431 != 6'h0;
  assign T431 = idxPagesOH_51 & pageHit;
  assign idxPagesOH_51 = T432[3'h5:1'h0];
  assign T432 = 1'h1 << T433;
  assign T433 = idxPages[6'h33];
  assign T434 = T435 != 6'h0;
  assign T435 = idxPagesOH_52 & pageHit;
  assign idxPagesOH_52 = T436[3'h5:1'h0];
  assign T436 = 1'h1 << T437;
  assign T437 = idxPages[6'h34];
  assign T438 = {T443, T439};
  assign T439 = T440 != 6'h0;
  assign T440 = idxPagesOH_53 & pageHit;
  assign idxPagesOH_53 = T441[3'h5:1'h0];
  assign T441 = 1'h1 << T442;
  assign T442 = idxPages[6'h35];
  assign T443 = T444 != 6'h0;
  assign T444 = idxPagesOH_54 & pageHit;
  assign idxPagesOH_54 = T445[3'h5:1'h0];
  assign T445 = 1'h1 << T446;
  assign T446 = idxPages[6'h36];
  assign T447 = {T467, T448};
  assign T448 = {T458, T449};
  assign T449 = {T454, T450};
  assign T450 = T451 != 6'h0;
  assign T451 = idxPagesOH_55 & pageHit;
  assign idxPagesOH_55 = T452[3'h5:1'h0];
  assign T452 = 1'h1 << T453;
  assign T453 = idxPages[6'h37];
  assign T454 = T455 != 6'h0;
  assign T455 = idxPagesOH_56 & pageHit;
  assign idxPagesOH_56 = T456[3'h5:1'h0];
  assign T456 = 1'h1 << T457;
  assign T457 = idxPages[6'h38];
  assign T458 = {T463, T459};
  assign T459 = T460 != 6'h0;
  assign T460 = idxPagesOH_57 & pageHit;
  assign idxPagesOH_57 = T461[3'h5:1'h0];
  assign T461 = 1'h1 << T462;
  assign T462 = idxPages[6'h39];
  assign T463 = T464 != 6'h0;
  assign T464 = idxPagesOH_58 & pageHit;
  assign idxPagesOH_58 = T465[3'h5:1'h0];
  assign T465 = 1'h1 << T466;
  assign T466 = idxPages[6'h3a];
  assign T467 = {T477, T468};
  assign T468 = {T473, T469};
  assign T469 = T470 != 6'h0;
  assign T470 = idxPagesOH_59 & pageHit;
  assign idxPagesOH_59 = T471[3'h5:1'h0];
  assign T471 = 1'h1 << T472;
  assign T472 = idxPages[6'h3b];
  assign T473 = T474 != 6'h0;
  assign T474 = idxPagesOH_60 & pageHit;
  assign idxPagesOH_60 = T475[3'h5:1'h0];
  assign T475 = 1'h1 << T476;
  assign T476 = idxPages[6'h3c];
  assign T477 = T478 != 6'h0;
  assign T478 = idxPagesOH_61 & pageHit;
  assign idxPagesOH_61 = T479[3'h5:1'h0];
  assign T479 = 1'h1 << T480;
  assign T480 = idxPages[6'h3d];
  assign T481 = idxValid & T482;
  assign T482 = T483;
  assign T483 = {T580, T484};
  assign T484 = {T536, T485};
  assign T485 = {T513, T486};
  assign T486 = {T502, T487};
  assign T487 = {T497, T488};
  assign T488 = {T495, T489};
  assign T489 = T491 == T490;
  assign T490 = io_req_bits_addr[4'hc:1'h0];
  assign T491 = idxs[6'h0];
  assign T1617 = R101[4'hc:1'h0];
  assign T493 = T7 & T494;
  assign T494 = T54 < 6'h3e;
  assign T495 = T496 == T490;
  assign T496 = idxs[6'h1];
  assign T497 = {T500, T498};
  assign T498 = T499 == T490;
  assign T499 = idxs[6'h2];
  assign T500 = T501 == T490;
  assign T501 = idxs[6'h3];
  assign T502 = {T508, T503};
  assign T503 = {T506, T504};
  assign T504 = T505 == T490;
  assign T505 = idxs[6'h4];
  assign T506 = T507 == T490;
  assign T507 = idxs[6'h5];
  assign T508 = {T511, T509};
  assign T509 = T510 == T490;
  assign T510 = idxs[6'h6];
  assign T511 = T512 == T490;
  assign T512 = idxs[6'h7];
  assign T513 = {T525, T514};
  assign T514 = {T520, T515};
  assign T515 = {T518, T516};
  assign T516 = T517 == T490;
  assign T517 = idxs[6'h8];
  assign T518 = T519 == T490;
  assign T519 = idxs[6'h9];
  assign T520 = {T523, T521};
  assign T521 = T522 == T490;
  assign T522 = idxs[6'ha];
  assign T523 = T524 == T490;
  assign T524 = idxs[6'hb];
  assign T525 = {T531, T526};
  assign T526 = {T529, T527};
  assign T527 = T528 == T490;
  assign T528 = idxs[6'hc];
  assign T529 = T530 == T490;
  assign T530 = idxs[6'hd];
  assign T531 = {T534, T532};
  assign T532 = T533 == T490;
  assign T533 = idxs[6'he];
  assign T534 = T535 == T490;
  assign T535 = idxs[6'hf];
  assign T536 = {T560, T537};
  assign T537 = {T549, T538};
  assign T538 = {T544, T539};
  assign T539 = {T542, T540};
  assign T540 = T541 == T490;
  assign T541 = idxs[6'h10];
  assign T542 = T543 == T490;
  assign T543 = idxs[6'h11];
  assign T544 = {T547, T545};
  assign T545 = T546 == T490;
  assign T546 = idxs[6'h12];
  assign T547 = T548 == T490;
  assign T548 = idxs[6'h13];
  assign T549 = {T555, T550};
  assign T550 = {T553, T551};
  assign T551 = T552 == T490;
  assign T552 = idxs[6'h14];
  assign T553 = T554 == T490;
  assign T554 = idxs[6'h15];
  assign T555 = {T558, T556};
  assign T556 = T557 == T490;
  assign T557 = idxs[6'h16];
  assign T558 = T559 == T490;
  assign T559 = idxs[6'h17];
  assign T560 = {T572, T561};
  assign T561 = {T567, T562};
  assign T562 = {T565, T563};
  assign T563 = T564 == T490;
  assign T564 = idxs[6'h18];
  assign T565 = T566 == T490;
  assign T566 = idxs[6'h19];
  assign T567 = {T570, T568};
  assign T568 = T569 == T490;
  assign T569 = idxs[6'h1a];
  assign T570 = T571 == T490;
  assign T571 = idxs[6'h1b];
  assign T572 = {T578, T573};
  assign T573 = {T576, T574};
  assign T574 = T575 == T490;
  assign T575 = idxs[6'h1c];
  assign T576 = T577 == T490;
  assign T577 = idxs[6'h1d];
  assign T578 = T579 == T490;
  assign T579 = idxs[6'h1e];
  assign T580 = {T628, T581};
  assign T581 = {T605, T582};
  assign T582 = {T594, T583};
  assign T583 = {T589, T584};
  assign T584 = {T587, T585};
  assign T585 = T586 == T490;
  assign T586 = idxs[6'h1f];
  assign T587 = T588 == T490;
  assign T588 = idxs[6'h20];
  assign T589 = {T592, T590};
  assign T590 = T591 == T490;
  assign T591 = idxs[6'h21];
  assign T592 = T593 == T490;
  assign T593 = idxs[6'h22];
  assign T594 = {T600, T595};
  assign T595 = {T598, T596};
  assign T596 = T597 == T490;
  assign T597 = idxs[6'h23];
  assign T598 = T599 == T490;
  assign T599 = idxs[6'h24];
  assign T600 = {T603, T601};
  assign T601 = T602 == T490;
  assign T602 = idxs[6'h25];
  assign T603 = T604 == T490;
  assign T604 = idxs[6'h26];
  assign T605 = {T617, T606};
  assign T606 = {T612, T607};
  assign T607 = {T610, T608};
  assign T608 = T609 == T490;
  assign T609 = idxs[6'h27];
  assign T610 = T611 == T490;
  assign T611 = idxs[6'h28];
  assign T612 = {T615, T613};
  assign T613 = T614 == T490;
  assign T614 = idxs[6'h29];
  assign T615 = T616 == T490;
  assign T616 = idxs[6'h2a];
  assign T617 = {T623, T618};
  assign T618 = {T621, T619};
  assign T619 = T620 == T490;
  assign T620 = idxs[6'h2b];
  assign T621 = T622 == T490;
  assign T622 = idxs[6'h2c];
  assign T623 = {T626, T624};
  assign T624 = T625 == T490;
  assign T625 = idxs[6'h2d];
  assign T626 = T627 == T490;
  assign T627 = idxs[6'h2e];
  assign T628 = {T652, T629};
  assign T629 = {T641, T630};
  assign T630 = {T636, T631};
  assign T631 = {T634, T632};
  assign T632 = T633 == T490;
  assign T633 = idxs[6'h2f];
  assign T634 = T635 == T490;
  assign T635 = idxs[6'h30];
  assign T636 = {T639, T637};
  assign T637 = T638 == T490;
  assign T638 = idxs[6'h31];
  assign T639 = T640 == T490;
  assign T640 = idxs[6'h32];
  assign T641 = {T647, T642};
  assign T642 = {T645, T643};
  assign T643 = T644 == T490;
  assign T644 = idxs[6'h33];
  assign T645 = T646 == T490;
  assign T646 = idxs[6'h34];
  assign T647 = {T650, T648};
  assign T648 = T649 == T490;
  assign T649 = idxs[6'h35];
  assign T650 = T651 == T490;
  assign T651 = idxs[6'h36];
  assign T652 = {T664, T653};
  assign T653 = {T659, T654};
  assign T654 = {T657, T655};
  assign T655 = T656 == T490;
  assign T656 = idxs[6'h37];
  assign T657 = T658 == T490;
  assign T658 = idxs[6'h38];
  assign T659 = {T662, T660};
  assign T660 = T661 == T490;
  assign T661 = idxs[6'h39];
  assign T662 = T663 == T490;
  assign T663 = idxs[6'h3a];
  assign T664 = {T670, T665};
  assign T665 = {T668, T666};
  assign T666 = T667 == T490;
  assign T667 = idxs[6'h3b];
  assign T668 = T669 == T490;
  assign T669 = idxs[6'h3c];
  assign T670 = T671 == T490;
  assign T671 = idxs[6'h3d];
  assign T1618 = T1619[6'h3d:1'h0];
  assign T1619 = reset ? 64'h0 : T672;
  assign T672 = io_invalidate ? 64'h0 : T673;
  assign T673 = T14 ? T1053 : T1620;
  assign T1620 = {2'h0, T674};
  assign T674 = T14 ? T675 : idxValid;
  assign T675 = idxValid & T676;
  assign T676 = ~ T677;
  assign T677 = T678;
  assign T678 = {T868, T679};
  assign T679 = {T779, T680};
  assign T680 = {T732, T681};
  assign T681 = {T709, T682};
  assign T682 = {T698, T683};
  assign T683 = {T693, T684};
  assign T684 = T685 != 8'h0;
  assign T685 = pageReplEn & T1621;
  assign T1621 = {2'h0, T686};
  assign T686 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T687[3'h5:1'h0];
  assign T687 = 1'h1 << T688;
  assign T688 = tgtPages[6'h0];
  assign T1622 = {T1633, T1623};
  assign T1623 = {T1632, T1624};
  assign T1624 = T1625[1'h1:1'h1];
  assign T1625 = T1631 | T1626;
  assign T1626 = T1627[1'h1:1'h0];
  assign T1627 = T1630 | T1628;
  assign T1628 = T690[2'h3:1'h0];
  assign T690 = usePageHit ? T1629 : tgtPageRepl;
  assign T1629 = {2'h0, pageHit};
  assign T1630 = T690[3'h7:3'h4];
  assign T1631 = T1627[2'h3:2'h2];
  assign T1632 = T1631 != 2'h0;
  assign T1633 = T1630 != 4'h0;
  assign T691 = T7 & T692;
  assign T692 = T54 < 6'h3e;
  assign T693 = T694 != 8'h0;
  assign T694 = pageReplEn & T1634;
  assign T1634 = {2'h0, T695};
  assign T695 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T696[3'h5:1'h0];
  assign T696 = 1'h1 << T697;
  assign T697 = tgtPages[6'h1];
  assign T698 = {T704, T699};
  assign T699 = T700 != 8'h0;
  assign T700 = pageReplEn & T1635;
  assign T1635 = {2'h0, T701};
  assign T701 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T702[3'h5:1'h0];
  assign T702 = 1'h1 << T703;
  assign T703 = tgtPages[6'h2];
  assign T704 = T705 != 8'h0;
  assign T705 = pageReplEn & T1636;
  assign T1636 = {2'h0, T706};
  assign T706 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T707[3'h5:1'h0];
  assign T707 = 1'h1 << T708;
  assign T708 = tgtPages[6'h3];
  assign T709 = {T721, T710};
  assign T710 = {T716, T711};
  assign T711 = T712 != 8'h0;
  assign T712 = pageReplEn & T1637;
  assign T1637 = {2'h0, T713};
  assign T713 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T714[3'h5:1'h0];
  assign T714 = 1'h1 << T715;
  assign T715 = tgtPages[6'h4];
  assign T716 = T717 != 8'h0;
  assign T717 = pageReplEn & T1638;
  assign T1638 = {2'h0, T718};
  assign T718 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T719[3'h5:1'h0];
  assign T719 = 1'h1 << T720;
  assign T720 = tgtPages[6'h5];
  assign T721 = {T727, T722};
  assign T722 = T723 != 8'h0;
  assign T723 = pageReplEn & T1639;
  assign T1639 = {2'h0, T724};
  assign T724 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T725[3'h5:1'h0];
  assign T725 = 1'h1 << T726;
  assign T726 = tgtPages[6'h6];
  assign T727 = T728 != 8'h0;
  assign T728 = pageReplEn & T1640;
  assign T1640 = {2'h0, T729};
  assign T729 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T730[3'h5:1'h0];
  assign T730 = 1'h1 << T731;
  assign T731 = tgtPages[6'h7];
  assign T732 = {T756, T733};
  assign T733 = {T745, T734};
  assign T734 = {T740, T735};
  assign T735 = T736 != 8'h0;
  assign T736 = pageReplEn & T1641;
  assign T1641 = {2'h0, T737};
  assign T737 = idxPagesOH_8 | tgtPagesOH_8;
  assign tgtPagesOH_8 = T738[3'h5:1'h0];
  assign T738 = 1'h1 << T739;
  assign T739 = tgtPages[6'h8];
  assign T740 = T741 != 8'h0;
  assign T741 = pageReplEn & T1642;
  assign T1642 = {2'h0, T742};
  assign T742 = idxPagesOH_9 | tgtPagesOH_9;
  assign tgtPagesOH_9 = T743[3'h5:1'h0];
  assign T743 = 1'h1 << T744;
  assign T744 = tgtPages[6'h9];
  assign T745 = {T751, T746};
  assign T746 = T747 != 8'h0;
  assign T747 = pageReplEn & T1643;
  assign T1643 = {2'h0, T748};
  assign T748 = idxPagesOH_10 | tgtPagesOH_10;
  assign tgtPagesOH_10 = T749[3'h5:1'h0];
  assign T749 = 1'h1 << T750;
  assign T750 = tgtPages[6'ha];
  assign T751 = T752 != 8'h0;
  assign T752 = pageReplEn & T1644;
  assign T1644 = {2'h0, T753};
  assign T753 = idxPagesOH_11 | tgtPagesOH_11;
  assign tgtPagesOH_11 = T754[3'h5:1'h0];
  assign T754 = 1'h1 << T755;
  assign T755 = tgtPages[6'hb];
  assign T756 = {T768, T757};
  assign T757 = {T763, T758};
  assign T758 = T759 != 8'h0;
  assign T759 = pageReplEn & T1645;
  assign T1645 = {2'h0, T760};
  assign T760 = idxPagesOH_12 | tgtPagesOH_12;
  assign tgtPagesOH_12 = T761[3'h5:1'h0];
  assign T761 = 1'h1 << T762;
  assign T762 = tgtPages[6'hc];
  assign T763 = T764 != 8'h0;
  assign T764 = pageReplEn & T1646;
  assign T1646 = {2'h0, T765};
  assign T765 = idxPagesOH_13 | tgtPagesOH_13;
  assign tgtPagesOH_13 = T766[3'h5:1'h0];
  assign T766 = 1'h1 << T767;
  assign T767 = tgtPages[6'hd];
  assign T768 = {T774, T769};
  assign T769 = T770 != 8'h0;
  assign T770 = pageReplEn & T1647;
  assign T1647 = {2'h0, T771};
  assign T771 = idxPagesOH_14 | tgtPagesOH_14;
  assign tgtPagesOH_14 = T772[3'h5:1'h0];
  assign T772 = 1'h1 << T773;
  assign T773 = tgtPages[6'he];
  assign T774 = T775 != 8'h0;
  assign T775 = pageReplEn & T1648;
  assign T1648 = {2'h0, T776};
  assign T776 = idxPagesOH_15 | tgtPagesOH_15;
  assign tgtPagesOH_15 = T777[3'h5:1'h0];
  assign T777 = 1'h1 << T778;
  assign T778 = tgtPages[6'hf];
  assign T779 = {T827, T780};
  assign T780 = {T804, T781};
  assign T781 = {T793, T782};
  assign T782 = {T788, T783};
  assign T783 = T784 != 8'h0;
  assign T784 = pageReplEn & T1649;
  assign T1649 = {2'h0, T785};
  assign T785 = idxPagesOH_16 | tgtPagesOH_16;
  assign tgtPagesOH_16 = T786[3'h5:1'h0];
  assign T786 = 1'h1 << T787;
  assign T787 = tgtPages[6'h10];
  assign T788 = T789 != 8'h0;
  assign T789 = pageReplEn & T1650;
  assign T1650 = {2'h0, T790};
  assign T790 = idxPagesOH_17 | tgtPagesOH_17;
  assign tgtPagesOH_17 = T791[3'h5:1'h0];
  assign T791 = 1'h1 << T792;
  assign T792 = tgtPages[6'h11];
  assign T793 = {T799, T794};
  assign T794 = T795 != 8'h0;
  assign T795 = pageReplEn & T1651;
  assign T1651 = {2'h0, T796};
  assign T796 = idxPagesOH_18 | tgtPagesOH_18;
  assign tgtPagesOH_18 = T797[3'h5:1'h0];
  assign T797 = 1'h1 << T798;
  assign T798 = tgtPages[6'h12];
  assign T799 = T800 != 8'h0;
  assign T800 = pageReplEn & T1652;
  assign T1652 = {2'h0, T801};
  assign T801 = idxPagesOH_19 | tgtPagesOH_19;
  assign tgtPagesOH_19 = T802[3'h5:1'h0];
  assign T802 = 1'h1 << T803;
  assign T803 = tgtPages[6'h13];
  assign T804 = {T816, T805};
  assign T805 = {T811, T806};
  assign T806 = T807 != 8'h0;
  assign T807 = pageReplEn & T1653;
  assign T1653 = {2'h0, T808};
  assign T808 = idxPagesOH_20 | tgtPagesOH_20;
  assign tgtPagesOH_20 = T809[3'h5:1'h0];
  assign T809 = 1'h1 << T810;
  assign T810 = tgtPages[6'h14];
  assign T811 = T812 != 8'h0;
  assign T812 = pageReplEn & T1654;
  assign T1654 = {2'h0, T813};
  assign T813 = idxPagesOH_21 | tgtPagesOH_21;
  assign tgtPagesOH_21 = T814[3'h5:1'h0];
  assign T814 = 1'h1 << T815;
  assign T815 = tgtPages[6'h15];
  assign T816 = {T822, T817};
  assign T817 = T818 != 8'h0;
  assign T818 = pageReplEn & T1655;
  assign T1655 = {2'h0, T819};
  assign T819 = idxPagesOH_22 | tgtPagesOH_22;
  assign tgtPagesOH_22 = T820[3'h5:1'h0];
  assign T820 = 1'h1 << T821;
  assign T821 = tgtPages[6'h16];
  assign T822 = T823 != 8'h0;
  assign T823 = pageReplEn & T1656;
  assign T1656 = {2'h0, T824};
  assign T824 = idxPagesOH_23 | tgtPagesOH_23;
  assign tgtPagesOH_23 = T825[3'h5:1'h0];
  assign T825 = 1'h1 << T826;
  assign T826 = tgtPages[6'h17];
  assign T827 = {T851, T828};
  assign T828 = {T840, T829};
  assign T829 = {T835, T830};
  assign T830 = T831 != 8'h0;
  assign T831 = pageReplEn & T1657;
  assign T1657 = {2'h0, T832};
  assign T832 = idxPagesOH_24 | tgtPagesOH_24;
  assign tgtPagesOH_24 = T833[3'h5:1'h0];
  assign T833 = 1'h1 << T834;
  assign T834 = tgtPages[6'h18];
  assign T835 = T836 != 8'h0;
  assign T836 = pageReplEn & T1658;
  assign T1658 = {2'h0, T837};
  assign T837 = idxPagesOH_25 | tgtPagesOH_25;
  assign tgtPagesOH_25 = T838[3'h5:1'h0];
  assign T838 = 1'h1 << T839;
  assign T839 = tgtPages[6'h19];
  assign T840 = {T846, T841};
  assign T841 = T842 != 8'h0;
  assign T842 = pageReplEn & T1659;
  assign T1659 = {2'h0, T843};
  assign T843 = idxPagesOH_26 | tgtPagesOH_26;
  assign tgtPagesOH_26 = T844[3'h5:1'h0];
  assign T844 = 1'h1 << T845;
  assign T845 = tgtPages[6'h1a];
  assign T846 = T847 != 8'h0;
  assign T847 = pageReplEn & T1660;
  assign T1660 = {2'h0, T848};
  assign T848 = idxPagesOH_27 | tgtPagesOH_27;
  assign tgtPagesOH_27 = T849[3'h5:1'h0];
  assign T849 = 1'h1 << T850;
  assign T850 = tgtPages[6'h1b];
  assign T851 = {T863, T852};
  assign T852 = {T858, T853};
  assign T853 = T854 != 8'h0;
  assign T854 = pageReplEn & T1661;
  assign T1661 = {2'h0, T855};
  assign T855 = idxPagesOH_28 | tgtPagesOH_28;
  assign tgtPagesOH_28 = T856[3'h5:1'h0];
  assign T856 = 1'h1 << T857;
  assign T857 = tgtPages[6'h1c];
  assign T858 = T859 != 8'h0;
  assign T859 = pageReplEn & T1662;
  assign T1662 = {2'h0, T860};
  assign T860 = idxPagesOH_29 | tgtPagesOH_29;
  assign tgtPagesOH_29 = T861[3'h5:1'h0];
  assign T861 = 1'h1 << T862;
  assign T862 = tgtPages[6'h1d];
  assign T863 = T864 != 8'h0;
  assign T864 = pageReplEn & T1663;
  assign T1663 = {2'h0, T865};
  assign T865 = idxPagesOH_30 | tgtPagesOH_30;
  assign tgtPagesOH_30 = T866[3'h5:1'h0];
  assign T866 = 1'h1 << T867;
  assign T867 = tgtPages[6'h1e];
  assign T868 = {T964, T869};
  assign T869 = {T917, T870};
  assign T870 = {T894, T871};
  assign T871 = {T883, T872};
  assign T872 = {T878, T873};
  assign T873 = T874 != 8'h0;
  assign T874 = pageReplEn & T1664;
  assign T1664 = {2'h0, T875};
  assign T875 = idxPagesOH_31 | tgtPagesOH_31;
  assign tgtPagesOH_31 = T876[3'h5:1'h0];
  assign T876 = 1'h1 << T877;
  assign T877 = tgtPages[6'h1f];
  assign T878 = T879 != 8'h0;
  assign T879 = pageReplEn & T1665;
  assign T1665 = {2'h0, T880};
  assign T880 = idxPagesOH_32 | tgtPagesOH_32;
  assign tgtPagesOH_32 = T881[3'h5:1'h0];
  assign T881 = 1'h1 << T882;
  assign T882 = tgtPages[6'h20];
  assign T883 = {T889, T884};
  assign T884 = T885 != 8'h0;
  assign T885 = pageReplEn & T1666;
  assign T1666 = {2'h0, T886};
  assign T886 = idxPagesOH_33 | tgtPagesOH_33;
  assign tgtPagesOH_33 = T887[3'h5:1'h0];
  assign T887 = 1'h1 << T888;
  assign T888 = tgtPages[6'h21];
  assign T889 = T890 != 8'h0;
  assign T890 = pageReplEn & T1667;
  assign T1667 = {2'h0, T891};
  assign T891 = idxPagesOH_34 | tgtPagesOH_34;
  assign tgtPagesOH_34 = T892[3'h5:1'h0];
  assign T892 = 1'h1 << T893;
  assign T893 = tgtPages[6'h22];
  assign T894 = {T906, T895};
  assign T895 = {T901, T896};
  assign T896 = T897 != 8'h0;
  assign T897 = pageReplEn & T1668;
  assign T1668 = {2'h0, T898};
  assign T898 = idxPagesOH_35 | tgtPagesOH_35;
  assign tgtPagesOH_35 = T899[3'h5:1'h0];
  assign T899 = 1'h1 << T900;
  assign T900 = tgtPages[6'h23];
  assign T901 = T902 != 8'h0;
  assign T902 = pageReplEn & T1669;
  assign T1669 = {2'h0, T903};
  assign T903 = idxPagesOH_36 | tgtPagesOH_36;
  assign tgtPagesOH_36 = T904[3'h5:1'h0];
  assign T904 = 1'h1 << T905;
  assign T905 = tgtPages[6'h24];
  assign T906 = {T912, T907};
  assign T907 = T908 != 8'h0;
  assign T908 = pageReplEn & T1670;
  assign T1670 = {2'h0, T909};
  assign T909 = idxPagesOH_37 | tgtPagesOH_37;
  assign tgtPagesOH_37 = T910[3'h5:1'h0];
  assign T910 = 1'h1 << T911;
  assign T911 = tgtPages[6'h25];
  assign T912 = T913 != 8'h0;
  assign T913 = pageReplEn & T1671;
  assign T1671 = {2'h0, T914};
  assign T914 = idxPagesOH_38 | tgtPagesOH_38;
  assign tgtPagesOH_38 = T915[3'h5:1'h0];
  assign T915 = 1'h1 << T916;
  assign T916 = tgtPages[6'h26];
  assign T917 = {T941, T918};
  assign T918 = {T930, T919};
  assign T919 = {T925, T920};
  assign T920 = T921 != 8'h0;
  assign T921 = pageReplEn & T1672;
  assign T1672 = {2'h0, T922};
  assign T922 = idxPagesOH_39 | tgtPagesOH_39;
  assign tgtPagesOH_39 = T923[3'h5:1'h0];
  assign T923 = 1'h1 << T924;
  assign T924 = tgtPages[6'h27];
  assign T925 = T926 != 8'h0;
  assign T926 = pageReplEn & T1673;
  assign T1673 = {2'h0, T927};
  assign T927 = idxPagesOH_40 | tgtPagesOH_40;
  assign tgtPagesOH_40 = T928[3'h5:1'h0];
  assign T928 = 1'h1 << T929;
  assign T929 = tgtPages[6'h28];
  assign T930 = {T936, T931};
  assign T931 = T932 != 8'h0;
  assign T932 = pageReplEn & T1674;
  assign T1674 = {2'h0, T933};
  assign T933 = idxPagesOH_41 | tgtPagesOH_41;
  assign tgtPagesOH_41 = T934[3'h5:1'h0];
  assign T934 = 1'h1 << T935;
  assign T935 = tgtPages[6'h29];
  assign T936 = T937 != 8'h0;
  assign T937 = pageReplEn & T1675;
  assign T1675 = {2'h0, T938};
  assign T938 = idxPagesOH_42 | tgtPagesOH_42;
  assign tgtPagesOH_42 = T939[3'h5:1'h0];
  assign T939 = 1'h1 << T940;
  assign T940 = tgtPages[6'h2a];
  assign T941 = {T953, T942};
  assign T942 = {T948, T943};
  assign T943 = T944 != 8'h0;
  assign T944 = pageReplEn & T1676;
  assign T1676 = {2'h0, T945};
  assign T945 = idxPagesOH_43 | tgtPagesOH_43;
  assign tgtPagesOH_43 = T946[3'h5:1'h0];
  assign T946 = 1'h1 << T947;
  assign T947 = tgtPages[6'h2b];
  assign T948 = T949 != 8'h0;
  assign T949 = pageReplEn & T1677;
  assign T1677 = {2'h0, T950};
  assign T950 = idxPagesOH_44 | tgtPagesOH_44;
  assign tgtPagesOH_44 = T951[3'h5:1'h0];
  assign T951 = 1'h1 << T952;
  assign T952 = tgtPages[6'h2c];
  assign T953 = {T959, T954};
  assign T954 = T955 != 8'h0;
  assign T955 = pageReplEn & T1678;
  assign T1678 = {2'h0, T956};
  assign T956 = idxPagesOH_45 | tgtPagesOH_45;
  assign tgtPagesOH_45 = T957[3'h5:1'h0];
  assign T957 = 1'h1 << T958;
  assign T958 = tgtPages[6'h2d];
  assign T959 = T960 != 8'h0;
  assign T960 = pageReplEn & T1679;
  assign T1679 = {2'h0, T961};
  assign T961 = idxPagesOH_46 | tgtPagesOH_46;
  assign tgtPagesOH_46 = T962[3'h5:1'h0];
  assign T962 = 1'h1 << T963;
  assign T963 = tgtPages[6'h2e];
  assign T964 = {T1012, T965};
  assign T965 = {T989, T966};
  assign T966 = {T978, T967};
  assign T967 = {T973, T968};
  assign T968 = T969 != 8'h0;
  assign T969 = pageReplEn & T1680;
  assign T1680 = {2'h0, T970};
  assign T970 = idxPagesOH_47 | tgtPagesOH_47;
  assign tgtPagesOH_47 = T971[3'h5:1'h0];
  assign T971 = 1'h1 << T972;
  assign T972 = tgtPages[6'h2f];
  assign T973 = T974 != 8'h0;
  assign T974 = pageReplEn & T1681;
  assign T1681 = {2'h0, T975};
  assign T975 = idxPagesOH_48 | tgtPagesOH_48;
  assign tgtPagesOH_48 = T976[3'h5:1'h0];
  assign T976 = 1'h1 << T977;
  assign T977 = tgtPages[6'h30];
  assign T978 = {T984, T979};
  assign T979 = T980 != 8'h0;
  assign T980 = pageReplEn & T1682;
  assign T1682 = {2'h0, T981};
  assign T981 = idxPagesOH_49 | tgtPagesOH_49;
  assign tgtPagesOH_49 = T982[3'h5:1'h0];
  assign T982 = 1'h1 << T983;
  assign T983 = tgtPages[6'h31];
  assign T984 = T985 != 8'h0;
  assign T985 = pageReplEn & T1683;
  assign T1683 = {2'h0, T986};
  assign T986 = idxPagesOH_50 | tgtPagesOH_50;
  assign tgtPagesOH_50 = T987[3'h5:1'h0];
  assign T987 = 1'h1 << T988;
  assign T988 = tgtPages[6'h32];
  assign T989 = {T1001, T990};
  assign T990 = {T996, T991};
  assign T991 = T992 != 8'h0;
  assign T992 = pageReplEn & T1684;
  assign T1684 = {2'h0, T993};
  assign T993 = idxPagesOH_51 | tgtPagesOH_51;
  assign tgtPagesOH_51 = T994[3'h5:1'h0];
  assign T994 = 1'h1 << T995;
  assign T995 = tgtPages[6'h33];
  assign T996 = T997 != 8'h0;
  assign T997 = pageReplEn & T1685;
  assign T1685 = {2'h0, T998};
  assign T998 = idxPagesOH_52 | tgtPagesOH_52;
  assign tgtPagesOH_52 = T999[3'h5:1'h0];
  assign T999 = 1'h1 << T1000;
  assign T1000 = tgtPages[6'h34];
  assign T1001 = {T1007, T1002};
  assign T1002 = T1003 != 8'h0;
  assign T1003 = pageReplEn & T1686;
  assign T1686 = {2'h0, T1004};
  assign T1004 = idxPagesOH_53 | tgtPagesOH_53;
  assign tgtPagesOH_53 = T1005[3'h5:1'h0];
  assign T1005 = 1'h1 << T1006;
  assign T1006 = tgtPages[6'h35];
  assign T1007 = T1008 != 8'h0;
  assign T1008 = pageReplEn & T1687;
  assign T1687 = {2'h0, T1009};
  assign T1009 = idxPagesOH_54 | tgtPagesOH_54;
  assign tgtPagesOH_54 = T1010[3'h5:1'h0];
  assign T1010 = 1'h1 << T1011;
  assign T1011 = tgtPages[6'h36];
  assign T1012 = {T1036, T1013};
  assign T1013 = {T1025, T1014};
  assign T1014 = {T1020, T1015};
  assign T1015 = T1016 != 8'h0;
  assign T1016 = pageReplEn & T1688;
  assign T1688 = {2'h0, T1017};
  assign T1017 = idxPagesOH_55 | tgtPagesOH_55;
  assign tgtPagesOH_55 = T1018[3'h5:1'h0];
  assign T1018 = 1'h1 << T1019;
  assign T1019 = tgtPages[6'h37];
  assign T1020 = T1021 != 8'h0;
  assign T1021 = pageReplEn & T1689;
  assign T1689 = {2'h0, T1022};
  assign T1022 = idxPagesOH_56 | tgtPagesOH_56;
  assign tgtPagesOH_56 = T1023[3'h5:1'h0];
  assign T1023 = 1'h1 << T1024;
  assign T1024 = tgtPages[6'h38];
  assign T1025 = {T1031, T1026};
  assign T1026 = T1027 != 8'h0;
  assign T1027 = pageReplEn & T1690;
  assign T1690 = {2'h0, T1028};
  assign T1028 = idxPagesOH_57 | tgtPagesOH_57;
  assign tgtPagesOH_57 = T1029[3'h5:1'h0];
  assign T1029 = 1'h1 << T1030;
  assign T1030 = tgtPages[6'h39];
  assign T1031 = T1032 != 8'h0;
  assign T1032 = pageReplEn & T1691;
  assign T1691 = {2'h0, T1033};
  assign T1033 = idxPagesOH_58 | tgtPagesOH_58;
  assign tgtPagesOH_58 = T1034[3'h5:1'h0];
  assign T1034 = 1'h1 << T1035;
  assign T1035 = tgtPages[6'h3a];
  assign T1036 = {T1048, T1037};
  assign T1037 = {T1043, T1038};
  assign T1038 = T1039 != 8'h0;
  assign T1039 = pageReplEn & T1692;
  assign T1692 = {2'h0, T1040};
  assign T1040 = idxPagesOH_59 | tgtPagesOH_59;
  assign tgtPagesOH_59 = T1041[3'h5:1'h0];
  assign T1041 = 1'h1 << T1042;
  assign T1042 = tgtPages[6'h3b];
  assign T1043 = T1044 != 8'h0;
  assign T1044 = pageReplEn & T1693;
  assign T1693 = {2'h0, T1045};
  assign T1045 = idxPagesOH_60 | tgtPagesOH_60;
  assign tgtPagesOH_60 = T1046[3'h5:1'h0];
  assign T1046 = 1'h1 << T1047;
  assign T1047 = tgtPages[6'h3c];
  assign T1048 = T1049 != 8'h0;
  assign T1049 = pageReplEn & T1694;
  assign T1694 = {2'h0, T1050};
  assign T1050 = idxPagesOH_61 | tgtPagesOH_61;
  assign tgtPagesOH_61 = T1051[3'h5:1'h0];
  assign T1051 = 1'h1 << T1052;
  assign T1052 = tgtPages[6'h3d];
  assign T1053 = T1060 | T1054;
  assign T1054 = T1696 & T1055;
  assign T1055 = T1057 | T1695;
  assign T1695 = {2'h0, T1056};
  assign T1056 = idxValid ^ idxValid;
  assign T1057 = 1'h1 << T54;
  assign T1696 = T1058 ? 64'hffffffffffffffff : 64'h0;
  assign T1058 = T1059;
  assign T1059 = updateValid;
  assign T1060 = T1697 & T1061;
  assign T1061 = ~ T1055;
  assign T1697 = {2'h0, T674};
  assign T1062 = io_req_valid & T1063;
  assign T1063 = hits != 62'h0;
  assign T1064 = {io_update_bits_taken, T1065};
  assign T1065 = io_update_bits_prediction_bits_bht_history[3'h6:1'h1];
  assign T1066 = T32 & io_update_bits_mispredict;
  assign T1067 = io_req_bits_addr[4'h8:2'h2];
  assign io_resp_bits_bht_history = T1068;
  assign T1068 = R38;
  assign io_resp_bits_entry = T1698;
  assign T1698 = {T1723, T1699};
  assign T1699 = {T1722, T1700};
  assign T1700 = {T1721, T1701};
  assign T1701 = {T1720, T1702};
  assign T1702 = {T1719, T1703};
  assign T1703 = T1704[1'h1:1'h1];
  assign T1704 = T1718 | T1705;
  assign T1705 = T1706[1'h1:1'h0];
  assign T1706 = T1717 | T1707;
  assign T1707 = T1708[2'h3:1'h0];
  assign T1708 = T1716 | T1709;
  assign T1709 = T1710[3'h7:1'h0];
  assign T1710 = T1715 | T1711;
  assign T1711 = T1712[4'hf:1'h0];
  assign T1712 = T1714 | T1713;
  assign T1713 = hits[5'h1f:1'h0];
  assign T1714 = hits[6'h3d:6'h20];
  assign T1715 = T1712[5'h1f:5'h10];
  assign T1716 = T1710[4'hf:4'h8];
  assign T1717 = T1708[3'h7:3'h4];
  assign T1718 = T1706[2'h3:2'h2];
  assign T1719 = T1718 != 2'h0;
  assign T1720 = T1717 != 4'h0;
  assign T1721 = T1716 != 8'h0;
  assign T1722 = T1715 != 16'h0;
  assign T1723 = T1714 != 30'h0;
  assign io_resp_bits_target = T1070;
  assign T1070 = T1581 ? io_update_bits_returnAddr : T1071;
  assign T1071 = T1564 ? T1531 : T1072;
  assign T1072 = {T1323, T1073};
  assign T1073 = T1080 | T1074;
  assign T1074 = T1079 ? T1075 : 13'h0;
  assign T1075 = tgts[6'h3d];
  assign T1724 = io_req_bits_addr[4'hc:1'h0];
  assign T1077 = T7 & T1078;
  assign T1078 = T54 < 6'h3e;
  assign T1079 = hits[6'h3d:6'h3d];
  assign T1080 = T1084 | T1081;
  assign T1081 = T1083 ? T1082 : 13'h0;
  assign T1082 = tgts[6'h3c];
  assign T1083 = hits[6'h3c:6'h3c];
  assign T1084 = T1088 | T1085;
  assign T1085 = T1087 ? T1086 : 13'h0;
  assign T1086 = tgts[6'h3b];
  assign T1087 = hits[6'h3b:6'h3b];
  assign T1088 = T1092 | T1089;
  assign T1089 = T1091 ? T1090 : 13'h0;
  assign T1090 = tgts[6'h3a];
  assign T1091 = hits[6'h3a:6'h3a];
  assign T1092 = T1096 | T1093;
  assign T1093 = T1095 ? T1094 : 13'h0;
  assign T1094 = tgts[6'h39];
  assign T1095 = hits[6'h39:6'h39];
  assign T1096 = T1100 | T1097;
  assign T1097 = T1099 ? T1098 : 13'h0;
  assign T1098 = tgts[6'h38];
  assign T1099 = hits[6'h38:6'h38];
  assign T1100 = T1104 | T1101;
  assign T1101 = T1103 ? T1102 : 13'h0;
  assign T1102 = tgts[6'h37];
  assign T1103 = hits[6'h37:6'h37];
  assign T1104 = T1108 | T1105;
  assign T1105 = T1107 ? T1106 : 13'h0;
  assign T1106 = tgts[6'h36];
  assign T1107 = hits[6'h36:6'h36];
  assign T1108 = T1112 | T1109;
  assign T1109 = T1111 ? T1110 : 13'h0;
  assign T1110 = tgts[6'h35];
  assign T1111 = hits[6'h35:6'h35];
  assign T1112 = T1116 | T1113;
  assign T1113 = T1115 ? T1114 : 13'h0;
  assign T1114 = tgts[6'h34];
  assign T1115 = hits[6'h34:6'h34];
  assign T1116 = T1120 | T1117;
  assign T1117 = T1119 ? T1118 : 13'h0;
  assign T1118 = tgts[6'h33];
  assign T1119 = hits[6'h33:6'h33];
  assign T1120 = T1124 | T1121;
  assign T1121 = T1123 ? T1122 : 13'h0;
  assign T1122 = tgts[6'h32];
  assign T1123 = hits[6'h32:6'h32];
  assign T1124 = T1128 | T1125;
  assign T1125 = T1127 ? T1126 : 13'h0;
  assign T1126 = tgts[6'h31];
  assign T1127 = hits[6'h31:6'h31];
  assign T1128 = T1132 | T1129;
  assign T1129 = T1131 ? T1130 : 13'h0;
  assign T1130 = tgts[6'h30];
  assign T1131 = hits[6'h30:6'h30];
  assign T1132 = T1136 | T1133;
  assign T1133 = T1135 ? T1134 : 13'h0;
  assign T1134 = tgts[6'h2f];
  assign T1135 = hits[6'h2f:6'h2f];
  assign T1136 = T1140 | T1137;
  assign T1137 = T1139 ? T1138 : 13'h0;
  assign T1138 = tgts[6'h2e];
  assign T1139 = hits[6'h2e:6'h2e];
  assign T1140 = T1144 | T1141;
  assign T1141 = T1143 ? T1142 : 13'h0;
  assign T1142 = tgts[6'h2d];
  assign T1143 = hits[6'h2d:6'h2d];
  assign T1144 = T1148 | T1145;
  assign T1145 = T1147 ? T1146 : 13'h0;
  assign T1146 = tgts[6'h2c];
  assign T1147 = hits[6'h2c:6'h2c];
  assign T1148 = T1152 | T1149;
  assign T1149 = T1151 ? T1150 : 13'h0;
  assign T1150 = tgts[6'h2b];
  assign T1151 = hits[6'h2b:6'h2b];
  assign T1152 = T1156 | T1153;
  assign T1153 = T1155 ? T1154 : 13'h0;
  assign T1154 = tgts[6'h2a];
  assign T1155 = hits[6'h2a:6'h2a];
  assign T1156 = T1160 | T1157;
  assign T1157 = T1159 ? T1158 : 13'h0;
  assign T1158 = tgts[6'h29];
  assign T1159 = hits[6'h29:6'h29];
  assign T1160 = T1164 | T1161;
  assign T1161 = T1163 ? T1162 : 13'h0;
  assign T1162 = tgts[6'h28];
  assign T1163 = hits[6'h28:6'h28];
  assign T1164 = T1168 | T1165;
  assign T1165 = T1167 ? T1166 : 13'h0;
  assign T1166 = tgts[6'h27];
  assign T1167 = hits[6'h27:6'h27];
  assign T1168 = T1172 | T1169;
  assign T1169 = T1171 ? T1170 : 13'h0;
  assign T1170 = tgts[6'h26];
  assign T1171 = hits[6'h26:6'h26];
  assign T1172 = T1176 | T1173;
  assign T1173 = T1175 ? T1174 : 13'h0;
  assign T1174 = tgts[6'h25];
  assign T1175 = hits[6'h25:6'h25];
  assign T1176 = T1180 | T1177;
  assign T1177 = T1179 ? T1178 : 13'h0;
  assign T1178 = tgts[6'h24];
  assign T1179 = hits[6'h24:6'h24];
  assign T1180 = T1184 | T1181;
  assign T1181 = T1183 ? T1182 : 13'h0;
  assign T1182 = tgts[6'h23];
  assign T1183 = hits[6'h23:6'h23];
  assign T1184 = T1188 | T1185;
  assign T1185 = T1187 ? T1186 : 13'h0;
  assign T1186 = tgts[6'h22];
  assign T1187 = hits[6'h22:6'h22];
  assign T1188 = T1192 | T1189;
  assign T1189 = T1191 ? T1190 : 13'h0;
  assign T1190 = tgts[6'h21];
  assign T1191 = hits[6'h21:6'h21];
  assign T1192 = T1196 | T1193;
  assign T1193 = T1195 ? T1194 : 13'h0;
  assign T1194 = tgts[6'h20];
  assign T1195 = hits[6'h20:6'h20];
  assign T1196 = T1200 | T1197;
  assign T1197 = T1199 ? T1198 : 13'h0;
  assign T1198 = tgts[6'h1f];
  assign T1199 = hits[5'h1f:5'h1f];
  assign T1200 = T1204 | T1201;
  assign T1201 = T1203 ? T1202 : 13'h0;
  assign T1202 = tgts[6'h1e];
  assign T1203 = hits[5'h1e:5'h1e];
  assign T1204 = T1208 | T1205;
  assign T1205 = T1207 ? T1206 : 13'h0;
  assign T1206 = tgts[6'h1d];
  assign T1207 = hits[5'h1d:5'h1d];
  assign T1208 = T1212 | T1209;
  assign T1209 = T1211 ? T1210 : 13'h0;
  assign T1210 = tgts[6'h1c];
  assign T1211 = hits[5'h1c:5'h1c];
  assign T1212 = T1216 | T1213;
  assign T1213 = T1215 ? T1214 : 13'h0;
  assign T1214 = tgts[6'h1b];
  assign T1215 = hits[5'h1b:5'h1b];
  assign T1216 = T1220 | T1217;
  assign T1217 = T1219 ? T1218 : 13'h0;
  assign T1218 = tgts[6'h1a];
  assign T1219 = hits[5'h1a:5'h1a];
  assign T1220 = T1224 | T1221;
  assign T1221 = T1223 ? T1222 : 13'h0;
  assign T1222 = tgts[6'h19];
  assign T1223 = hits[5'h19:5'h19];
  assign T1224 = T1228 | T1225;
  assign T1225 = T1227 ? T1226 : 13'h0;
  assign T1226 = tgts[6'h18];
  assign T1227 = hits[5'h18:5'h18];
  assign T1228 = T1232 | T1229;
  assign T1229 = T1231 ? T1230 : 13'h0;
  assign T1230 = tgts[6'h17];
  assign T1231 = hits[5'h17:5'h17];
  assign T1232 = T1236 | T1233;
  assign T1233 = T1235 ? T1234 : 13'h0;
  assign T1234 = tgts[6'h16];
  assign T1235 = hits[5'h16:5'h16];
  assign T1236 = T1240 | T1237;
  assign T1237 = T1239 ? T1238 : 13'h0;
  assign T1238 = tgts[6'h15];
  assign T1239 = hits[5'h15:5'h15];
  assign T1240 = T1244 | T1241;
  assign T1241 = T1243 ? T1242 : 13'h0;
  assign T1242 = tgts[6'h14];
  assign T1243 = hits[5'h14:5'h14];
  assign T1244 = T1248 | T1245;
  assign T1245 = T1247 ? T1246 : 13'h0;
  assign T1246 = tgts[6'h13];
  assign T1247 = hits[5'h13:5'h13];
  assign T1248 = T1252 | T1249;
  assign T1249 = T1251 ? T1250 : 13'h0;
  assign T1250 = tgts[6'h12];
  assign T1251 = hits[5'h12:5'h12];
  assign T1252 = T1256 | T1253;
  assign T1253 = T1255 ? T1254 : 13'h0;
  assign T1254 = tgts[6'h11];
  assign T1255 = hits[5'h11:5'h11];
  assign T1256 = T1260 | T1257;
  assign T1257 = T1259 ? T1258 : 13'h0;
  assign T1258 = tgts[6'h10];
  assign T1259 = hits[5'h10:5'h10];
  assign T1260 = T1264 | T1261;
  assign T1261 = T1263 ? T1262 : 13'h0;
  assign T1262 = tgts[6'hf];
  assign T1263 = hits[4'hf:4'hf];
  assign T1264 = T1268 | T1265;
  assign T1265 = T1267 ? T1266 : 13'h0;
  assign T1266 = tgts[6'he];
  assign T1267 = hits[4'he:4'he];
  assign T1268 = T1272 | T1269;
  assign T1269 = T1271 ? T1270 : 13'h0;
  assign T1270 = tgts[6'hd];
  assign T1271 = hits[4'hd:4'hd];
  assign T1272 = T1276 | T1273;
  assign T1273 = T1275 ? T1274 : 13'h0;
  assign T1274 = tgts[6'hc];
  assign T1275 = hits[4'hc:4'hc];
  assign T1276 = T1280 | T1277;
  assign T1277 = T1279 ? T1278 : 13'h0;
  assign T1278 = tgts[6'hb];
  assign T1279 = hits[4'hb:4'hb];
  assign T1280 = T1284 | T1281;
  assign T1281 = T1283 ? T1282 : 13'h0;
  assign T1282 = tgts[6'ha];
  assign T1283 = hits[4'ha:4'ha];
  assign T1284 = T1288 | T1285;
  assign T1285 = T1287 ? T1286 : 13'h0;
  assign T1286 = tgts[6'h9];
  assign T1287 = hits[4'h9:4'h9];
  assign T1288 = T1292 | T1289;
  assign T1289 = T1291 ? T1290 : 13'h0;
  assign T1290 = tgts[6'h8];
  assign T1291 = hits[4'h8:4'h8];
  assign T1292 = T1296 | T1293;
  assign T1293 = T1295 ? T1294 : 13'h0;
  assign T1294 = tgts[6'h7];
  assign T1295 = hits[3'h7:3'h7];
  assign T1296 = T1300 | T1297;
  assign T1297 = T1299 ? T1298 : 13'h0;
  assign T1298 = tgts[6'h6];
  assign T1299 = hits[3'h6:3'h6];
  assign T1300 = T1304 | T1301;
  assign T1301 = T1303 ? T1302 : 13'h0;
  assign T1302 = tgts[6'h5];
  assign T1303 = hits[3'h5:3'h5];
  assign T1304 = T1308 | T1305;
  assign T1305 = T1307 ? T1306 : 13'h0;
  assign T1306 = tgts[6'h4];
  assign T1307 = hits[3'h4:3'h4];
  assign T1308 = T1312 | T1309;
  assign T1309 = T1311 ? T1310 : 13'h0;
  assign T1310 = tgts[6'h3];
  assign T1311 = hits[2'h3:2'h3];
  assign T1312 = T1316 | T1313;
  assign T1313 = T1315 ? T1314 : 13'h0;
  assign T1314 = tgts[6'h2];
  assign T1315 = hits[2'h2:2'h2];
  assign T1316 = T1320 | T1317;
  assign T1317 = T1319 ? T1318 : 13'h0;
  assign T1318 = tgts[6'h1];
  assign T1319 = hits[1'h1:1'h1];
  assign T1320 = T1322 ? T1321 : 13'h0;
  assign T1321 = tgts[6'h0];
  assign T1322 = hits[1'h0:1'h0];
  assign T1323 = T1512 | T1324;
  assign T1324 = T1326 ? T1325 : 30'h0;
  assign T1325 = pages[3'h5];
  assign T1326 = T1327[3'h5:3'h5];
  assign T1327 = T1330 | T1328;
  assign T1328 = T1329 ? tgtPagesOH_61 : 6'h0;
  assign T1329 = hits[6'h3d:6'h3d];
  assign T1330 = T1333 | T1331;
  assign T1331 = T1332 ? tgtPagesOH_60 : 6'h0;
  assign T1332 = hits[6'h3c:6'h3c];
  assign T1333 = T1336 | T1334;
  assign T1334 = T1335 ? tgtPagesOH_59 : 6'h0;
  assign T1335 = hits[6'h3b:6'h3b];
  assign T1336 = T1339 | T1337;
  assign T1337 = T1338 ? tgtPagesOH_58 : 6'h0;
  assign T1338 = hits[6'h3a:6'h3a];
  assign T1339 = T1342 | T1340;
  assign T1340 = T1341 ? tgtPagesOH_57 : 6'h0;
  assign T1341 = hits[6'h39:6'h39];
  assign T1342 = T1345 | T1343;
  assign T1343 = T1344 ? tgtPagesOH_56 : 6'h0;
  assign T1344 = hits[6'h38:6'h38];
  assign T1345 = T1348 | T1346;
  assign T1346 = T1347 ? tgtPagesOH_55 : 6'h0;
  assign T1347 = hits[6'h37:6'h37];
  assign T1348 = T1351 | T1349;
  assign T1349 = T1350 ? tgtPagesOH_54 : 6'h0;
  assign T1350 = hits[6'h36:6'h36];
  assign T1351 = T1354 | T1352;
  assign T1352 = T1353 ? tgtPagesOH_53 : 6'h0;
  assign T1353 = hits[6'h35:6'h35];
  assign T1354 = T1357 | T1355;
  assign T1355 = T1356 ? tgtPagesOH_52 : 6'h0;
  assign T1356 = hits[6'h34:6'h34];
  assign T1357 = T1360 | T1358;
  assign T1358 = T1359 ? tgtPagesOH_51 : 6'h0;
  assign T1359 = hits[6'h33:6'h33];
  assign T1360 = T1363 | T1361;
  assign T1361 = T1362 ? tgtPagesOH_50 : 6'h0;
  assign T1362 = hits[6'h32:6'h32];
  assign T1363 = T1366 | T1364;
  assign T1364 = T1365 ? tgtPagesOH_49 : 6'h0;
  assign T1365 = hits[6'h31:6'h31];
  assign T1366 = T1369 | T1367;
  assign T1367 = T1368 ? tgtPagesOH_48 : 6'h0;
  assign T1368 = hits[6'h30:6'h30];
  assign T1369 = T1372 | T1370;
  assign T1370 = T1371 ? tgtPagesOH_47 : 6'h0;
  assign T1371 = hits[6'h2f:6'h2f];
  assign T1372 = T1375 | T1373;
  assign T1373 = T1374 ? tgtPagesOH_46 : 6'h0;
  assign T1374 = hits[6'h2e:6'h2e];
  assign T1375 = T1378 | T1376;
  assign T1376 = T1377 ? tgtPagesOH_45 : 6'h0;
  assign T1377 = hits[6'h2d:6'h2d];
  assign T1378 = T1381 | T1379;
  assign T1379 = T1380 ? tgtPagesOH_44 : 6'h0;
  assign T1380 = hits[6'h2c:6'h2c];
  assign T1381 = T1384 | T1382;
  assign T1382 = T1383 ? tgtPagesOH_43 : 6'h0;
  assign T1383 = hits[6'h2b:6'h2b];
  assign T1384 = T1387 | T1385;
  assign T1385 = T1386 ? tgtPagesOH_42 : 6'h0;
  assign T1386 = hits[6'h2a:6'h2a];
  assign T1387 = T1390 | T1388;
  assign T1388 = T1389 ? tgtPagesOH_41 : 6'h0;
  assign T1389 = hits[6'h29:6'h29];
  assign T1390 = T1393 | T1391;
  assign T1391 = T1392 ? tgtPagesOH_40 : 6'h0;
  assign T1392 = hits[6'h28:6'h28];
  assign T1393 = T1396 | T1394;
  assign T1394 = T1395 ? tgtPagesOH_39 : 6'h0;
  assign T1395 = hits[6'h27:6'h27];
  assign T1396 = T1399 | T1397;
  assign T1397 = T1398 ? tgtPagesOH_38 : 6'h0;
  assign T1398 = hits[6'h26:6'h26];
  assign T1399 = T1402 | T1400;
  assign T1400 = T1401 ? tgtPagesOH_37 : 6'h0;
  assign T1401 = hits[6'h25:6'h25];
  assign T1402 = T1405 | T1403;
  assign T1403 = T1404 ? tgtPagesOH_36 : 6'h0;
  assign T1404 = hits[6'h24:6'h24];
  assign T1405 = T1408 | T1406;
  assign T1406 = T1407 ? tgtPagesOH_35 : 6'h0;
  assign T1407 = hits[6'h23:6'h23];
  assign T1408 = T1411 | T1409;
  assign T1409 = T1410 ? tgtPagesOH_34 : 6'h0;
  assign T1410 = hits[6'h22:6'h22];
  assign T1411 = T1414 | T1412;
  assign T1412 = T1413 ? tgtPagesOH_33 : 6'h0;
  assign T1413 = hits[6'h21:6'h21];
  assign T1414 = T1417 | T1415;
  assign T1415 = T1416 ? tgtPagesOH_32 : 6'h0;
  assign T1416 = hits[6'h20:6'h20];
  assign T1417 = T1420 | T1418;
  assign T1418 = T1419 ? tgtPagesOH_31 : 6'h0;
  assign T1419 = hits[5'h1f:5'h1f];
  assign T1420 = T1423 | T1421;
  assign T1421 = T1422 ? tgtPagesOH_30 : 6'h0;
  assign T1422 = hits[5'h1e:5'h1e];
  assign T1423 = T1426 | T1424;
  assign T1424 = T1425 ? tgtPagesOH_29 : 6'h0;
  assign T1425 = hits[5'h1d:5'h1d];
  assign T1426 = T1429 | T1427;
  assign T1427 = T1428 ? tgtPagesOH_28 : 6'h0;
  assign T1428 = hits[5'h1c:5'h1c];
  assign T1429 = T1432 | T1430;
  assign T1430 = T1431 ? tgtPagesOH_27 : 6'h0;
  assign T1431 = hits[5'h1b:5'h1b];
  assign T1432 = T1435 | T1433;
  assign T1433 = T1434 ? tgtPagesOH_26 : 6'h0;
  assign T1434 = hits[5'h1a:5'h1a];
  assign T1435 = T1438 | T1436;
  assign T1436 = T1437 ? tgtPagesOH_25 : 6'h0;
  assign T1437 = hits[5'h19:5'h19];
  assign T1438 = T1441 | T1439;
  assign T1439 = T1440 ? tgtPagesOH_24 : 6'h0;
  assign T1440 = hits[5'h18:5'h18];
  assign T1441 = T1444 | T1442;
  assign T1442 = T1443 ? tgtPagesOH_23 : 6'h0;
  assign T1443 = hits[5'h17:5'h17];
  assign T1444 = T1447 | T1445;
  assign T1445 = T1446 ? tgtPagesOH_22 : 6'h0;
  assign T1446 = hits[5'h16:5'h16];
  assign T1447 = T1450 | T1448;
  assign T1448 = T1449 ? tgtPagesOH_21 : 6'h0;
  assign T1449 = hits[5'h15:5'h15];
  assign T1450 = T1453 | T1451;
  assign T1451 = T1452 ? tgtPagesOH_20 : 6'h0;
  assign T1452 = hits[5'h14:5'h14];
  assign T1453 = T1456 | T1454;
  assign T1454 = T1455 ? tgtPagesOH_19 : 6'h0;
  assign T1455 = hits[5'h13:5'h13];
  assign T1456 = T1459 | T1457;
  assign T1457 = T1458 ? tgtPagesOH_18 : 6'h0;
  assign T1458 = hits[5'h12:5'h12];
  assign T1459 = T1462 | T1460;
  assign T1460 = T1461 ? tgtPagesOH_17 : 6'h0;
  assign T1461 = hits[5'h11:5'h11];
  assign T1462 = T1465 | T1463;
  assign T1463 = T1464 ? tgtPagesOH_16 : 6'h0;
  assign T1464 = hits[5'h10:5'h10];
  assign T1465 = T1468 | T1466;
  assign T1466 = T1467 ? tgtPagesOH_15 : 6'h0;
  assign T1467 = hits[4'hf:4'hf];
  assign T1468 = T1471 | T1469;
  assign T1469 = T1470 ? tgtPagesOH_14 : 6'h0;
  assign T1470 = hits[4'he:4'he];
  assign T1471 = T1474 | T1472;
  assign T1472 = T1473 ? tgtPagesOH_13 : 6'h0;
  assign T1473 = hits[4'hd:4'hd];
  assign T1474 = T1477 | T1475;
  assign T1475 = T1476 ? tgtPagesOH_12 : 6'h0;
  assign T1476 = hits[4'hc:4'hc];
  assign T1477 = T1480 | T1478;
  assign T1478 = T1479 ? tgtPagesOH_11 : 6'h0;
  assign T1479 = hits[4'hb:4'hb];
  assign T1480 = T1483 | T1481;
  assign T1481 = T1482 ? tgtPagesOH_10 : 6'h0;
  assign T1482 = hits[4'ha:4'ha];
  assign T1483 = T1486 | T1484;
  assign T1484 = T1485 ? tgtPagesOH_9 : 6'h0;
  assign T1485 = hits[4'h9:4'h9];
  assign T1486 = T1489 | T1487;
  assign T1487 = T1488 ? tgtPagesOH_8 : 6'h0;
  assign T1488 = hits[4'h8:4'h8];
  assign T1489 = T1492 | T1490;
  assign T1490 = T1491 ? tgtPagesOH_7 : 6'h0;
  assign T1491 = hits[3'h7:3'h7];
  assign T1492 = T1495 | T1493;
  assign T1493 = T1494 ? tgtPagesOH_6 : 6'h0;
  assign T1494 = hits[3'h6:3'h6];
  assign T1495 = T1498 | T1496;
  assign T1496 = T1497 ? tgtPagesOH_5 : 6'h0;
  assign T1497 = hits[3'h5:3'h5];
  assign T1498 = T1501 | T1499;
  assign T1499 = T1500 ? tgtPagesOH_4 : 6'h0;
  assign T1500 = hits[3'h4:3'h4];
  assign T1501 = T1504 | T1502;
  assign T1502 = T1503 ? tgtPagesOH_3 : 6'h0;
  assign T1503 = hits[2'h3:2'h3];
  assign T1504 = T1507 | T1505;
  assign T1505 = T1506 ? tgtPagesOH_2 : 6'h0;
  assign T1506 = hits[2'h2:2'h2];
  assign T1507 = T1510 | T1508;
  assign T1508 = T1509 ? tgtPagesOH_1 : 6'h0;
  assign T1509 = hits[1'h1:1'h1];
  assign T1510 = T1511 ? tgtPagesOH_0 : 6'h0;
  assign T1511 = hits[1'h0:1'h0];
  assign T1512 = T1516 | T1513;
  assign T1513 = T1515 ? T1514 : 30'h0;
  assign T1514 = pages[3'h4];
  assign T1515 = T1327[3'h4:3'h4];
  assign T1516 = T1520 | T1517;
  assign T1517 = T1519 ? T1518 : 30'h0;
  assign T1518 = pages[3'h3];
  assign T1519 = T1327[2'h3:2'h3];
  assign T1520 = T1524 | T1521;
  assign T1521 = T1523 ? T1522 : 30'h0;
  assign T1522 = pages[3'h2];
  assign T1523 = T1327[2'h2:2'h2];
  assign T1524 = T1528 | T1525;
  assign T1525 = T1527 ? T1526 : 30'h0;
  assign T1526 = pages[3'h1];
  assign T1527 = T1327[1'h1:1'h1];
  assign T1528 = T1530 ? T1529 : 30'h0;
  assign T1529 = pages[3'h0];
  assign T1530 = T1327[1'h0:1'h0];
  assign T1531 = T1563 ? R1559 : R1532;
  assign T1533 = T1534 ? io_update_bits_returnAddr : R1532;
  assign T1534 = T1558 & T1535;
  assign T1535 = T1536[1'h0:1'h0];
  assign T1536 = 1'h1 << T1537;
  assign T1537 = T1538;
  assign T1538 = R1539 + 1'h1;
  assign T1725 = reset ? 1'h0 : T1540;
  assign T1540 = T1543 ? T1542 : T1541;
  assign T1541 = T1558 ? T1538 : R1539;
  assign T1542 = R1539 - 1'h1;
  assign T1543 = T1554 & T1544;
  assign T1544 = T1545 ^ 1'h1;
  assign T1545 = R1546 == 2'h0;
  assign T1726 = reset ? 2'h0 : T1547;
  assign T1547 = io_invalidate ? 2'h0 : T1548;
  assign T1548 = T1543 ? T1553 : T1549;
  assign T1549 = T1551 ? T1550 : R1546;
  assign T1550 = R1546 + 2'h1;
  assign T1551 = T1558 & T1552;
  assign T1552 = R1546 < 2'h2;
  assign T1553 = R1546 - 2'h1;
  assign T1554 = io_update_valid & T1555;
  assign T1555 = T1557 & T1556;
  assign T1556 = io_update_bits_isReturn & io_update_bits_prediction_valid;
  assign T1557 = io_update_bits_isCall ^ 1'h1;
  assign T1558 = io_update_valid & io_update_bits_isCall;
  assign T1560 = T1561 ? io_update_bits_returnAddr : R1559;
  assign T1561 = T1558 & T1562;
  assign T1562 = T1536[1'h1:1'h1];
  assign T1563 = R1539;
  assign T1564 = T1579 & T1565;
  assign T1565 = T1566 != 62'h0;
  assign T1566 = hits & useRAS;
  assign T1727 = T1567[6'h3d:1'h0];
  assign T1567 = T7 ? T1568 : T1728;
  assign T1728 = {2'h0, useRAS};
  assign T1568 = T1577 | T1569;
  assign T1569 = T1730 & T1570;
  assign T1570 = T1572 | T1729;
  assign T1729 = {2'h0, T1571};
  assign T1571 = useRAS ^ useRAS;
  assign T1572 = 1'h1 << T54;
  assign T1730 = T1573 ? 64'hffffffffffffffff : 64'h0;
  assign T1573 = T1574;
  assign T1574 = R1575;
  assign T1576 = io_update_valid ? io_update_bits_isReturn : R1575;
  assign T1577 = T1731 & T1578;
  assign T1578 = ~ T1570;
  assign T1731 = {2'h0, useRAS};
  assign T1579 = T1580 ^ 1'h1;
  assign T1580 = R1546 == 2'h0;
  assign T1581 = T1558 & T1565;
  assign io_resp_bits_taken = T1582;
  assign T1582 = T1583 ? 1'h0 : io_resp_valid;
  assign T1583 = T1587 & T1584;
  assign T1584 = T1585 ^ 1'h1;
  assign T1585 = T1586 != 62'h0;
  assign T1586 = hits & isJump;
  assign T1587 = T1588 ^ 1'h1;
  assign T1588 = T19[1'h0:1'h0];
  assign io_resp_valid = T1589;
  assign T1589 = hits != 62'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
`endif
    if(io_update_valid) begin
      R4 <= io_update_bits_target;
    end
    if(io_update_valid) begin
      R8 <= io_update_bits_taken;
    end
    if(io_update_valid) begin
      R11 <= io_update_bits_mispredict;
    end
    if(io_update_valid) begin
      updateHit <= io_update_bits_prediction_valid;
    end
    if(reset) begin
      R18 <= 1'h0;
    end else begin
      R18 <= io_update_valid;
    end
    if (T32)
      T21[T35] <= T23;
    if(T1066) begin
      R38 <= T1064;
    end else if(T44) begin
      R38 <= T41;
    end
    isJump <= T1591;
    if(reset) begin
      R55 <= 6'h0;
    end else if(T60) begin
      R55 <= T57;
    end
    if(io_update_valid) begin
      R63 <= io_update_bits_prediction_bits_entry;
    end
    if(io_update_valid) begin
      R67 <= io_update_bits_isJump;
    end
    pageValid <= T1597;
    if(reset) begin
      R88 <= 3'h0;
    end else if(T93) begin
      R88 <= T90;
    end
    if(io_update_valid) begin
      R101 <= io_update_bits_pc;
    end
    if (T110)
      pages[3'h5] <= T105;
    if (T115)
      pages[3'h3] <= T105;
    if (T119)
      pages[3'h1] <= T105;
    if (T126)
      pages[3'h4] <= T123;
    if (T131)
      pages[3'h2] <= T123;
    if (T135)
      pages[3'h0] <= T123;
    if (T180)
      idxPages[T54] <= T1606;
    if (T493)
      idxs[T54] <= T1617;
    idxValid <= T1618;
    if (T691)
      tgtPages[T54] <= T1622;
    if (T1077)
      tgts[T54] <= T1724;
    if(T1534) begin
      R1532 <= io_update_bits_returnAddr;
    end
    if(reset) begin
      R1539 <= 1'h0;
    end else if(T1543) begin
      R1539 <= T1542;
    end else if(T1558) begin
      R1539 <= T1538;
    end
    if(reset) begin
      R1546 <= 2'h0;
    end else if(io_invalidate) begin
      R1546 <= 2'h0;
    end else if(T1543) begin
      R1546 <= T1553;
    end else if(T1551) begin
      R1546 <= T1550;
    end
    if(T1561) begin
      R1559 <= io_update_bits_returnAddr;
    end
    useRAS <= T1727;
    if(io_update_valid) begin
      R1575 <= io_update_bits_isReturn;
    end
  end
endmodule

module FlowThroughSerializer_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T36;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T37;
  wire T4;
  wire T5;
  reg  active;
  wire T38;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire T9;
  wire[3:0] T10;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T39;
  wire[3:0] T11;
  wire[2:0] T12;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T40;
  wire[2:0] T13;
  wire[1:0] T14;
  reg [1:0] rbits_payload_client_xact_id;
  wire[1:0] T41;
  wire[1:0] T15;
  wire[511:0] T16;
  wire[511:0] T17;
  reg [511:0] rbits_payload_data;
  wire[511:0] T42;
  wire[511:0] T18;
  wire[511:0] T43;
  wire[127:0] T19;
  wire[127:0] T20;
  wire[127:0] shifter_0;
  wire[127:0] T21;
  wire[127:0] shifter_1;
  wire[127:0] T22;
  wire T23;
  wire[1:0] T24;
  wire[127:0] T25;
  wire[127:0] shifter_2;
  wire[127:0] T26;
  wire[127:0] shifter_3;
  wire[127:0] T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  reg [1:0] rbits_header_dst;
  wire[1:0] T44;
  wire[1:0] T31;
  wire[1:0] T32;
  reg [1:0] rbits_header_src;
  wire[1:0] T45;
  wire[1:0] T33;
  wire T34;
  wire T35;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cnt = {1{$random}};
    active = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T9 & wrap;
  assign wrap = cnt == 2'h3;
  assign T36 = reset ? 2'h0 : T1;
  assign T1 = T0 ? 2'h0 : T2;
  assign T2 = T9 ? T8 : T3;
  assign T3 = T4 ? T37 : cnt;
  assign T37 = {1'h0, io_out_ready};
  assign T4 = T5 & io_in_valid;
  assign T5 = active ^ 1'h1;
  assign T38 = reset ? 1'h0 : T6;
  assign T6 = T0 ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : active;
  assign T8 = cnt + 2'h1;
  assign T9 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T10;
  assign T10 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T39 = reset ? io_in_bits_payload_g_type : T11;
  assign T11 = T4 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T12;
  assign T12 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T40 = reset ? io_in_bits_payload_master_xact_id : T13;
  assign T13 = T4 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T14;
  assign T14 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T41 = reset ? io_in_bits_payload_client_xact_id : T15;
  assign T15 = T4 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T16;
  assign T16 = active ? T43 : T17;
  assign T17 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T42 = reset ? io_in_bits_payload_data : T18;
  assign T18 = T4 ? io_in_bits_payload_data : rbits_payload_data;
  assign T43 = {384'h0, T19};
  assign T19 = T29 ? T25 : T20;
  assign T20 = T23 ? shifter_1 : shifter_0;
  assign shifter_0 = T21;
  assign T21 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T22;
  assign T22 = rbits_payload_data[8'hff:8'h80];
  assign T23 = T24[1'h0:1'h0];
  assign T24 = cnt;
  assign T25 = T28 ? shifter_3 : shifter_2;
  assign shifter_2 = T26;
  assign T26 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T27;
  assign T27 = rbits_payload_data[9'h1ff:9'h180];
  assign T28 = T24[1'h0:1'h0];
  assign T29 = T24[1'h1:1'h1];
  assign io_out_bits_header_dst = T30;
  assign T30 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T44 = reset ? io_in_bits_header_dst : T31;
  assign T31 = T4 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T32;
  assign T32 = active ? rbits_header_src : io_in_bits_header_src;
  assign T45 = reset ? io_in_bits_header_src : T33;
  assign T33 = T4 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T34;
  assign T34 = active | io_in_valid;
  assign io_in_ready = T35;
  assign T35 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      cnt <= 2'h0;
    end else if(T0) begin
      cnt <= 2'h0;
    end else if(T9) begin
      cnt <= T8;
    end else if(T4) begin
      cnt <= T37;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T0) begin
      active <= 1'h0;
    end else if(T4) begin
      active <= 1'h1;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T4) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T4) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T4) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T4) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T4) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T4) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output io_count
);

  wire T13;
  wire[1:0] T0;
  reg  full;
  wire T14;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[2:0] T3;
  wire[6:0] T4;
  reg [6:0] ram [0:0];
  wire[6:0] T5;
  wire[6:0] T6;
  wire[6:0] T7;
  wire[4:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire empty;
  wire T12;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T13;
  assign T13 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T14 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T3;
  assign T3 = T4[2'h2:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign io_deq_bits_header_dst = T9;
  assign T9 = T4[3'h4:2'h3];
  assign io_deq_bits_header_src = T10;
  assign T10 = T4[3'h6:3'h5];
  assign io_deq_valid = T11;
  assign T11 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [12:0] io_req_bits_idx,
    input [18:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire T209;
  wire T210;
  wire[3:0] T0;
  wire[2:0] T1;
  wire[5:0] T2;
  wire[2:0] T3;
  wire[511:0] T4;
  wire[1:0] T5;
  wire[25:0] T6;
  wire[25:0] T7;
  reg [31:0] s2_addr;
  wire[31:0] T8;
  wire[31:0] s1_addr;
  wire[31:0] T9;
  reg [12:0] s1_pgoff;
  wire[12:0] T10;
  wire T11;
  wire rdy;
  wire T12;
  wire T13;
  wire s2_miss;
  wire T14;
  wire s2_any_tag_hit;
  wire T15;
  wire T16;
  wire T17;
  wire s2_disparity_1;
  wire T18;
  reg  R19;
  wire T20;
  wire T21;
  wire T22;
  wire stall;
  wire T23;
  reg  s1_valid;
  wire T197;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  R29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[6:0] T38;
  wire T39;
  reg [255:0] vb_array;
  wire[255:0] T198;
  wire[255:0] T40;
  wire[255:0] T41;
  wire[255:0] T42;
  wire[255:0] T43;
  wire[255:0] T44;
  wire[255:0] T45;
  wire[255:0] T46;
  wire[7:0] T47;
  wire[6:0] s2_idx;
  wire repl_way;
  reg [15:0] R48;
  wire[15:0] T199;
  wire[15:0] T49;
  wire[15:0] T50;
  wire[14:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[255:0] T200;
  wire T59;
  wire[255:0] T60;
  wire[255:0] T61;
  wire T62;
  wire T63;
  reg  invalidated;
  wire T64;
  wire T65;
  wire T66;
  reg [1:0] state;
  wire[1:0] T201;
  wire[1:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire[255:0] T79;
  wire[255:0] T80;
  wire[255:0] T81;
  wire[7:0] T82;
  wire[255:0] T202;
  wire T83;
  wire[255:0] T84;
  wire[255:0] T85;
  wire T86;
  wire[255:0] T87;
  wire[255:0] T88;
  wire[255:0] T89;
  wire[7:0] T90;
  wire[255:0] T203;
  wire T91;
  wire[255:0] T92;
  wire[255:0] T93;
  wire T94;
  wire s2_disparity_0;
  wire T95;
  reg  R96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg  R101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[7:0] T109;
  wire[6:0] T110;
  wire T111;
  wire T112;
  wire s2_tag_hit_1;
  wire T113;
  reg  R114;
  wire T115;
  wire s1_tag_match_1;
  wire T116;
  wire[18:0] s1_tag;
  wire[18:0] T117;
  wire[18:0] T118;
  wire[37:0] T119;
  wire T133;
  wire s0_valid;
  wire T134;
  wire T135;
  wire[6:0] T131;
  wire[12:0] s0_pgoff;
  wire T132;
  wire[37:0] T120;
  wire[37:0] T121;
  wire[37:0] T122;
  wire[18:0] T123;
  wire[18:0] T204;
  wire T124;
  wire[1:0] T125;
  wire[18:0] T126;
  wire[18:0] T205;
  wire T127;
  wire[37:0] T128;
  wire[18:0] T129;
  wire[18:0] s2_tag;
  reg [6:0] tag_raddr;
  wire[6:0] T130;
  wire s2_tag_hit_0;
  wire T136;
  reg  R137;
  wire T138;
  wire s1_tag_match_0;
  wire T139;
  wire[18:0] T140;
  wire[18:0] T141;
  reg  s2_valid;
  wire T206;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire[127:0] T153;
  wire[127:0] T154;
  reg [127:0] s2_dout_1;
  wire[127:0] T155;
  wire[127:0] T156;
  wire T165;
  wire T166;
  wire T159;
  wire T160;
  wire[8:0] T164;
  wire[127:0] T158;
  wire[127:0] T207;
  wire[8:0] T161;
  reg [8:0] R162;
  wire[8:0] T163;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire[127:0] T171;
  reg [127:0] s2_dout_0;
  wire[127:0] T172;
  wire[127:0] T173;
  wire T182;
  wire T183;
  wire T176;
  wire T177;
  wire[8:0] T181;
  wire[127:0] T175;
  wire[127:0] T208;
  wire[8:0] T178;
  reg [8:0] R179;
  wire[8:0] T180;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire[31:0] T188;
  wire[31:0] T189;
  wire[31:0] s2_dout_word_1;
  wire[127:0] T190;
  wire[6:0] T191;
  wire[1:0] T192;
  wire[5:0] s2_offset;
  wire[31:0] T193;
  wire[31:0] s2_dout_word_0;
  wire[127:0] T194;
  wire[6:0] T195;
  wire[1:0] T196;
  wire s2_hit;
  wire FlowThroughSerializer_1_io_in_ready;
  wire FlowThroughSerializer_1_io_out_valid;
  wire[1:0] FlowThroughSerializer_1_io_out_bits_header_src;
  wire[511:0] FlowThroughSerializer_1_io_out_bits_payload_data;
  wire[2:0] FlowThroughSerializer_1_io_out_bits_payload_master_xact_id;
  wire[3:0] FlowThroughSerializer_1_io_out_bits_payload_g_type;
  wire[1:0] FlowThroughSerializer_1_io_cnt;
  wire FlowThroughSerializer_1_io_done;
  wire ack_q_io_enq_ready;
  wire ack_q_io_deq_valid;
  wire[1:0] ack_q_io_deq_bits_header_src;
  wire[1:0] ack_q_io_deq_bits_header_dst;
  wire[2:0] ack_q_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R19 = {1{$random}};
    s1_valid = {1{$random}};
    R29 = {1{$random}};
    vb_array = {8{$random}};
    R48 = {1{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    R96 = {1{$random}};
    R101 = {1{$random}};
    R114 = {1{$random}};
    tag_raddr = {1{$random}};
    R137 = {1{$random}};
    s2_valid = {1{$random}};
    s2_dout_1 = {4{$random}};
    R162 = {1{$random}};
    s2_dout_0 = {4{$random}};
    R179 = {1{$random}};
  end
`endif

  assign T209 = FlowThroughSerializer_1_io_done & T210;
  assign T210 = FlowThroughSerializer_1_io_out_bits_payload_g_type != 4'h0;
  assign io_mem_finish_bits_payload_master_xact_id = ack_q_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ack_q_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ack_q_io_deq_bits_header_src;
  assign io_mem_finish_valid = ack_q_io_deq_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T0;
  assign T0 = 4'h0;
  assign io_mem_acquire_bits_payload_subword_addr = T1;
  assign T1 = 3'h0;
  assign io_mem_acquire_bits_payload_write_mask = T2;
  assign T2 = 6'h0;
  assign io_mem_acquire_bits_payload_a_type = T3;
  assign T3 = 3'h2;
  assign io_mem_acquire_bits_payload_data = T4;
  assign T4 = 512'h0;
  assign io_mem_acquire_bits_payload_client_xact_id = T5;
  assign T5 = 2'h0;
  assign io_mem_acquire_bits_payload_addr = T6;
  assign T6 = T7;
  assign T7 = s2_addr >> 3'h6;
  assign T8 = T148 ? s1_addr : s2_addr;
  assign s1_addr = T9;
  assign T9 = {io_req_bits_ppn, s1_pgoff};
  assign T10 = T11 ? io_req_bits_idx : s1_pgoff;
  assign T11 = io_req_valid & rdy;
  assign rdy = T12;
  assign T12 = T147 & T13;
  assign T13 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T14;
  assign T14 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T15;
  assign T15 = T112 & T16;
  assign T16 = T17 ^ 1'h1;
  assign T17 = s2_disparity_0 | s2_disparity_1;
  assign s2_disparity_1 = T18;
  assign T18 = R29 & R19;
  assign T20 = T21 ? 1'h0 : R19;
  assign T21 = T23 & T22;
  assign T22 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T23 = s1_valid & rdy;
  assign T197 = reset ? 1'h0 : T24;
  assign T24 = T28 | T25;
  assign T25 = T27 & T26;
  assign T26 = io_req_bits_kill ^ 1'h1;
  assign T27 = s1_valid & stall;
  assign T28 = io_req_valid & rdy;
  assign T30 = T21 ? T31 : R29;
  assign T31 = T32;
  assign T32 = T39 & T33;
  assign T33 = T34 - 1'h1;
  assign T34 = 1'h1 << T35;
  assign T35 = T36 + 8'h1;
  assign T36 = T37 - T37;
  assign T37 = {1'h1, T38};
  assign T38 = s1_pgoff[4'hc:3'h6];
  assign T39 = vb_array >> T37;
  assign T198 = reset ? 256'h0 : T40;
  assign T40 = T94 ? T87 : T41;
  assign T41 = T86 ? T79 : T42;
  assign T42 = io_invalidate ? 256'h0 : T43;
  assign T43 = T62 ? T44 : vb_array;
  assign T44 = T60 | T45;
  assign T45 = T200 & T46;
  assign T46 = 1'h1 << T47;
  assign T47 = {repl_way, s2_idx};
  assign s2_idx = s2_addr[4'hc:3'h6];
  assign repl_way = R48[1'h0:1'h0];
  assign T199 = reset ? 16'h1 : T49;
  assign T49 = s2_miss ? T50 : R48;
  assign T50 = {T52, T51};
  assign T51 = R48[4'hf:1'h1];
  assign T52 = T54 ^ T53;
  assign T53 = R48[3'h5:3'h5];
  assign T54 = T56 ^ T55;
  assign T55 = R48[2'h3:2'h3];
  assign T56 = T58 ^ T57;
  assign T57 = R48[2'h2:2'h2];
  assign T58 = R48[1'h0:1'h0];
  assign T200 = T59 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T59 = 1'h1;
  assign T60 = vb_array & T61;
  assign T61 = ~ T46;
  assign T62 = FlowThroughSerializer_1_io_done & T63;
  assign T63 = invalidated ^ 1'h1;
  assign T64 = T66 ? 1'h0 : T65;
  assign T65 = io_invalidate ? 1'h1 : invalidated;
  assign T66 = 2'h0 == state;
  assign T201 = reset ? 2'h0 : T67;
  assign T67 = T77 ? 2'h0 : T68;
  assign T68 = T75 ? 2'h3 : T69;
  assign T69 = T72 ? 2'h2 : T70;
  assign T70 = T71 ? 2'h1 : state;
  assign T71 = T66 & s2_miss;
  assign T72 = T74 & T73;
  assign T73 = io_mem_acquire_ready & ack_q_io_enq_ready;
  assign T74 = 2'h1 == state;
  assign T75 = T76 & io_mem_grant_valid;
  assign T76 = 2'h2 == state;
  assign T77 = T78 & FlowThroughSerializer_1_io_done;
  assign T78 = 2'h3 == state;
  assign T79 = T84 | T80;
  assign T80 = T202 & T81;
  assign T81 = 1'h1 << T82;
  assign T82 = {1'h0, s2_idx};
  assign T202 = T83 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T83 = 1'h0;
  assign T84 = vb_array & T85;
  assign T85 = ~ T81;
  assign T86 = s2_valid & s2_disparity_0;
  assign T87 = T92 | T88;
  assign T88 = T203 & T89;
  assign T89 = 1'h1 << T90;
  assign T90 = {1'h1, s2_idx};
  assign T203 = T91 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T91 = 1'h0;
  assign T92 = vb_array & T93;
  assign T93 = ~ T89;
  assign T94 = s2_valid & s2_disparity_1;
  assign s2_disparity_0 = T95;
  assign T95 = R101 & R96;
  assign T97 = T98 ? 1'h0 : R96;
  assign T98 = T100 & T99;
  assign T99 = stall ^ 1'h1;
  assign T100 = s1_valid & rdy;
  assign T102 = T98 ? T103 : R101;
  assign T103 = T104;
  assign T104 = T111 & T105;
  assign T105 = T106 - 1'h1;
  assign T106 = 1'h1 << T107;
  assign T107 = T108 + 8'h1;
  assign T108 = T109 - T109;
  assign T109 = {1'h0, T110};
  assign T110 = s1_pgoff[4'hc:3'h6];
  assign T111 = vb_array >> T109;
  assign T112 = s2_tag_hit_0 | s2_tag_hit_1;
  assign s2_tag_hit_1 = T113;
  assign T113 = R29 & R114;
  assign T115 = T21 ? s1_tag_match_1 : R114;
  assign s1_tag_match_1 = T116;
  assign T116 = T117 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hd];
  assign T117 = T118[5'h12:1'h0];
  assign T118 = T119[6'h25:5'h13];
  assign T133 = T135 & s0_valid;
  assign s0_valid = io_req_valid | T134;
  assign T134 = s1_valid & stall;
  assign T135 = FlowThroughSerializer_1_io_done ^ 1'h1;
  assign T131 = s0_pgoff[4'hc:3'h6];
  assign s0_pgoff = T132 ? s1_pgoff : io_req_bits_idx;
  assign T132 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_1_io_done ? s2_idx : T131),
    .RW0E(T133 || FlowThroughSerializer_1_io_done),
    .RW0W(FlowThroughSerializer_1_io_done),
    .RW0I(T128),
    .RW0M(T121),
    .RW0O(T119)
  );
  assign T121 = T122;
  assign T122 = {T126, T123};
  assign T123 = 19'h0 - T204;
  assign T204 = {18'h0, T124};
  assign T124 = T125[1'h0:1'h0];
  assign T125 = 1'h1 << repl_way;
  assign T126 = 19'h0 - T205;
  assign T205 = {18'h0, T127};
  assign T127 = T125[1'h1:1'h1];
  assign T128 = {T129, T129};
  assign T129 = s2_tag;
  assign s2_tag = s2_addr[5'h1f:4'hd];
  assign T130 = T133 ? T131 : tag_raddr;
  assign s2_tag_hit_0 = T136;
  assign T136 = R101 & R137;
  assign T138 = T98 ? s1_tag_match_0 : R137;
  assign s1_tag_match_0 = T139;
  assign T139 = T140 == s1_tag;
  assign T140 = T141[5'h12:1'h0];
  assign T141 = T119[5'h12:1'h0];
  assign T206 = reset ? 1'h0 : T142;
  assign T142 = T144 | T143;
  assign T143 = io_resp_valid & stall;
  assign T144 = T146 & T145;
  assign T145 = io_req_bits_kill ^ 1'h1;
  assign T146 = s1_valid & rdy;
  assign T147 = state == 2'h0;
  assign T148 = T150 & T149;
  assign T149 = stall ^ 1'h1;
  assign T150 = s1_valid & rdy;
  assign io_mem_acquire_valid = T151;
  assign T151 = T152 & ack_q_io_enq_ready;
  assign T152 = state == 2'h1;
  assign io_resp_bits_datablock = T153;
  assign T153 = T171 | T154;
  assign T154 = s2_tag_hit_1 ? s2_dout_1 : 128'h0;
  assign T155 = T167 ? T156 : s2_dout_1;
  assign T165 = T166 & s0_valid;
  assign T166 = T159 ^ 1'h1;
  assign T159 = FlowThroughSerializer_1_io_out_valid & T160;
  assign T160 = repl_way == 1'h1;
  assign T164 = s0_pgoff[4'hc:3'h4];
  ICache_T157 T157 (
    .CLK(clk),
    .RW0A(T159 ? T161 : T164),
    .RW0E(T165 || T159),
    .RW0W(T159),
    .RW0I(T207),
    .RW0O(T156)
  );
  assign T207 = FlowThroughSerializer_1_io_out_bits_payload_data[7'h7f:1'h0];
  assign T161 = {s2_idx, FlowThroughSerializer_1_io_cnt};
  assign T163 = T165 ? T164 : R162;
  assign T167 = T168 & s1_tag_match_1;
  assign T168 = T170 & T169;
  assign T169 = stall ^ 1'h1;
  assign T170 = s1_valid & rdy;
  assign T171 = s2_tag_hit_0 ? s2_dout_0 : 128'h0;
  assign T172 = T184 ? T173 : s2_dout_0;
  assign T182 = T183 & s0_valid;
  assign T183 = T176 ^ 1'h1;
  assign T176 = FlowThroughSerializer_1_io_out_valid & T177;
  assign T177 = repl_way == 1'h0;
  assign T181 = s0_pgoff[4'hc:3'h4];
  ICache_T157 T174 (
    .CLK(clk),
    .RW0A(T176 ? T178 : T181),
    .RW0E(T182 || T176),
    .RW0W(T176),
    .RW0I(T208),
    .RW0O(T173)
  );
  assign T208 = FlowThroughSerializer_1_io_out_bits_payload_data[7'h7f:1'h0];
  assign T178 = {s2_idx, FlowThroughSerializer_1_io_cnt};
  assign T180 = T182 ? T181 : R179;
  assign T184 = T185 & s1_tag_match_0;
  assign T185 = T187 & T186;
  assign T186 = stall ^ 1'h1;
  assign T187 = s1_valid & rdy;
  assign io_resp_bits_data = T188;
  assign T188 = T193 | T189;
  assign T189 = s2_tag_hit_1 ? s2_dout_word_1 : 32'h0;
  assign s2_dout_word_1 = T190[5'h1f:1'h0];
  assign T190 = s2_dout_1 >> T191;
  assign T191 = T192 << 3'h5;
  assign T192 = s2_offset[2'h3:2'h2];
  assign s2_offset = s2_addr[3'h5:1'h0];
  assign T193 = s2_tag_hit_0 ? s2_dout_word_0 : 32'h0;
  assign s2_dout_word_0 = T194[5'h1f:1'h0];
  assign T194 = s2_dout_0 >> T195;
  assign T195 = T196 << 3'h5;
  assign T196 = s2_offset[2'h3:2'h2];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer_1 FlowThroughSerializer_1(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_1_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_1_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_1_io_out_bits_header_src ),
       //.io_out_bits_header_dst(  )
       .io_out_bits_payload_data( FlowThroughSerializer_1_io_out_bits_payload_data ),
       //.io_out_bits_payload_client_xact_id(  )
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_1_io_out_bits_payload_g_type ),
       .io_cnt( FlowThroughSerializer_1_io_cnt ),
       .io_done( FlowThroughSerializer_1_io_done )
  );
  Queue_9 ack_q(.clk(clk), .reset(reset),
       .io_enq_ready( ack_q_io_enq_ready ),
       .io_enq_valid( T209 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( FlowThroughSerializer_1_io_out_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( FlowThroughSerializer_1_io_out_bits_payload_master_xact_id ),
       .io_deq_ready( io_mem_finish_ready ),
       .io_deq_valid( ack_q_io_deq_valid ),
       .io_deq_bits_header_src( ack_q_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ack_q_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ack_q_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ack_q.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(T148) begin
      s2_addr <= s1_addr;
    end
    if(T11) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T21) begin
      R19 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T24;
    end
    if(T21) begin
      R29 <= T31;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else if(T94) begin
      vb_array <= T87;
    end else if(T86) begin
      vb_array <= T79;
    end else if(io_invalidate) begin
      vb_array <= 256'h0;
    end else if(T62) begin
      vb_array <= T44;
    end
    if(reset) begin
      R48 <= 16'h1;
    end else if(s2_miss) begin
      R48 <= T50;
    end
    if(T66) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T77) begin
      state <= 2'h0;
    end else if(T75) begin
      state <= 2'h3;
    end else if(T72) begin
      state <= 2'h2;
    end else if(T71) begin
      state <= 2'h1;
    end
    if(T98) begin
      R96 <= 1'h0;
    end
    if(T98) begin
      R101 <= T103;
    end
    if(T21) begin
      R114 <= s1_tag_match_1;
    end
    if(T133) begin
      tag_raddr <= T131;
    end
    if(T98) begin
      R137 <= s1_tag_match_0;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T142;
    end
    if(T167) begin
      s2_dout_1 <= T156;
    end
    if(T165) begin
      R162 <= T164;
    end
    if(T184) begin
      s2_dout_0 <= T173;
    end
    if(T182) begin
      R179 <= T181;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input  io_clear_hit,
    input [36:0] io_tag,
    output io_hit,
    output[7:0] io_hits,
    output[7:0] io_valid_bits,
    input  io_write,
    input [36:0] io_write_tag,
    input [2:0] io_write_addr
);

  reg [7:0] vb_array;
  wire[7:0] T47;
  wire[7:0] T0;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[7:0] T4;
  wire[7:0] T5;
  wire[7:0] T48;
  wire T6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire T11;
  wire T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[3:0] T15;
  wire[1:0] T16;
  wire hits_0;
  wire T17;
  wire[36:0] T18;
  reg [36:0] cam_tags [7:0];
  wire[36:0] T19;
  wire T20;
  wire hits_1;
  wire T21;
  wire[36:0] T22;
  wire T23;
  wire[1:0] T24;
  wire hits_2;
  wire T25;
  wire[36:0] T26;
  wire T27;
  wire hits_3;
  wire T28;
  wire[36:0] T29;
  wire T30;
  wire[3:0] T31;
  wire[1:0] T32;
  wire hits_4;
  wire T33;
  wire[36:0] T34;
  wire T35;
  wire hits_5;
  wire T36;
  wire[36:0] T37;
  wire T38;
  wire[1:0] T39;
  wire hits_6;
  wire T40;
  wire[36:0] T41;
  wire T42;
  wire hits_7;
  wire T43;
  wire[36:0] T44;
  wire T45;
  wire T46;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
`endif

  assign io_valid_bits = vb_array;
  assign T47 = reset ? 8'h0 : T0;
  assign T0 = T11 ? T9 : T1;
  assign T1 = io_clear ? 8'h0 : T2;
  assign T2 = io_write ? T3 : vb_array;
  assign T3 = T7 | T4;
  assign T4 = T48 & T5;
  assign T5 = 1'h1 << io_write_addr;
  assign T48 = T6 ? 8'hff : 8'h0;
  assign T6 = 1'h1;
  assign T7 = vb_array & T8;
  assign T8 = ~ T5;
  assign T9 = vb_array & T10;
  assign T10 = ~ io_hits;
  assign T11 = T12 & io_clear_hit;
  assign T12 = io_clear ^ 1'h1;
  assign io_hits = T13;
  assign T13 = T14;
  assign T14 = {T31, T15};
  assign T15 = {T24, T16};
  assign T16 = {hits_1, hits_0};
  assign hits_0 = T20 & T17;
  assign T17 = T18 == io_tag;
  assign T18 = cam_tags[3'h0];
  assign T20 = vb_array[1'h0:1'h0];
  assign hits_1 = T23 & T21;
  assign T21 = T22 == io_tag;
  assign T22 = cam_tags[3'h1];
  assign T23 = vb_array[1'h1:1'h1];
  assign T24 = {hits_3, hits_2};
  assign hits_2 = T27 & T25;
  assign T25 = T26 == io_tag;
  assign T26 = cam_tags[3'h2];
  assign T27 = vb_array[2'h2:2'h2];
  assign hits_3 = T30 & T28;
  assign T28 = T29 == io_tag;
  assign T29 = cam_tags[3'h3];
  assign T30 = vb_array[2'h3:2'h3];
  assign T31 = {T39, T32};
  assign T32 = {hits_5, hits_4};
  assign hits_4 = T35 & T33;
  assign T33 = T34 == io_tag;
  assign T34 = cam_tags[3'h4];
  assign T35 = vb_array[3'h4:3'h4];
  assign hits_5 = T38 & T36;
  assign T36 = T37 == io_tag;
  assign T37 = cam_tags[3'h5];
  assign T38 = vb_array[3'h5:3'h5];
  assign T39 = {hits_7, hits_6};
  assign hits_6 = T42 & T40;
  assign T40 = T41 == io_tag;
  assign T41 = cam_tags[3'h6];
  assign T42 = vb_array[3'h6:3'h6];
  assign hits_7 = T45 & T43;
  assign T43 = T44 == io_tag;
  assign T44 = cam_tags[3'h7];
  assign T45 = vb_array[3'h7:3'h7];
  assign io_hit = T46;
  assign T46 = io_hits != 8'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 8'h0;
    end else if(T11) begin
      vb_array <= T9;
    end else if(io_clear) begin
      vb_array <= 8'h0;
    end else if(io_write) begin
      vb_array <= T3;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [30:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    output io_resp_miss,
    output[7:0] io_resp_hit_idx,
    output[18:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[29:0] io_ptw_req_bits,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [18:0] io_ptw_resp_bits_ppn,
    input [5:0] io_ptw_resp_bits_perm,
    input [7:0] io_ptw_status_ip,
    input [7:0] io_ptw_status_im,
    input [6:0] io_ptw_status_zero,
    input  io_ptw_status_er,
    input  io_ptw_status_vm,
    input  io_ptw_status_s64,
    input  io_ptw_status_u64,
    input  io_ptw_status_ef,
    input  io_ptw_status_pei,
    input  io_ptw_status_ei,
    input  io_ptw_status_ps,
    input  io_ptw_status_s,
    input  io_ptw_invalidate,
    input  io_ptw_sret
);

  reg [2:0] r_refill_waddr;
  wire[2:0] T32;
  wire[2:0] repl_waddr;
  wire[2:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[2:0] T38;
  wire[2:0] T39;
  wire T40;
  reg [7:0] R41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[14:0] T46;
  wire[2:0] T47;
  wire T48;
  wire[2:0] T180;
  wire[1:0] T181;
  wire T182;
  wire[1:0] T183;
  wire[1:0] T184;
  wire[3:0] T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[1:0] T188;
  wire T189;
  wire T190;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[10:0] T58;
  wire[7:0] T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire T64;
  wire tlb_hit;
  wire[2:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[1:0] T72;
  wire T73;
  wire[2:0] T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[2:0] T196;
  wire[2:0] T197;
  wire T198;
  wire[7:0] T74;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire has_invalid_entry;
  wire T75;
  wire T2;
  wire tlb_miss;
  wire T3;
  wire bad_va;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[36:0] T212;
  reg [37:0] r_refill_tag;
  wire[37:0] T0;
  wire[37:0] lookup_tag;
  wire[37:0] T1;
  wire T213;
  wire T214;
  reg [1:0] state;
  wire[1:0] T179;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[36:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[29:0] T178;
  wire T9;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[7:0] T27;
  reg [7:0] ux_array;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T205;
  wire T76;
  wire T77;
  wire[5:0] T78;
  wire[5:0] T206;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire T83;
  wire[7:0] T84;
  reg [7:0] sx_array;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T207;
  wire T89;
  wire T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[7:0] T98;
  reg [7:0] uw_array;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T208;
  wire T103;
  wire T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire T107;
  wire[7:0] T108;
  reg [7:0] sw_array;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T209;
  wire T113;
  wire T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[7:0] T122;
  reg [7:0] ur_array;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire[7:0] T210;
  wire T127;
  wire T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire T131;
  wire[7:0] T132;
  reg [7:0] sr_array;
  wire[7:0] T133;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[7:0] T211;
  wire T137;
  wire T138;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[18:0] T141;
  wire[18:0] T142;
  wire[18:0] T143;
  wire[18:0] T144;
  wire[18:0] T145;
  reg [18:0] tag_ram [7:0];
  wire[18:0] T146;
  wire T147;
  wire[18:0] T148;
  wire[18:0] T149;
  wire[18:0] T150;
  wire T151;
  wire[18:0] T152;
  wire[18:0] T153;
  wire[18:0] T154;
  wire T155;
  wire[18:0] T156;
  wire[18:0] T157;
  wire[18:0] T158;
  wire T159;
  wire[18:0] T160;
  wire[18:0] T161;
  wire[18:0] T162;
  wire T163;
  wire[18:0] T164;
  wire[18:0] T165;
  wire[18:0] T166;
  wire T167;
  wire[18:0] T168;
  wire[18:0] T169;
  wire[18:0] T170;
  wire T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire tag_cam_io_hit;
  wire[7:0] tag_cam_io_hits;
  wire[7:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R41 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    ux_array = {1{$random}};
    sx_array = {1{$random}};
    uw_array = {1{$random}};
    sw_array = {1{$random}};
    ur_array = {1{$random}};
    sr_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
`endif

  assign T32 = T2 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T191 : T33;
  assign T33 = T34[2'h2:1'h0];
  assign T34 = {T65, T35};
  assign T35 = T40 & T36;
  assign T36 = T37 - 1'h1;
  assign T37 = 1'h1 << T38;
  assign T38 = T39 + 3'h1;
  assign T39 = T65 - T65;
  assign T40 = R41 >> T65;
  assign T42 = T64 ? T43 : R41;
  assign T43 = T53 | T44;
  assign T44 = T52 ? 8'h0 : T45;
  assign T45 = T46[3'h7:1'h0];
  assign T46 = 8'h1 << T47;
  assign T47 = {T50, T48};
  assign T48 = T180[1'h1:1'h1];
  assign T180 = {T190, T181};
  assign T181 = {T189, T182};
  assign T182 = T183[1'h1:1'h1];
  assign T183 = T188 | T184;
  assign T184 = T185[1'h1:1'h0];
  assign T185 = T187 | T186;
  assign T186 = tag_cam_io_hits[2'h3:1'h0];
  assign T187 = tag_cam_io_hits[3'h7:3'h4];
  assign T188 = T185[2'h3:2'h2];
  assign T189 = T188 != 2'h0;
  assign T190 = T187 != 4'h0;
  assign T50 = {1'h1, T51};
  assign T51 = T180[2'h2:2'h2];
  assign T52 = T180[1'h0:1'h0];
  assign T53 = T55 & T54;
  assign T54 = ~ T45;
  assign T55 = T59 | T56;
  assign T56 = T48 ? 8'h0 : T57;
  assign T57 = T58[3'h7:1'h0];
  assign T58 = 8'h1 << T50;
  assign T59 = T61 & T60;
  assign T60 = ~ T57;
  assign T61 = T63 | T62;
  assign T62 = T51 ? 8'h0 : 8'h2;
  assign T63 = R41 & 8'hfd;
  assign T64 = io_req_valid & tlb_hit;
  assign tlb_hit = io_ptw_status_vm & tag_cam_io_hit;
  assign T65 = {T72, T66};
  assign T66 = T71 & T67;
  assign T67 = T68 - 1'h1;
  assign T68 = 1'h1 << T69;
  assign T69 = T70 + 2'h1;
  assign T70 = T72 - T72;
  assign T71 = R41 >> T72;
  assign T72 = {1'h1, T73};
  assign T73 = R41[1'h1:1'h1];
  assign T191 = T204 ? 1'h0 : T192;
  assign T192 = T203 ? 1'h1 : T193;
  assign T193 = T202 ? 2'h2 : T194;
  assign T194 = T201 ? 2'h3 : T195;
  assign T195 = T200 ? 3'h4 : T196;
  assign T196 = T199 ? 3'h5 : T197;
  assign T197 = T198 ? 3'h6 : 3'h7;
  assign T198 = T74[3'h6:3'h6];
  assign T74 = ~ tag_cam_io_valid_bits;
  assign T199 = T74[3'h5:3'h5];
  assign T200 = T74[3'h4:3'h4];
  assign T201 = T74[2'h3:2'h3];
  assign T202 = T74[2'h2:2'h2];
  assign T203 = T74[1'h1:1'h1];
  assign T204 = T74[1'h0:1'h0];
  assign has_invalid_entry = T75 ^ 1'h1;
  assign T75 = tag_cam_io_valid_bits == 8'hff;
  assign T2 = T8 & tlb_miss;
  assign tlb_miss = T6 & T3;
  assign T3 = bad_va ^ 1'h1;
  assign bad_va = T5 != T4;
  assign T4 = io_req_bits_vpn[5'h1d:5'h1d];
  assign T5 = io_req_bits_vpn[5'h1e:5'h1e];
  assign T6 = io_ptw_status_vm & T7;
  assign T7 = tag_cam_io_hit ^ 1'h1;
  assign T8 = io_req_ready & io_req_valid;
  assign T212 = r_refill_tag[6'h24:1'h0];
  assign T0 = T2 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T1;
  assign T1 = {io_req_bits_asid, io_req_bits_vpn};
  assign T213 = T214 & io_ptw_resp_valid;
  assign T214 = state == 2'h2;
  assign T179 = reset ? 2'h0 : T10;
  assign T10 = io_ptw_resp_valid ? 2'h0 : T11;
  assign T11 = T20 ? 2'h3 : T12;
  assign T12 = T19 ? 2'h3 : T13;
  assign T13 = T18 ? 2'h2 : T14;
  assign T14 = T16 ? 2'h0 : T15;
  assign T15 = T2 ? 2'h1 : state;
  assign T16 = T17 & io_ptw_invalidate;
  assign T17 = state == 2'h1;
  assign T18 = T17 & io_ptw_req_ready;
  assign T19 = T18 & io_ptw_invalidate;
  assign T20 = T21 & io_ptw_invalidate;
  assign T21 = state == 2'h2;
  assign T215 = lookup_tag[6'h24:1'h0];
  assign T216 = T219 & T217;
  assign T217 = io_req_bits_instruction ? io_resp_xcpt_if : T218;
  assign T218 = io_resp_xcpt_ld & io_resp_xcpt_st;
  assign T219 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits = T178;
  assign T178 = r_refill_tag[5'h1d:1'h0];
  assign io_ptw_req_valid = T9;
  assign T9 = state == 2'h1;
  assign io_resp_xcpt_if = T22;
  assign T22 = bad_va | T23;
  assign T23 = tlb_hit & T24;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_ptw_status_s ? T83 : T26;
  assign T26 = T27 != 8'h0;
  assign T27 = ux_array & tag_cam_io_hits;
  assign T28 = io_ptw_resp_valid ? T29 : ux_array;
  assign T29 = T81 | T30;
  assign T30 = T205 & T31;
  assign T31 = 1'h1 << r_refill_waddr;
  assign T205 = T76 ? 8'hff : 8'h0;
  assign T76 = T77;
  assign T77 = T78[2'h2:2'h2];
  assign T78 = T206 & io_ptw_resp_bits_perm;
  assign T206 = T79 ? 6'h3f : 6'h0;
  assign T79 = T80;
  assign T80 = io_ptw_resp_bits_error ^ 1'h1;
  assign T81 = ux_array & T82;
  assign T82 = ~ T31;
  assign T83 = T84 != 8'h0;
  assign T84 = sx_array & tag_cam_io_hits;
  assign T85 = io_ptw_resp_valid ? T86 : sx_array;
  assign T86 = T91 | T87;
  assign T87 = T207 & T88;
  assign T88 = 1'h1 << r_refill_waddr;
  assign T207 = T89 ? 8'hff : 8'h0;
  assign T89 = T90;
  assign T90 = T78[3'h5:3'h5];
  assign T91 = sx_array & T92;
  assign T92 = ~ T88;
  assign io_resp_xcpt_st = T93;
  assign T93 = bad_va | T94;
  assign T94 = tlb_hit & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = io_ptw_status_s ? T107 : T97;
  assign T97 = T98 != 8'h0;
  assign T98 = uw_array & tag_cam_io_hits;
  assign T99 = io_ptw_resp_valid ? T100 : uw_array;
  assign T100 = T105 | T101;
  assign T101 = T208 & T102;
  assign T102 = 1'h1 << r_refill_waddr;
  assign T208 = T103 ? 8'hff : 8'h0;
  assign T103 = T104;
  assign T104 = T78[1'h1:1'h1];
  assign T105 = uw_array & T106;
  assign T106 = ~ T102;
  assign T107 = T108 != 8'h0;
  assign T108 = sw_array & tag_cam_io_hits;
  assign T109 = io_ptw_resp_valid ? T110 : sw_array;
  assign T110 = T115 | T111;
  assign T111 = T209 & T112;
  assign T112 = 1'h1 << r_refill_waddr;
  assign T209 = T113 ? 8'hff : 8'h0;
  assign T113 = T114;
  assign T114 = T78[3'h4:3'h4];
  assign T115 = sw_array & T116;
  assign T116 = ~ T112;
  assign io_resp_xcpt_ld = T117;
  assign T117 = bad_va | T118;
  assign T118 = tlb_hit & T119;
  assign T119 = T120 ^ 1'h1;
  assign T120 = io_ptw_status_s ? T131 : T121;
  assign T121 = T122 != 8'h0;
  assign T122 = ur_array & tag_cam_io_hits;
  assign T123 = io_ptw_resp_valid ? T124 : ur_array;
  assign T124 = T129 | T125;
  assign T125 = T210 & T126;
  assign T126 = 1'h1 << r_refill_waddr;
  assign T210 = T127 ? 8'hff : 8'h0;
  assign T127 = T128;
  assign T128 = T78[1'h0:1'h0];
  assign T129 = ur_array & T130;
  assign T130 = ~ T126;
  assign T131 = T132 != 8'h0;
  assign T132 = sr_array & tag_cam_io_hits;
  assign T133 = io_ptw_resp_valid ? T134 : sr_array;
  assign T134 = T139 | T135;
  assign T135 = T211 & T136;
  assign T136 = 1'h1 << r_refill_waddr;
  assign T211 = T137 ? 8'hff : 8'h0;
  assign T137 = T138;
  assign T138 = T78[2'h3:2'h3];
  assign T139 = sr_array & T140;
  assign T140 = ~ T136;
  assign io_resp_ppn = T141;
  assign T141 = T175 ? T143 : T142;
  assign T142 = io_req_bits_vpn[5'h12:1'h0];
  assign T143 = T148 | T144;
  assign T144 = T147 ? T145 : 19'h0;
  assign T145 = tag_ram[3'h7];
  assign T147 = tag_cam_io_hits[3'h7:3'h7];
  assign T148 = T152 | T149;
  assign T149 = T151 ? T150 : 19'h0;
  assign T150 = tag_ram[3'h6];
  assign T151 = tag_cam_io_hits[3'h6:3'h6];
  assign T152 = T156 | T153;
  assign T153 = T155 ? T154 : 19'h0;
  assign T154 = tag_ram[3'h5];
  assign T155 = tag_cam_io_hits[3'h5:3'h5];
  assign T156 = T160 | T157;
  assign T157 = T159 ? T158 : 19'h0;
  assign T158 = tag_ram[3'h4];
  assign T159 = tag_cam_io_hits[3'h4:3'h4];
  assign T160 = T164 | T161;
  assign T161 = T163 ? T162 : 19'h0;
  assign T162 = tag_ram[3'h3];
  assign T163 = tag_cam_io_hits[2'h3:2'h3];
  assign T164 = T168 | T165;
  assign T165 = T167 ? T166 : 19'h0;
  assign T166 = tag_ram[3'h2];
  assign T167 = tag_cam_io_hits[2'h2:2'h2];
  assign T168 = T172 | T169;
  assign T169 = T171 ? T170 : 19'h0;
  assign T170 = tag_ram[3'h1];
  assign T171 = tag_cam_io_hits[1'h1:1'h1];
  assign T172 = T174 ? T173 : 19'h0;
  assign T173 = tag_ram[3'h0];
  assign T174 = tag_cam_io_hits[1'h0:1'h0];
  assign T175 = io_ptw_status_vm & T176;
  assign T176 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T177;
  assign T177 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( io_ptw_invalidate ),
       .io_clear_hit( T216 ),
       .io_tag( T215 ),
       .io_hit( tag_cam_io_hit ),
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T213 ),
       .io_write_tag( T212 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T2) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T64) begin
      R41 <= T43;
    end
    if(T2) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T20) begin
      state <= 2'h3;
    end else if(T19) begin
      state <= 2'h3;
    end else if(T18) begin
      state <= 2'h2;
    end else if(T16) begin
      state <= 2'h0;
    end else if(T2) begin
      state <= 2'h1;
    end
    if(io_ptw_resp_valid) begin
      ux_array <= T29;
    end
    if(io_ptw_resp_valid) begin
      sx_array <= T86;
    end
    if(io_ptw_resp_valid) begin
      uw_array <= T100;
    end
    if(io_ptw_resp_valid) begin
      sw_array <= T110;
    end
    if(io_ptw_resp_valid) begin
      ur_array <= T124;
    end
    if(io_ptw_resp_valid) begin
      sr_array <= T134;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [43:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[43:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_xcpt_ma,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output[42:0] io_cpu_btb_resp_bits_target,
    output[5:0] io_cpu_btb_resp_bits_entry,
    output[6:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input [42:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_btb_update_bits_pc,
    input [42:0] io_cpu_btb_update_bits_target,
    input [42:0] io_cpu_btb_update_bits_returnAddr,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isCall,
    input  io_cpu_btb_update_bits_isReturn,
    input  io_cpu_btb_update_bits_mispredict,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    input  io_cpu_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[30:0] T38;
  wire[43:0] s1_pc;
  reg [43:0] s1_pc_;
  wire[43:0] T19;
  wire[43:0] T20;
  wire[43:0] npc;
  wire[43:0] T21;
  wire[43:0] predicted_npc;
  wire[43:0] pcp4;
  wire[42:0] T22;
  wire[43:0] pcp4_0;
  wire T23;
  wire T24;
  wire T25;
  wire[43:0] btbTarget;
  wire T26;
  reg [43:0] s2_pc;
  wire[43:0] T36;
  wire[43:0] T18;
  wire T2;
  wire T3;
  wire icmiss;
  wire T4;
  reg  s2_valid;
  wire T33;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire stall;
  wire T9;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg  s1_same_block;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire s0_same_block;
  wire T48;
  wire[43:0] T49;
  wire[43:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[12:0] T59;
  wire[43:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[42:0] T65;
  wire[43:0] T66;
  wire T67;
  wire T68;
  wire T69;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T0;
  wire T1;
  reg [6:0] s2_btb_resp_bits_bht_history;
  wire[6:0] T10;
  reg [5:0] s2_btb_resp_bits_entry;
  wire[5:0] T11;
  reg [42:0] s2_btb_resp_bits_target;
  wire[42:0] T12;
  reg  s2_btb_resp_bits_taken;
  wire T13;
  reg  s2_btb_resp_valid;
  wire T34;
  wire T14;
  reg  s2_xcpt_if;
  wire T35;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire[31:0] T37;
  wire[127:0] T27;
  wire[6:0] T28;
  wire[1:0] T29;
  wire[43:0] T30;
  wire T31;
  wire T32;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire[42:0] btb_io_resp_bits_target;
  wire[5:0] btb_io_resp_bits_entry;
  wire[6:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire tlb_io_resp_miss;
  wire[18:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[29:0] tlb_io_ptw_req_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
`endif

  assign T38 = s1_pc >> 4'hd;
  assign s1_pc = s1_pc_ & 44'hffffffffffe;
  assign T19 = io_cpu_req_valid ? io_cpu_req_bits_pc : T20;
  assign T20 = T8 ? npc : s1_pc_;
  assign npc = T21;
  assign T21 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : pcp4;
  assign pcp4 = {T23, T22};
  assign T22 = pcp4_0[6'h2a:1'h0];
  assign pcp4_0 = s1_pc + 44'h4;
  assign T23 = T25 & T24;
  assign T24 = pcp4_0[6'h2a:6'h2a];
  assign T25 = s1_pc[6'h2a:6'h2a];
  assign btbTarget = {T26, btb_io_resp_bits_target};
  assign T26 = btb_io_resp_bits_target[6'h2a:6'h2a];
  assign T36 = reset ? 44'h2000 : T18;
  assign T18 = T2 ? s1_pc : s2_pc;
  assign T2 = T8 & T3;
  assign T3 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T4;
  assign T4 = icache_io_resp_valid ^ 1'h1;
  assign T33 = reset ? 1'h1 : T5;
  assign T5 = io_cpu_req_valid ? 1'h0 : T6;
  assign T6 = T8 ? T7 : s2_valid;
  assign T7 = icmiss ^ 1'h1;
  assign T8 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T9;
  assign T9 = io_cpu_resp_ready ^ 1'h1;
  assign T39 = T41 & T40;
  assign T40 = icmiss ^ 1'h1;
  assign T41 = stall ^ 1'h1;
  assign T42 = T56 & T43;
  assign T43 = s1_same_block ^ 1'h1;
  assign T44 = io_cpu_req_valid ? 1'h0 : T45;
  assign T45 = T8 ? T46 : s1_same_block;
  assign T46 = s0_same_block & T47;
  assign T47 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T51 & T48;
  assign T48 = T50 == T49;
  assign T49 = s1_pc & 44'h10;
  assign T50 = pcp4 & 44'h10;
  assign T51 = T53 & T52;
  assign T52 = btb_io_resp_bits_taken ^ 1'h1;
  assign T53 = T55 & T54;
  assign T54 = io_cpu_req_valid ^ 1'h1;
  assign T55 = icmiss ^ 1'h1;
  assign T56 = stall ^ 1'h1;
  assign T57 = T58 | icmiss;
  assign T58 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T59 = T60[4'hc:1'h0];
  assign T60 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T61 = T63 & T62;
  assign T62 = s0_same_block ^ 1'h1;
  assign T63 = stall ^ 1'h1;
  assign T64 = io_cpu_invalidate | io_cpu_ptw_invalidate;
  assign T65 = T66[6'h2a:1'h0];
  assign T66 = s1_pc & 44'hffffffffffc;
  assign T67 = T69 & T68;
  assign T68 = icmiss ^ 1'h1;
  assign T69 = stall ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = icache_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = icache_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = icache_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = icache_io_mem_finish_valid;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = icache_io_mem_acquire_bits_payload_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = icache_io_mem_acquire_bits_payload_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = icache_io_mem_acquire_bits_payload_write_mask;
  assign io_mem_acquire_bits_payload_a_type = icache_io_mem_acquire_bits_payload_a_type;
  assign io_mem_acquire_bits_payload_data = icache_io_mem_acquire_bits_payload_data;
  assign io_mem_acquire_bits_payload_client_xact_id = icache_io_mem_acquire_bits_payload_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = icache_io_mem_acquire_bits_payload_addr;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cpu_ptw_req_bits = tlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T0 = T1 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T1 = T2 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T10 = T1 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T11 = T1 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T12 = T1 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T13 = T1 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T34 = reset ? 1'h0 : T14;
  assign T14 = T2 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T35 = reset ? 1'h0 : T15;
  assign T15 = T2 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_xcpt_ma = T16;
  assign T16 = T17 != 2'h0;
  assign T17 = s2_pc[1'h1:1'h0];
  assign io_cpu_resp_bits_data = T37;
  assign T37 = T27[5'h1f:1'h0];
  assign T27 = icache_io_resp_bits_datablock >> T28;
  assign T28 = T29 << 3'h5;
  assign T29 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = T30;
  assign T30 = s2_pc & 44'hffffffffffc;
  assign io_cpu_resp_valid = T31;
  assign T31 = s2_valid & T32;
  assign T32 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T67 ),
       .io_req_bits_addr( T65 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_update_valid( io_cpu_btb_update_valid ),
       .io_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_update_bits_returnAddr( io_cpu_btb_update_bits_returnAddr ),
       .io_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_update_bits_isCall( io_cpu_btb_update_bits_isCall ),
       .io_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_update_bits_mispredict( io_cpu_btb_update_bits_mispredict ),
       .io_invalidate( T64 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T61 ),
       .io_req_bits_idx( T59 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T57 ),
       .io_resp_ready( T42 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T39 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T38 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_resp_miss( tlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits( tlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T8) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 44'h2000;
    end else if(T2) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T8) begin
      s2_valid <= T7;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T8) begin
      s1_same_block <= T46;
    end
    if(T1) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T1) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T1) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T1) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T1) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T2) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T2) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [18:0] io_req_bits_tag,
    input [6:0] io_req_bits_idx,
    input [3:0] io_req_bits_way_en,
    input [1:0] io_req_bits_client_xact_id,
    input [2:0] io_req_bits_master_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output[3:0] io_data_req_bits_way_en,
    output[12:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr,
    output[1:0] io_release_bits_client_xact_id,
    output[2:0] io_release_bits_master_xact_id,
    output[511:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg [511:0] R2;
  wire[511:0] T3;
  wire[511:0] T4;
  wire[383:0] T5;
  wire T6;
  reg  r2_data_req_fired;
  wire T38;
  wire T7;
  reg  r1_data_req_fired;
  wire T39;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  reg  active;
  wire T40;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [2:0] cnt;
  wire[2:0] T41;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  reg [2:0] req_master_xact_id;
  wire[2:0] T26;
  reg [1:0] req_client_xact_id;
  wire[1:0] T27;
  wire[25:0] T28;
  wire[25:0] T29;
  reg [6:0] req_idx;
  wire[6:0] T30;
  reg [18:0] req_tag;
  wire[18:0] T31;
  wire[12:0] T32;
  wire[8:0] T33;
  wire[1:0] T34;
  reg [3:0] req_way_en;
  wire[3:0] T35;
  wire fire;
  wire T36;
  wire T37;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    R2 = {16{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    cnt = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_idx = {1{$random}};
    req_tag = {1{$random}};
    req_way_en = {1{$random}};
  end
`endif

  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_data = R2;
  assign T3 = T6 ? T4 : R2;
  assign T4 = {io_data_resp, T5};
  assign T5 = R2[9'h1ff:8'h80];
  assign T6 = active & r2_data_req_fired;
  assign T38 = reset ? 1'h0 : T7;
  assign T7 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T39 = reset ? 1'h0 : T8;
  assign T8 = T10 ? 1'h1 : T9;
  assign T9 = active ? 1'h0 : r1_data_req_fired;
  assign T10 = active & T11;
  assign T11 = T13 & T12;
  assign T12 = io_meta_read_ready & io_meta_read_valid;
  assign T13 = io_data_req_ready & io_data_req_valid;
  assign T40 = reset ? 1'h0 : T14;
  assign T14 = T1 ? 1'h1 : T15;
  assign T15 = T17 ? T16 : active;
  assign T16 = io_release_ready ^ 1'h1;
  assign T17 = active & T18;
  assign T18 = T23 & T19;
  assign T19 = cnt == 3'h4;
  assign T41 = reset ? 3'h0 : T20;
  assign T20 = T1 ? 3'h0 : T21;
  assign T21 = T10 ? T22 : cnt;
  assign T22 = cnt + 3'h1;
  assign T23 = T25 & T24;
  assign T24 = r2_data_req_fired ^ 1'h1;
  assign T25 = r1_data_req_fired ^ 1'h1;
  assign io_release_bits_master_xact_id = req_master_xact_id;
  assign T26 = T1 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T27 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr = T28;
  assign T28 = T29;
  assign T29 = {req_tag, req_idx};
  assign T30 = T1 ? io_req_bits_idx : req_idx;
  assign T31 = T1 ? io_req_bits_tag : req_tag;
  assign io_release_valid = T17;
  assign io_data_req_bits_addr = T32;
  assign T32 = T33 << 3'h4;
  assign T33 = {req_idx, T34};
  assign T34 = cnt[1'h1:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T35 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T36;
  assign T36 = cnt < 3'h4;
  assign io_meta_read_bits_tag = req_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T37;
  assign T37 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T6) begin
      R2 <= T4;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T10) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T17) begin
      active <= T16;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else if(T1) begin
      cnt <= 3'h0;
    end else if(T10) begin
      cnt <= T22;
    end
    if(T1) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_idx <= io_req_bits_idx;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr,
    input [2:0] io_req_bits_master_xact_id,
    input [1:0] io_req_bits_p_type,
    input [1:0] io_req_bits_client_xact_id,
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr,
    output[1:0] io_rep_bits_client_xact_id,
    output[2:0] io_rep_bits_master_xact_id,
    output[511:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    input [3:0] io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_line_state_state
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  reg [1:0] req_p_type;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [3:0] state;
  wire[3:0] T93;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  reg [1:0] line_state_state;
  wire[1:0] T29;
  wire T30;
  wire hit;
  reg [3:0] way_en;
  wire[3:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  reg [2:0] req_master_xact_id;
  wire[2:0] T50;
  reg [1:0] req_client_xact_id;
  wire[1:0] T51;
  wire[6:0] T94;
  reg [25:0] req_addr;
  wire[25:0] T52;
  wire[18:0] T53;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[18:0] T62;
  wire[6:0] T95;
  wire T63;
  wire[18:0] T64;
  wire[6:0] T96;
  wire T65;
  wire[2:0] T66;
  wire[2:0] T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire[2:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire[511:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[25:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_p_type = {1{$random}};
    state = {1{$random}};
    line_state_state = {1{$random}};
    way_en = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr = {1{$random}};
  end
`endif

  assign io_wb_req_bits_r_type = T0;
  assign T0 = T47 ? T41 : T1;
  assign T1 = T40 ? 3'h4 : T2;
  assign T2 = T39 ? 3'h5 : T3;
  assign T3 = T4 ? 3'h6 : 3'h4;
  assign T4 = req_p_type == 2'h2;
  assign T5 = T6 ? io_req_bits_p_type : req_p_type;
  assign T6 = T7 & io_req_valid;
  assign T7 = state == 4'h1;
  assign T93 = reset ? 4'h1 : T8;
  assign T8 = T38 ? 4'h1 : T9;
  assign T9 = T6 ? 4'h2 : T10;
  assign T10 = T36 ? 4'h3 : T11;
  assign T11 = T35 ? 4'h4 : T12;
  assign T12 = T33 ? 4'h2 : T13;
  assign T13 = T32 ? 4'h5 : T14;
  assign T14 = T30 ? T27 : T15;
  assign T15 = T25 ? 4'h1 : T16;
  assign T16 = T23 ? 4'h7 : T17;
  assign T17 = T21 ? 4'h8 : T18;
  assign T18 = T19 ? 4'h1 : state;
  assign T19 = T20 & io_meta_write_ready;
  assign T20 = state == 4'h8;
  assign T21 = T22 & io_wb_req_ready;
  assign T22 = state == 4'h7;
  assign T23 = T24 & io_wb_req_ready;
  assign T24 = state == 4'h6;
  assign T25 = T26 & io_rep_ready;
  assign T26 = state == 4'h5;
  assign T27 = T28 ? 4'h6 : 4'h8;
  assign T28 = line_state_state == 2'h2;
  assign T29 = T32 ? io_line_state_state : line_state_state;
  assign T30 = T25 & hit;
  assign hit = way_en != 4'h0;
  assign T31 = T32 ? io_way_en : way_en;
  assign T32 = state == 4'h4;
  assign T33 = T32 & T34;
  assign T34 = io_mshr_rdy ^ 1'h1;
  assign T35 = state == 4'h3;
  assign T36 = T37 & io_meta_read_ready;
  assign T37 = state == 4'h2;
  assign T38 = state == 4'h0;
  assign T39 = req_p_type == 2'h1;
  assign T40 = req_p_type == 2'h0;
  assign T41 = T46 ? 3'h1 : T42;
  assign T42 = T45 ? 3'h2 : T43;
  assign T43 = T44 ? 3'h3 : 3'h1;
  assign T44 = req_p_type == 2'h2;
  assign T45 = req_p_type == 2'h1;
  assign T46 = req_p_type == 2'h0;
  assign T47 = T48 == 2'h2;
  assign T48 = hit ? line_state_state : T49;
  assign T49 = 2'h0;
  assign io_wb_req_bits_master_xact_id = req_master_xact_id;
  assign T50 = T6 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_wb_req_bits_client_xact_id = req_client_xact_id;
  assign T51 = T6 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_wb_req_bits_way_en = way_en;
  assign io_wb_req_bits_idx = T94;
  assign T94 = req_addr[3'h6:1'h0];
  assign T52 = T6 ? io_req_bits_addr : req_addr;
  assign io_wb_req_bits_tag = T53;
  assign T53 = req_addr >> 3'h7;
  assign io_wb_req_valid = T54;
  assign T54 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T55;
  assign T55 = T56;
  assign T56 = T61 ? 2'h0 : T57;
  assign T57 = T60 ? 2'h1 : T58;
  assign T58 = T59 ? line_state_state : line_state_state;
  assign T59 = req_p_type == 2'h2;
  assign T60 = req_p_type == 2'h1;
  assign T61 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T62;
  assign T62 = req_addr >> 3'h7;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T95;
  assign T95 = req_addr[3'h6:1'h0];
  assign io_meta_write_valid = T63;
  assign T63 = state == 4'h8;
  assign io_meta_read_bits_tag = T64;
  assign T64 = req_addr >> 3'h7;
  assign io_meta_read_bits_idx = T96;
  assign T96 = req_addr[3'h6:1'h0];
  assign io_meta_read_valid = T65;
  assign T65 = state == 4'h2;
  assign io_rep_bits_r_type = T66;
  assign T66 = T67;
  assign T67 = T80 ? T74 : T68;
  assign T68 = T73 ? 3'h4 : T69;
  assign T69 = T72 ? 3'h5 : T70;
  assign T70 = T71 ? 3'h6 : 3'h4;
  assign T71 = req_p_type == 2'h2;
  assign T72 = req_p_type == 2'h1;
  assign T73 = req_p_type == 2'h0;
  assign T74 = T79 ? 3'h1 : T75;
  assign T75 = T78 ? 3'h2 : T76;
  assign T76 = T77 ? 3'h3 : 3'h1;
  assign T77 = req_p_type == 2'h2;
  assign T78 = req_p_type == 2'h1;
  assign T79 = req_p_type == 2'h0;
  assign T80 = T81 == 2'h2;
  assign T81 = hit ? line_state_state : T82;
  assign T82 = 2'h0;
  assign io_rep_bits_data = T83;
  assign T83 = 512'h0;
  assign io_rep_bits_master_xact_id = T84;
  assign T84 = req_master_xact_id;
  assign io_rep_bits_client_xact_id = T85;
  assign T85 = req_client_xact_id;
  assign io_rep_bits_addr = T86;
  assign T86 = req_addr;
  assign io_rep_valid = T87;
  assign T87 = T91 & T88;
  assign T88 = T89 ^ 1'h1;
  assign T89 = hit & T90;
  assign T90 = line_state_state == 2'h2;
  assign T91 = state == 4'h5;
  assign io_req_ready = T92;
  assign T92 = state == 4'h1;

  always @(posedge clk) begin
    if(T6) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(reset) begin
      state <= 4'h1;
    end else if(T38) begin
      state <= 4'h1;
    end else if(T6) begin
      state <= 4'h2;
    end else if(T36) begin
      state <= 4'h3;
    end else if(T35) begin
      state <= 4'h4;
    end else if(T33) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T30) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T23) begin
      state <= 4'h7;
    end else if(T21) begin
      state <= 4'h8;
    end else if(T19) begin
      state <= 4'h1;
    end
    if(T32) begin
      line_state_state <= io_line_state_state;
    end
    if(T32) begin
      way_en <= io_way_en;
    end
    if(T6) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T6) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T6) begin
      req_addr <= io_req_bits_addr;
    end
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    input [18:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input [18:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[18:0] io_out_bits_tag,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[18:0] T2;
  wire T3;
  wire[6:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T2;
  assign T2 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T3 = T0;
  assign io_out_bits_idx = T4;
  assign T4 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [18:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [18:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[18:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[1:0] T2;
  wire T3;
  wire[18:0] T4;
  wire[3:0] T5;
  wire[6:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T2;
  assign T2 = T3 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T3 = T0;
  assign io_out_bits_data_tag = T4;
  assign T4 = T3 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T5;
  assign T5 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T6;
  assign T6 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_a_type,
    input [5:0] io_in_1_bits_write_mask,
    input [2:0] io_in_1_bits_subword_addr,
    input [3:0] io_in_1_bits_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_a_type,
    input [5:0] io_in_0_bits_write_mask,
    input [2:0] io_in_0_bits_subword_addr,
    input [3:0] io_in_0_bits_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_a_type,
    output[5:0] io_out_bits_write_mask,
    output[2:0] io_out_bits_subword_addr,
    output[3:0] io_out_bits_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[2:0] T6;
  wire[511:0] T7;
  wire[1:0] T8;
  wire[25:0] T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_atomic_opcode = T2;
  assign T2 = T3 ? io_in_1_bits_atomic_opcode : io_in_0_bits_atomic_opcode;
  assign T3 = T0;
  assign io_out_bits_subword_addr = T4;
  assign T4 = T3 ? io_in_1_bits_subword_addr : io_in_0_bits_subword_addr;
  assign io_out_bits_write_mask = T5;
  assign T5 = T3 ? io_in_1_bits_write_mask : io_in_0_bits_write_mask;
  assign io_out_bits_a_type = T6;
  assign T6 = T3 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_data = T7;
  assign T7 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T8;
  assign T8 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T9;
  assign T9 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_payload_master_xact_id = T2;
  assign T2 = T3 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T3 = T0;
  assign io_out_bits_header_dst = T4;
  assign T4 = T3 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T5;
  assign T5 = T3 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T6;
  assign T6 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [18:0] io_in_1_bits_tag,
    input [6:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_master_xact_id,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [18:0] io_in_0_bits_tag,
    input [6:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_master_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[18:0] io_out_bits_tag,
    output[6:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_master_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire[3:0] T6;
  wire[6:0] T7;
  wire[18:0] T8;
  wire T9;
  wire T10;
  wire T11;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_master_xact_id = T4;
  assign T4 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T7;
  assign T7 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_bits_tag = T8;
  assign T8 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_valid = T9;
  assign T9 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_9(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    input [7:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input [7:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[2:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output[7:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[4:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[7:0] T5;
  wire[63:0] T6;
  wire[43:0] T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T2;
  assign T2 = T3 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T3 = T0;
  assign io_out_bits_cmd = T4;
  assign T4 = T3 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T5;
  assign T5 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_data = T6;
  assign T6 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T8;
  assign T8 = T3 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T9;
  assign T9 = T3 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T10;
  assign T10 = T3 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T11;
  assign T11 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_10(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits = T2;
  assign T2 = T3 ? io_in_1_bits : io_in_0_bits;
  assign T3 = T0;
  assign io_out_valid = T4;
  assign T4 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input [7:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[7:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T31;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T32;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[130:0] T11;
  reg [130:0] ram [15:0];
  wire[130:0] T12;
  wire[130:0] T13;
  wire[130:0] T14;
  wire[81:0] T15;
  wire[9:0] T16;
  wire[71:0] T17;
  wire[48:0] T18;
  wire[44:0] T19;
  wire[3:0] T20;
  wire[4:0] T21;
  wire[7:0] T22;
  wire[63:0] T23;
  wire[43:0] T24;
  wire T25;
  wire[2:0] T26;
  wire T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_cmd, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_data, io_enq_bits_tag};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_phys, io_enq_bits_addr};
  assign T20 = {io_enq_bits_kill, io_enq_bits_typ};
  assign io_deq_bits_cmd = T21;
  assign T21 = T11[4'h9:3'h5];
  assign io_deq_bits_tag = T22;
  assign T22 = T11[5'h11:4'ha];
  assign io_deq_bits_data = T23;
  assign T23 = T11[7'h51:5'h12];
  assign io_deq_bits_addr = T24;
  assign T24 = T11[7'h7d:7'h52];
  assign io_deq_bits_phys = T25;
  assign T25 = T11[7'h7e:7'h7e];
  assign io_deq_bits_typ = T26;
  assign T26 = T11[8'h81:7'h7f];
  assign io_deq_bits_kill = T27;
  assign T27 = T11[8'h82:8'h82];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[18:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T198;
  wire can_finish;
  wire T77;
  reg [3:0] state;
  wire[3:0] T194;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire refill_done;
  wire T28;
  reg [1:0] refill_count;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire reply;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T78;
  wire T79;
  wire T80;
  wire T199;
  wire T200;
  wire T201;
  wire wb_done;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T82;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire sec_rdy;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire idx_match;
  wire[6:0] T70;
  wire[6:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T71;
  wire T215;
  wire T0;
  wire T1;
  wire T2;
  reg [1:0] meta_hazard;
  wire[1:0] T193;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg [3:0] req_way_en;
  wire[3:0] T72;
  reg [18:0] req_old_meta_tag;
  wire[18:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire[4:0] T81;
  wire[43:0] T195;
  wire[31:0] T83;
  wire[31:0] T84;
  wire[12:0] T85;
  wire[5:0] T86;
  wire T87;
  wire T88;
  wire[1:0] T89;
  reg [1:0] line_state_state;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[1:0] meta_on_flush_state;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[127:0] T196;
  reg [63:0] req_data;
  wire[63:0] T112;
  wire[12:0] T113;
  wire[8:0] T114;
  reg [2:0] acquire_type;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire[2:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire[25:0] T142;
  wire[25:0] T143;
  wire T144;
  wire T145;
  wire[18:0] T197;
  wire[30:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire T192;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[2:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[63:0] rpq_io_deq_bits_data;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T198 = io_mem_finish_ready & can_finish;
  assign can_finish = T78 | T77;
  assign T77 = state == 4'h5;
  assign T194 = reset ? 4'h0 : T10;
  assign T10 = T64 ? T62 : T11;
  assign T11 = T60 ? 4'h4 : T12;
  assign T12 = T42 ? 4'h6 : T13;
  assign T13 = T41 ? 4'h2 : T14;
  assign T14 = T39 ? 4'h3 : T15;
  assign T15 = T37 ? 4'h4 : T16;
  assign T16 = T36 ? 4'h5 : T17;
  assign T17 = T27 ? 4'h6 : T18;
  assign T18 = T25 ? 4'h7 : T19;
  assign T19 = T24 ? 4'h8 : T20;
  assign T20 = T21 ? 4'h0 : state;
  assign T21 = T23 & T22;
  assign T22 = rpq_io_deq_valid ^ 1'h1;
  assign T23 = state == 4'h8;
  assign T24 = state == 4'h7;
  assign T25 = T26 & io_meta_write_ready;
  assign T26 = state == 4'h6;
  assign T27 = T35 & refill_done;
  assign refill_done = reply & T28;
  assign T28 = refill_count == 2'h3;
  assign T29 = T33 ? 2'h0 : T30;
  assign T30 = T32 ? T31 : refill_count;
  assign T31 = refill_count + 2'h1;
  assign T32 = T35 & reply;
  assign T33 = io_req_pri_val & io_req_pri_rdy;
  assign reply = io_mem_grant_valid & T34;
  assign T34 = io_mem_grant_bits_payload_client_xact_id == 2'h0;
  assign T35 = state == 4'h5;
  assign T36 = io_mem_req_ready & io_mem_req_valid;
  assign T37 = T38 & io_meta_write_ready;
  assign T38 = state == 4'h3;
  assign T39 = T40 & reply;
  assign T40 = state == 4'h2;
  assign T41 = io_wb_req_ready & io_wb_req_valid;
  assign T42 = T59 & T43;
  assign T43 = T48 ? T47 : T44;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T46 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T47 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T33 & io_req_bits_tag_match;
  assign T60 = T59 & T61;
  assign T61 = T43 ^ 1'h1;
  assign T62 = T63 ? 4'h1 : 4'h3;
  assign T63 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T64 = T33 & T65;
  assign T65 = io_req_bits_tag_match ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = state == 4'h4;
  assign T80 = state == 4'h0;
  assign T199 = T201 & T200;
  assign T200 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T201 = wb_done | refill_done;
  assign wb_done = reply & T202;
  assign T202 = state == 4'h2;
  assign T203 = T82 ? 1'h0 : T204;
  assign T204 = T206 | T205;
  assign T205 = state == 4'h0;
  assign T206 = io_replay_ready & T207;
  assign T207 = state == 4'h8;
  assign T82 = io_meta_read_ready ^ 1'h1;
  assign T208 = T213 & T209;
  assign T209 = T210 ^ 1'h1;
  assign T210 = T212 | T211;
  assign T211 = io_req_bits_cmd == 5'h3;
  assign T212 = io_req_bits_cmd == 5'h2;
  assign T213 = T215 | T214;
  assign T214 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T150;
  assign T150 = T187 | T151;
  assign T151 = T184 & T152;
  assign T152 = T153 ^ 1'h1;
  assign T153 = T167 | T154;
  assign T154 = T156 & T155;
  assign T155 = io_mem_req_bits_a_type != 3'h1;
  assign T156 = T158 | T157;
  assign T157 = io_req_bits_cmd == 5'h6;
  assign T158 = T160 | T159;
  assign T159 = io_req_bits_cmd == 5'h3;
  assign T160 = T164 | T161;
  assign T161 = T163 | T162;
  assign T162 = io_req_bits_cmd == 5'h4;
  assign T163 = io_req_bits_cmd[2'h3:2'h3];
  assign T164 = T166 | T165;
  assign T165 = io_req_bits_cmd == 5'h7;
  assign T166 = io_req_bits_cmd == 5'h1;
  assign T167 = T177 & T168;
  assign T168 = T170 | T169;
  assign T169 = 3'h6 == io_mem_req_bits_a_type;
  assign T170 = T172 | T171;
  assign T171 = 3'h5 == io_mem_req_bits_a_type;
  assign T172 = T174 | T173;
  assign T173 = 3'h4 == io_mem_req_bits_a_type;
  assign T174 = T176 | T175;
  assign T175 = 3'h3 == io_mem_req_bits_a_type;
  assign T176 = 3'h2 == io_mem_req_bits_a_type;
  assign T177 = T181 | T178;
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h4;
  assign T180 = io_req_bits_cmd[2'h3:2'h3];
  assign T181 = T183 | T182;
  assign T182 = io_req_bits_cmd == 5'h6;
  assign T183 = io_req_bits_cmd == 5'h0;
  assign T184 = T186 | T185;
  assign T185 = state == 4'h5;
  assign T186 = state == 4'h4;
  assign T187 = T189 | T188;
  assign T188 = state == 4'h3;
  assign T189 = T191 | T190;
  assign T190 = state == 4'h2;
  assign T191 = state == 4'h1;
  assign idx_match = req_idx == T70;
  assign T70 = io_req_bits_addr[4'hc:3'h6];
  assign req_idx = req_addr[4'hc:3'h6];
  assign T71 = T33 ? io_req_bits_addr : req_addr;
  assign T215 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T0;
  assign T0 = T69 | T1;
  assign T1 = T8 & T2;
  assign T2 = meta_hazard == 2'h0;
  assign T193 = reset ? 2'h0 : T3;
  assign T3 = T7 ? 2'h1 : T4;
  assign T4 = T6 ? T5 : meta_hazard;
  assign T5 = meta_hazard + 2'h1;
  assign T6 = meta_hazard != 2'h0;
  assign T7 = io_meta_write_ready & io_meta_write_valid;
  assign T8 = T66 & T9;
  assign T9 = state != 4'h3;
  assign T66 = T68 & T67;
  assign T67 = state != 4'h2;
  assign T68 = state != 4'h1;
  assign T69 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h0;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T72 = T33 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T73 = T33 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T74;
  assign T74 = T75 & ackq_io_enq_ready;
  assign T75 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T76;
  assign T76 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T81;
  assign T81 = T82 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T195;
  assign T195 = {12'h0, T83};
  assign T83 = T84;
  assign T84 = {io_tag, T85};
  assign T85 = {req_idx, T86};
  assign T86 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T87;
  assign T87 = T88 & rpq_io_deq_valid;
  assign T88 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T89;
  assign T89 = T107 ? meta_on_flush_state : line_state_state;
  assign T90 = T42 ? meta_on_hit_state : T91;
  assign T91 = T33 ? meta_on_flush_state : T92;
  assign T92 = T32 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T93;
  assign T93 = T98 ? 2'h1 : T94;
  assign T94 = T97 ? 2'h2 : T95;
  assign T95 = T96 ? 2'h2 : 2'h0;
  assign T96 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T97 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T98 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_hit_state = T99;
  assign T99 = T100 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T107 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T108;
  assign T108 = T110 | T109;
  assign T109 = state == 4'h3;
  assign T110 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T111;
  assign T111 = state == 4'h8;
  assign io_mem_resp_data = T196;
  assign T196 = {64'h0, req_data};
  assign T112 = T33 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T113;
  assign T113 = T114 << 3'h4;
  assign T114 = {req_idx, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T115 = T33 ? T130 : T116;
  assign T116 = T129 ? T117 : acquire_type;
  assign T117 = T118 ? 3'h1 : io_mem_req_bits_a_type;
  assign T118 = T120 | T119;
  assign T119 = io_req_bits_cmd == 5'h6;
  assign T120 = T122 | T121;
  assign T121 = io_req_bits_cmd == 5'h3;
  assign T122 = T126 | T123;
  assign T123 = T125 | T124;
  assign T124 = io_req_bits_cmd == 5'h4;
  assign T125 = io_req_bits_cmd[2'h3:2'h3];
  assign T126 = T128 | T127;
  assign T127 = io_req_bits_cmd == 5'h7;
  assign T128 = io_req_bits_cmd == 5'h1;
  assign T129 = io_req_sec_val & io_req_sec_rdy;
  assign T130 = T131 ? 3'h1 : 3'h0;
  assign T131 = T133 | T132;
  assign T132 = io_req_bits_cmd == 5'h6;
  assign T133 = T135 | T134;
  assign T134 = io_req_bits_cmd == 5'h3;
  assign T135 = T139 | T136;
  assign T136 = T138 | T137;
  assign T137 = io_req_bits_cmd == 5'h4;
  assign T138 = io_req_bits_cmd[2'h3:2'h3];
  assign T139 = T141 | T140;
  assign T140 = io_req_bits_cmd == 5'h7;
  assign T141 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 2'h0;
  assign io_mem_req_bits_addr = T142;
  assign T142 = T143;
  assign T143 = {io_tag, req_idx};
  assign io_mem_req_valid = T144;
  assign T144 = T145 & ackq_io_enq_ready;
  assign T145 = state == 4'h4;
  assign io_tag = T197;
  assign T197 = T146[5'h12:1'h0];
  assign T146 = req_addr >> 4'hd;
  assign io_idx_match = T147;
  assign T147 = T148 & idx_match;
  assign T148 = state != 4'h0;
  assign io_req_sec_rdy = T149;
  assign T149 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T192;
  assign T192 = state == 4'h0;
  Queue_12 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T208 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T203 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_9 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T199 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T198 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T64) begin
      state <= T62;
    end else if(T60) begin
      state <= 4'h4;
    end else if(T42) begin
      state <= 4'h6;
    end else if(T41) begin
      state <= 4'h2;
    end else if(T39) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= 4'h5;
    end else if(T27) begin
      state <= 4'h6;
    end else if(T25) begin
      state <= 4'h7;
    end else if(T24) begin
      state <= 4'h8;
    end else if(T21) begin
      state <= 4'h0;
    end
    if(T33) begin
      refill_count <= 2'h0;
    end else if(T32) begin
      refill_count <= T31;
    end
    if(T33) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T7) begin
      meta_hazard <= 2'h1;
    end else if(T6) begin
      meta_hazard <= T5;
    end
    if(T33) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T33) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T42) begin
      line_state_state <= meta_on_hit_state;
    end else if(T33) begin
      line_state_state <= meta_on_flush_state;
    end else if(T32) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T33) begin
      req_data <= io_req_bits_data;
    end
    if(T33) begin
      acquire_type <= T130;
    end else if(T129) begin
      acquire_type <= T117;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[18:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T198;
  wire can_finish;
  wire T77;
  reg [3:0] state;
  wire[3:0] T194;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire refill_done;
  wire T28;
  reg [1:0] refill_count;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire reply;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T78;
  wire T79;
  wire T80;
  wire T199;
  wire T200;
  wire T201;
  wire wb_done;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T82;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire sec_rdy;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire idx_match;
  wire[6:0] T70;
  wire[6:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T71;
  wire T215;
  wire T0;
  wire T1;
  wire T2;
  reg [1:0] meta_hazard;
  wire[1:0] T193;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg [3:0] req_way_en;
  wire[3:0] T72;
  reg [18:0] req_old_meta_tag;
  wire[18:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire[4:0] T81;
  wire[43:0] T195;
  wire[31:0] T83;
  wire[31:0] T84;
  wire[12:0] T85;
  wire[5:0] T86;
  wire T87;
  wire T88;
  wire[1:0] T89;
  reg [1:0] line_state_state;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[1:0] meta_on_flush_state;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[127:0] T196;
  reg [63:0] req_data;
  wire[63:0] T112;
  wire[12:0] T113;
  wire[8:0] T114;
  reg [2:0] acquire_type;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire[2:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire[25:0] T142;
  wire[25:0] T143;
  wire T144;
  wire T145;
  wire[18:0] T197;
  wire[30:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire T192;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[2:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[63:0] rpq_io_deq_bits_data;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T198 = io_mem_finish_ready & can_finish;
  assign can_finish = T78 | T77;
  assign T77 = state == 4'h5;
  assign T194 = reset ? 4'h0 : T10;
  assign T10 = T64 ? T62 : T11;
  assign T11 = T60 ? 4'h4 : T12;
  assign T12 = T42 ? 4'h6 : T13;
  assign T13 = T41 ? 4'h2 : T14;
  assign T14 = T39 ? 4'h3 : T15;
  assign T15 = T37 ? 4'h4 : T16;
  assign T16 = T36 ? 4'h5 : T17;
  assign T17 = T27 ? 4'h6 : T18;
  assign T18 = T25 ? 4'h7 : T19;
  assign T19 = T24 ? 4'h8 : T20;
  assign T20 = T21 ? 4'h0 : state;
  assign T21 = T23 & T22;
  assign T22 = rpq_io_deq_valid ^ 1'h1;
  assign T23 = state == 4'h8;
  assign T24 = state == 4'h7;
  assign T25 = T26 & io_meta_write_ready;
  assign T26 = state == 4'h6;
  assign T27 = T35 & refill_done;
  assign refill_done = reply & T28;
  assign T28 = refill_count == 2'h3;
  assign T29 = T33 ? 2'h0 : T30;
  assign T30 = T32 ? T31 : refill_count;
  assign T31 = refill_count + 2'h1;
  assign T32 = T35 & reply;
  assign T33 = io_req_pri_val & io_req_pri_rdy;
  assign reply = io_mem_grant_valid & T34;
  assign T34 = io_mem_grant_bits_payload_client_xact_id == 2'h1;
  assign T35 = state == 4'h5;
  assign T36 = io_mem_req_ready & io_mem_req_valid;
  assign T37 = T38 & io_meta_write_ready;
  assign T38 = state == 4'h3;
  assign T39 = T40 & reply;
  assign T40 = state == 4'h2;
  assign T41 = io_wb_req_ready & io_wb_req_valid;
  assign T42 = T59 & T43;
  assign T43 = T48 ? T47 : T44;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T46 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T47 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T33 & io_req_bits_tag_match;
  assign T60 = T59 & T61;
  assign T61 = T43 ^ 1'h1;
  assign T62 = T63 ? 4'h1 : 4'h3;
  assign T63 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T64 = T33 & T65;
  assign T65 = io_req_bits_tag_match ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = state == 4'h4;
  assign T80 = state == 4'h0;
  assign T199 = T201 & T200;
  assign T200 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T201 = wb_done | refill_done;
  assign wb_done = reply & T202;
  assign T202 = state == 4'h2;
  assign T203 = T82 ? 1'h0 : T204;
  assign T204 = T206 | T205;
  assign T205 = state == 4'h0;
  assign T206 = io_replay_ready & T207;
  assign T207 = state == 4'h8;
  assign T82 = io_meta_read_ready ^ 1'h1;
  assign T208 = T213 & T209;
  assign T209 = T210 ^ 1'h1;
  assign T210 = T212 | T211;
  assign T211 = io_req_bits_cmd == 5'h3;
  assign T212 = io_req_bits_cmd == 5'h2;
  assign T213 = T215 | T214;
  assign T214 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T150;
  assign T150 = T187 | T151;
  assign T151 = T184 & T152;
  assign T152 = T153 ^ 1'h1;
  assign T153 = T167 | T154;
  assign T154 = T156 & T155;
  assign T155 = io_mem_req_bits_a_type != 3'h1;
  assign T156 = T158 | T157;
  assign T157 = io_req_bits_cmd == 5'h6;
  assign T158 = T160 | T159;
  assign T159 = io_req_bits_cmd == 5'h3;
  assign T160 = T164 | T161;
  assign T161 = T163 | T162;
  assign T162 = io_req_bits_cmd == 5'h4;
  assign T163 = io_req_bits_cmd[2'h3:2'h3];
  assign T164 = T166 | T165;
  assign T165 = io_req_bits_cmd == 5'h7;
  assign T166 = io_req_bits_cmd == 5'h1;
  assign T167 = T177 & T168;
  assign T168 = T170 | T169;
  assign T169 = 3'h6 == io_mem_req_bits_a_type;
  assign T170 = T172 | T171;
  assign T171 = 3'h5 == io_mem_req_bits_a_type;
  assign T172 = T174 | T173;
  assign T173 = 3'h4 == io_mem_req_bits_a_type;
  assign T174 = T176 | T175;
  assign T175 = 3'h3 == io_mem_req_bits_a_type;
  assign T176 = 3'h2 == io_mem_req_bits_a_type;
  assign T177 = T181 | T178;
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h4;
  assign T180 = io_req_bits_cmd[2'h3:2'h3];
  assign T181 = T183 | T182;
  assign T182 = io_req_bits_cmd == 5'h6;
  assign T183 = io_req_bits_cmd == 5'h0;
  assign T184 = T186 | T185;
  assign T185 = state == 4'h5;
  assign T186 = state == 4'h4;
  assign T187 = T189 | T188;
  assign T188 = state == 4'h3;
  assign T189 = T191 | T190;
  assign T190 = state == 4'h2;
  assign T191 = state == 4'h1;
  assign idx_match = req_idx == T70;
  assign T70 = io_req_bits_addr[4'hc:3'h6];
  assign req_idx = req_addr[4'hc:3'h6];
  assign T71 = T33 ? io_req_bits_addr : req_addr;
  assign T215 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T0;
  assign T0 = T69 | T1;
  assign T1 = T8 & T2;
  assign T2 = meta_hazard == 2'h0;
  assign T193 = reset ? 2'h0 : T3;
  assign T3 = T7 ? 2'h1 : T4;
  assign T4 = T6 ? T5 : meta_hazard;
  assign T5 = meta_hazard + 2'h1;
  assign T6 = meta_hazard != 2'h0;
  assign T7 = io_meta_write_ready & io_meta_write_valid;
  assign T8 = T66 & T9;
  assign T9 = state != 4'h3;
  assign T66 = T68 & T67;
  assign T67 = state != 4'h2;
  assign T68 = state != 4'h1;
  assign T69 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T72 = T33 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T73 = T33 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T74;
  assign T74 = T75 & ackq_io_enq_ready;
  assign T75 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T76;
  assign T76 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T81;
  assign T81 = T82 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T195;
  assign T195 = {12'h0, T83};
  assign T83 = T84;
  assign T84 = {io_tag, T85};
  assign T85 = {req_idx, T86};
  assign T86 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T87;
  assign T87 = T88 & rpq_io_deq_valid;
  assign T88 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T89;
  assign T89 = T107 ? meta_on_flush_state : line_state_state;
  assign T90 = T42 ? meta_on_hit_state : T91;
  assign T91 = T33 ? meta_on_flush_state : T92;
  assign T92 = T32 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T93;
  assign T93 = T98 ? 2'h1 : T94;
  assign T94 = T97 ? 2'h2 : T95;
  assign T95 = T96 ? 2'h2 : 2'h0;
  assign T96 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T97 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T98 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_hit_state = T99;
  assign T99 = T100 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T107 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T108;
  assign T108 = T110 | T109;
  assign T109 = state == 4'h3;
  assign T110 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T111;
  assign T111 = state == 4'h8;
  assign io_mem_resp_data = T196;
  assign T196 = {64'h0, req_data};
  assign T112 = T33 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T113;
  assign T113 = T114 << 3'h4;
  assign T114 = {req_idx, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T115 = T33 ? T130 : T116;
  assign T116 = T129 ? T117 : acquire_type;
  assign T117 = T118 ? 3'h1 : io_mem_req_bits_a_type;
  assign T118 = T120 | T119;
  assign T119 = io_req_bits_cmd == 5'h6;
  assign T120 = T122 | T121;
  assign T121 = io_req_bits_cmd == 5'h3;
  assign T122 = T126 | T123;
  assign T123 = T125 | T124;
  assign T124 = io_req_bits_cmd == 5'h4;
  assign T125 = io_req_bits_cmd[2'h3:2'h3];
  assign T126 = T128 | T127;
  assign T127 = io_req_bits_cmd == 5'h7;
  assign T128 = io_req_bits_cmd == 5'h1;
  assign T129 = io_req_sec_val & io_req_sec_rdy;
  assign T130 = T131 ? 3'h1 : 3'h0;
  assign T131 = T133 | T132;
  assign T132 = io_req_bits_cmd == 5'h6;
  assign T133 = T135 | T134;
  assign T134 = io_req_bits_cmd == 5'h3;
  assign T135 = T139 | T136;
  assign T136 = T138 | T137;
  assign T137 = io_req_bits_cmd == 5'h4;
  assign T138 = io_req_bits_cmd[2'h3:2'h3];
  assign T139 = T141 | T140;
  assign T140 = io_req_bits_cmd == 5'h7;
  assign T141 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 2'h1;
  assign io_mem_req_bits_addr = T142;
  assign T142 = T143;
  assign T143 = {io_tag, req_idx};
  assign io_mem_req_valid = T144;
  assign T144 = T145 & ackq_io_enq_ready;
  assign T145 = state == 4'h4;
  assign io_tag = T197;
  assign T197 = T146[5'h12:1'h0];
  assign T146 = req_addr >> 4'hd;
  assign io_idx_match = T147;
  assign T147 = T148 & idx_match;
  assign T148 = state != 4'h0;
  assign io_req_sec_rdy = T149;
  assign T149 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T192;
  assign T192 = state == 4'h0;
  Queue_12 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T208 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T203 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_9 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T199 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T198 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T64) begin
      state <= T62;
    end else if(T60) begin
      state <= 4'h4;
    end else if(T42) begin
      state <= 4'h6;
    end else if(T41) begin
      state <= 4'h2;
    end else if(T39) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= 4'h5;
    end else if(T27) begin
      state <= 4'h6;
    end else if(T25) begin
      state <= 4'h7;
    end else if(T24) begin
      state <= 4'h8;
    end else if(T21) begin
      state <= 4'h0;
    end
    if(T33) begin
      refill_count <= 2'h0;
    end else if(T32) begin
      refill_count <= T31;
    end
    if(T33) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T7) begin
      meta_hazard <= 2'h1;
    end else if(T6) begin
      meta_hazard <= T5;
    end
    if(T33) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T33) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T42) begin
      line_state_state <= meta_on_hit_state;
    end else if(T33) begin
      line_state_state <= meta_on_flush_state;
    end else if(T32) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T33) begin
      req_data <= io_req_bits_data;
    end
    if(T33) begin
      acquire_type <= T130;
    end else if(T129) begin
      acquire_type <= T117;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output[2:0] io_mem_req_bits_a_type,
    output[5:0] io_mem_req_bits_write_mask,
    output[2:0] io_mem_req_bits_subword_addr,
    output[3:0] io_mem_req_bits_atomic_opcode,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire[4:0] T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire[4:0] T95;
  wire[4:0] T96;
  wire[4:0] T97;
  wire[4:0] T98;
  wire[4:0] T99;
  wire[4:0] T100;
  wire[4:0] T101;
  wire[4:0] T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire[4:0] T106;
  wire[4:0] T107;
  wire T108;
  wire[16:0] T21;
  wire[16:0] T22;
  reg [16:0] sdq_val;
  wire[16:0] T109;
  wire[31:0] T110;
  wire[31:0] T23;
  wire[31:0] T111;
  wire[31:0] T24;
  wire[31:0] T112;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T113;
  wire sdq_enq;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire[16:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire[16:0] T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire[16:0] T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire[16:0] T41;
  wire[16:0] T42;
  wire[16:0] T43;
  wire T44;
  wire[16:0] T45;
  wire[16:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[31:0] T114;
  wire[16:0] T66;
  wire[16:0] T115;
  wire free_sdq;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[31:0] T75;
  wire[31:0] T116;
  wire T76;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T134;
  wire tag_match;
  wire[30:0] T88;
  wire[30:0] T133;
  wire[18:0] T89;
  wire[18:0] T90;
  wire[18:0] tagList_1;
  wire idxMatch_1;
  wire[18:0] T91;
  wire[18:0] tagList_0;
  wire idxMatch_0;
  wire T135;
  wire sdq_rdy;
  wire T85;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire idx_match;
  wire T140;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[63:0] T8;
  reg [63:0] sdq [16:0];
  wire[63:0] T9;
  wire T10;
  wire T11;
  wire[4:0] T12;
  reg [4:0] R77;
  wire[4:0] T78;
  wire[127:0] T79;
  wire[127:0] memRespMux_0_data;
  wire[127:0] memRespMux_1_data;
  wire T80;
  wire T132;
  wire[1:0] T81;
  wire[1:0] memRespMux_0_wmask;
  wire[1:0] memRespMux_1_wmask;
  wire[12:0] T82;
  wire[12:0] memRespMux_0_addr;
  wire[12:0] memRespMux_1_addr;
  wire[3:0] T83;
  wire[3:0] memRespMux_0_way_en;
  wire[3:0] memRespMux_1_way_en;
  wire T84;
  wire T86;
  wire pri_rdy;
  wire T87;
  wire sec_rdy;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[6:0] meta_read_arb_io_out_bits_idx;
  wire[18:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[6:0] meta_write_arb_io_out_bits_idx;
  wire[3:0] meta_write_arb_io_out_bits_way_en;
  wire[18:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr;
  wire[1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[511:0] mem_req_arb_io_out_bits_data;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[5:0] mem_req_arb_io_out_bits_write_mask;
  wire[2:0] mem_req_arb_io_out_bits_subword_addr;
  wire[3:0] mem_req_arb_io_out_bits_atomic_opcode;
  wire mem_finish_arb_io_in_1_ready;
  wire mem_finish_arb_io_in_0_ready;
  wire mem_finish_arb_io_out_valid;
  wire[1:0] mem_finish_arb_io_out_bits_header_src;
  wire[1:0] mem_finish_arb_io_out_bits_header_dst;
  wire[2:0] mem_finish_arb_io_out_bits_payload_master_xact_id;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[18:0] wb_req_arb_io_out_bits_tag;
  wire[6:0] wb_req_arb_io_out_bits_idx;
  wire[3:0] wb_req_arb_io_out_bits_way_en;
  wire[1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_master_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire replay_arb_io_out_bits_kill;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_phys;
  wire[43:0] replay_arb_io_out_bits_addr;
  wire[7:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire MSHR_0_io_req_pri_rdy;
  wire MSHR_0_io_req_sec_rdy;
  wire MSHR_0_io_idx_match;
  wire[18:0] MSHR_0_io_tag;
  wire MSHR_0_io_mem_req_valid;
  wire[25:0] MSHR_0_io_mem_req_bits_addr;
  wire[1:0] MSHR_0_io_mem_req_bits_client_xact_id;
  wire[2:0] MSHR_0_io_mem_req_bits_a_type;
  wire[3:0] MSHR_0_io_mem_resp_way_en;
  wire[12:0] MSHR_0_io_mem_resp_addr;
  wire[1:0] MSHR_0_io_mem_resp_wmask;
  wire[127:0] MSHR_0_io_mem_resp_data;
  wire MSHR_0_io_meta_read_valid;
  wire[6:0] MSHR_0_io_meta_read_bits_idx;
  wire[18:0] MSHR_0_io_meta_read_bits_tag;
  wire MSHR_0_io_meta_write_valid;
  wire[6:0] MSHR_0_io_meta_write_bits_idx;
  wire[3:0] MSHR_0_io_meta_write_bits_way_en;
  wire[18:0] MSHR_0_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_0_io_meta_write_bits_data_coh_state;
  wire MSHR_0_io_replay_valid;
  wire MSHR_0_io_replay_bits_kill;
  wire[2:0] MSHR_0_io_replay_bits_typ;
  wire MSHR_0_io_replay_bits_phys;
  wire[43:0] MSHR_0_io_replay_bits_addr;
  wire[63:0] MSHR_0_io_replay_bits_data;
  wire[7:0] MSHR_0_io_replay_bits_tag;
  wire[4:0] MSHR_0_io_replay_bits_cmd;
  wire[4:0] MSHR_0_io_replay_bits_sdq_id;
  wire MSHR_0_io_mem_finish_valid;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_dst;
  wire[2:0] MSHR_0_io_mem_finish_bits_payload_master_xact_id;
  wire MSHR_0_io_wb_req_valid;
  wire[18:0] MSHR_0_io_wb_req_bits_tag;
  wire[6:0] MSHR_0_io_wb_req_bits_idx;
  wire[3:0] MSHR_0_io_wb_req_bits_way_en;
  wire[1:0] MSHR_0_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_0_io_wb_req_bits_master_xact_id;
  wire[2:0] MSHR_0_io_wb_req_bits_r_type;
  wire MSHR_0_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[18:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr;
  wire[1:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[3:0] MSHR_1_io_mem_resp_way_en;
  wire[12:0] MSHR_1_io_mem_resp_addr;
  wire[1:0] MSHR_1_io_mem_resp_wmask;
  wire[127:0] MSHR_1_io_mem_resp_data;
  wire MSHR_1_io_meta_read_valid;
  wire[6:0] MSHR_1_io_meta_read_bits_idx;
  wire[18:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[6:0] MSHR_1_io_meta_write_bits_idx;
  wire[3:0] MSHR_1_io_meta_write_bits_way_en;
  wire[18:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire MSHR_1_io_replay_bits_kill;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_phys;
  wire[43:0] MSHR_1_io_replay_bits_addr;
  wire[63:0] MSHR_1_io_replay_bits_data;
  wire[7:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_mem_finish_valid;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_dst;
  wire[2:0] MSHR_1_io_mem_finish_bits_payload_master_xact_id;
  wire MSHR_1_io_wb_req_valid;
  wire[18:0] MSHR_1_io_wb_req_bits_tag;
  wire[6:0] MSHR_1_io_wb_req_bits_idx;
  wire[3:0] MSHR_1_io_wb_req_bits_way_en;
  wire[1:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_master_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R77 = {1{$random}};
  end
`endif

  assign T92 = T131 ? 1'h0 : T93;
  assign T93 = T130 ? 1'h1 : T94;
  assign T94 = T129 ? 2'h2 : T95;
  assign T95 = T128 ? 2'h3 : T96;
  assign T96 = T127 ? 3'h4 : T97;
  assign T97 = T126 ? 3'h5 : T98;
  assign T98 = T125 ? 3'h6 : T99;
  assign T99 = T124 ? 3'h7 : T100;
  assign T100 = T123 ? 4'h8 : T101;
  assign T101 = T122 ? 4'h9 : T102;
  assign T102 = T121 ? 4'ha : T103;
  assign T103 = T120 ? 4'hb : T104;
  assign T104 = T119 ? 4'hc : T105;
  assign T105 = T118 ? 4'hd : T106;
  assign T106 = T117 ? 4'he : T107;
  assign T107 = T108 ? 4'hf : 5'h10;
  assign T108 = T21[4'hf:4'hf];
  assign T21 = ~ T22;
  assign T22 = sdq_val[5'h10:1'h0];
  assign T109 = T110[5'h10:1'h0];
  assign T110 = reset ? 32'h0 : T23;
  assign T23 = T76 ? T24 : T111;
  assign T111 = {15'h0, sdq_val};
  assign T24 = T63 | T112;
  assign T112 = {15'h0, T25};
  assign T25 = T27 & T26;
  assign T26 = 17'h0 - T113;
  assign T113 = {16'h0, sdq_enq};
  assign sdq_enq = T20 & T13;
  assign T13 = T17 | T14;
  assign T14 = T16 | T15;
  assign T15 = io_req_bits_cmd == 5'h4;
  assign T16 = io_req_bits_cmd[2'h3:2'h3];
  assign T17 = T19 | T18;
  assign T18 = io_req_bits_cmd == 5'h7;
  assign T19 = io_req_bits_cmd == 5'h1;
  assign T20 = io_req_valid & io_req_ready;
  assign T27 = T62 ? 17'h1 : T28;
  assign T28 = T61 ? 17'h2 : T29;
  assign T29 = T60 ? 17'h4 : T30;
  assign T30 = T59 ? 17'h8 : T31;
  assign T31 = T58 ? 17'h10 : T32;
  assign T32 = T57 ? 17'h20 : T33;
  assign T33 = T56 ? 17'h40 : T34;
  assign T34 = T55 ? 17'h80 : T35;
  assign T35 = T54 ? 17'h100 : T36;
  assign T36 = T53 ? 17'h200 : T37;
  assign T37 = T52 ? 17'h400 : T38;
  assign T38 = T51 ? 17'h800 : T39;
  assign T39 = T50 ? 17'h1000 : T40;
  assign T40 = T49 ? 17'h2000 : T41;
  assign T41 = T48 ? 17'h4000 : T42;
  assign T42 = T47 ? 17'h8000 : T43;
  assign T43 = T44 ? 17'h10000 : 17'h0;
  assign T44 = T45[5'h10:5'h10];
  assign T45 = ~ T46;
  assign T46 = sdq_val[5'h10:1'h0];
  assign T47 = T45[4'hf:4'hf];
  assign T48 = T45[4'he:4'he];
  assign T49 = T45[4'hd:4'hd];
  assign T50 = T45[4'hc:4'hc];
  assign T51 = T45[4'hb:4'hb];
  assign T52 = T45[4'ha:4'ha];
  assign T53 = T45[4'h9:4'h9];
  assign T54 = T45[4'h8:4'h8];
  assign T55 = T45[3'h7:3'h7];
  assign T56 = T45[3'h6:3'h6];
  assign T57 = T45[3'h5:3'h5];
  assign T58 = T45[3'h4:3'h4];
  assign T59 = T45[2'h3:2'h3];
  assign T60 = T45[2'h2:2'h2];
  assign T61 = T45[1'h1:1'h1];
  assign T62 = T45[1'h0:1'h0];
  assign T63 = T116 & T64;
  assign T64 = ~ T65;
  assign T65 = T75 & T114;
  assign T114 = {15'h0, T66};
  assign T66 = 17'h0 - T115;
  assign T115 = {16'h0, free_sdq};
  assign free_sdq = T74 & T67;
  assign T67 = T71 | T68;
  assign T68 = T70 | T69;
  assign T69 = io_replay_bits_cmd == 5'h4;
  assign T70 = io_replay_bits_cmd[2'h3:2'h3];
  assign T71 = T73 | T72;
  assign T72 = io_replay_bits_cmd == 5'h7;
  assign T73 = io_replay_bits_cmd == 5'h1;
  assign T74 = io_replay_ready & io_replay_valid;
  assign T75 = 1'h1 << io_replay_bits_sdq_id;
  assign T116 = {15'h0, sdq_val};
  assign T76 = io_replay_valid | sdq_enq;
  assign T117 = T21[4'he:4'he];
  assign T118 = T21[4'hd:4'hd];
  assign T119 = T21[4'hc:4'hc];
  assign T120 = T21[4'hb:4'hb];
  assign T121 = T21[4'ha:4'ha];
  assign T122 = T21[4'h9:4'h9];
  assign T123 = T21[4'h8:4'h8];
  assign T124 = T21[3'h7:3'h7];
  assign T125 = T21[3'h6:3'h6];
  assign T126 = T21[3'h5:3'h5];
  assign T127 = T21[3'h4:3'h4];
  assign T128 = T21[2'h3:2'h3];
  assign T129 = T21[2'h2:2'h2];
  assign T130 = T21[1'h1:1'h1];
  assign T131 = T21[1'h0:1'h0];
  assign T134 = T135 & tag_match;
  assign tag_match = T133 == T88;
  assign T88 = io_req_bits_addr >> 4'hd;
  assign T133 = {12'h0, T89};
  assign T89 = T91 | T90;
  assign T90 = idxMatch_1 ? tagList_1 : 19'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T91 = idxMatch_0 ? tagList_0 : 19'h0;
  assign tagList_0 = MSHR_0_io_tag;
  assign idxMatch_0 = MSHR_0_io_idx_match;
  assign T135 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T85 ^ 1'h1;
  assign T85 = sdq_val == 17'h1ffff;
  assign T136 = T137 & tag_match;
  assign T137 = io_req_valid & sdq_rdy;
  assign T138 = T140 & T139;
  assign T139 = idx_match ^ 1'h1;
  assign idx_match = MSHR_0_io_idx_match | MSHR_1_io_idx_match;
  assign T140 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T0;
  assign T0 = T3 ? 1'h0 : T1;
  assign T1 = T2 == 1'h0;
  assign T2 = MSHR_0_io_req_pri_rdy ^ 1'h1;
  assign T3 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T4;
  assign T4 = T7 ? 1'h0 : T5;
  assign T5 = T6 == 1'h0;
  assign T6 = MSHR_0_io_probe_rdy ^ 1'h1;
  assign T7 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_master_xact_id = wb_req_arb_io_out_bits_master_xact_id;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_idx = wb_req_arb_io_out_bits_idx;
  assign io_wb_req_bits_tag = wb_req_arb_io_out_bits_tag;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_mem_finish_bits_payload_master_xact_id = mem_finish_arb_io_out_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mem_finish_arb_io_out_bits_header_dst;
  assign io_mem_finish_bits_header_src = mem_finish_arb_io_out_bits_header_src;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_replay_bits_sdq_id = replay_arb_io_out_bits_sdq_id;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_data = T8;
  assign T8 = sdq[R77];
  assign T10 = sdq_enq & T11;
  assign T11 = T12 < 5'h11;
  assign T12 = T92[3'h4:1'h0];
  assign T78 = free_sdq ? replay_arb_io_out_bits_sdq_id : R77;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_mem_resp_data = T79;
  assign T79 = T80 ? memRespMux_1_data : memRespMux_0_data;
  assign memRespMux_0_data = MSHR_0_io_mem_resp_data;
  assign memRespMux_1_data = MSHR_1_io_mem_resp_data;
  assign T80 = T132;
  assign T132 = io_mem_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_mem_resp_wmask = T81;
  assign T81 = T80 ? memRespMux_1_wmask : memRespMux_0_wmask;
  assign memRespMux_0_wmask = MSHR_0_io_mem_resp_wmask;
  assign memRespMux_1_wmask = MSHR_1_io_mem_resp_wmask;
  assign io_mem_resp_addr = T82;
  assign T82 = T80 ? memRespMux_1_addr : memRespMux_0_addr;
  assign memRespMux_0_addr = MSHR_0_io_mem_resp_addr;
  assign memRespMux_1_addr = MSHR_1_io_mem_resp_addr;
  assign io_mem_resp_way_en = T83;
  assign T83 = T80 ? memRespMux_1_way_en : memRespMux_0_way_en;
  assign memRespMux_0_way_en = MSHR_0_io_mem_resp_way_en;
  assign memRespMux_1_way_en = MSHR_1_io_mem_resp_way_en;
  assign io_mem_req_bits_atomic_opcode = mem_req_arb_io_out_bits_atomic_opcode;
  assign io_mem_req_bits_subword_addr = mem_req_arb_io_out_bits_subword_addr;
  assign io_mem_req_bits_write_mask = mem_req_arb_io_out_bits_write_mask;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr = mem_req_arb_io_out_bits_addr;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T84;
  assign T84 = T86 & sdq_rdy;
  assign T86 = idx_match ? T87 : pri_rdy;
  assign pri_rdy = MSHR_0_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T87 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_0_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_6 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  Arbiter_7 mem_req_arb(
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_in_1_bits_data(  )
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_in_1_bits_write_mask(  )
       //.io_in_1_bits_subword_addr(  )
       //.io_in_1_bits_atomic_opcode(  )
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_req_valid ),
       .io_in_0_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_in_0_bits_data(  )
       .io_in_0_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_in_0_bits_write_mask(  )
       //.io_in_0_bits_subword_addr(  )
       //.io_in_0_bits_atomic_opcode(  )
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr( mem_req_arb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_write_mask( mem_req_arb_io_out_bits_write_mask ),
       .io_out_bits_subword_addr( mem_req_arb_io_out_bits_subword_addr ),
       .io_out_bits_atomic_opcode( mem_req_arb_io_out_bits_atomic_opcode )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign mem_req_arb.io_in_1_bits_data = {16{$random}};
    assign mem_req_arb.io_in_1_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_1_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_1_bits_atomic_opcode = {1{$random}};
    assign mem_req_arb.io_in_0_bits_data = {16{$random}};
    assign mem_req_arb.io_in_0_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_0_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_0_bits_atomic_opcode = {1{$random}};
  `endif
  Arbiter_8 mem_finish_arb(
       .io_in_1_ready( mem_finish_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_finish_valid ),
       .io_in_1_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_in_1_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( mem_finish_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_finish_valid ),
       .io_in_0_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_in_0_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_mem_finish_ready ),
       .io_out_valid( mem_finish_arb_io_out_valid ),
       .io_out_bits_header_src( mem_finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( mem_finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( mem_finish_arb_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  Arbiter_5 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_wb_req_valid ),
       .io_in_0_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_tag( wb_req_arb_io_out_bits_tag ),
       .io_out_bits_idx( wb_req_arb_io_out_bits_idx ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wb_req_arb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  Arbiter_9 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_data( MSHR_1_io_replay_bits_data ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_replay_valid ),
       .io_in_0_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_in_0_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_in_0_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_in_0_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_in_0_bits_data( MSHR_0_io_replay_bits_data ),
       .io_in_0_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_in_0_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       //.io_out_bits_data(  )
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_10 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T138 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  MSHR_0 MSHR_0(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_0_io_req_pri_rdy ),
       .io_req_sec_val( T136 ),
       .io_req_sec_rdy( MSHR_0_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T92 ),
       .io_idx_match( MSHR_0_io_idx_match ),
       .io_tag( MSHR_0_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_0_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_0_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_0_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_0_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_0_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_0_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_0_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_0_io_replay_valid ),
       .io_replay_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_0_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_0_ready ),
       .io_mem_finish_valid( MSHR_0_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_0_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_0_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_0.io_mem_resp_wmask = {1{$random}};
  `endif
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T134 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T92 ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_1_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_1_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_1_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_1_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_1_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_1_ready ),
       .io_mem_finish_valid( MSHR_1_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_1.io_mem_resp_wmask = {1{$random}};
  `endif

  always @(posedge clk) begin
    sdq_val <= T109;
    if (T10)
      sdq[T92] <= io_req_bits_data;
    if(free_sdq) begin
      R77 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [6:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [6:0] io_write_bits_idx,
    input [3:0] io_write_bits_way_en,
    input [18:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[18:0] io_resp_3_tag,
    output[1:0] io_resp_3_coh_state,
    output[18:0] io_resp_2_tag,
    output[1:0] io_resp_2_coh_state,
    output[18:0] io_resp_1_tag,
    output[1:0] io_resp_1_coh_state,
    output[18:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[20:0] T1;
  wire[83:0] tags;
  wire[83:0] T2;
  wire[83:0] T3;
  wire[83:0] T4;
  wire[41:0] T5;
  wire[20:0] T6;
  wire[20:0] T40;
  wire T7;
  wire[3:0] wmask;
  wire rst;
  reg [7:0] rst_cnt;
  wire[7:0] T41;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[20:0] T10;
  wire[20:0] T42;
  wire T11;
  wire[41:0] T12;
  wire[20:0] T13;
  wire[20:0] T43;
  wire T14;
  wire[20:0] T15;
  wire[20:0] T44;
  wire T16;
  wire[83:0] T17;
  wire[41:0] T18;
  wire[20:0] wdata;
  wire[20:0] T19;
  wire[1:0] T20;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T21;
  wire[18:0] T22;
  wire[18:0] rstVal_tag;
  wire T23;
  wire[6:0] T45;
  wire[7:0] waddr;
  wire[7:0] T46;
  reg [6:0] R24;
  wire[6:0] T25;
  wire[18:0] T26;
  wire[1:0] T27;
  wire[20:0] T28;
  wire[18:0] T29;
  wire[1:0] T30;
  wire[20:0] T31;
  wire[18:0] T32;
  wire[1:0] T33;
  wire[20:0] T34;
  wire[18:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R24 = {1{$random}};
  end
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = tags[5'h14:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T45),
    .W0E(T23),
    .W0I(T17),
    .W0M(T3),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(tags)
  );
  assign T3 = T4;
  assign T4 = {T12, T5};
  assign T5 = {T10, T6};
  assign T6 = 21'h0 - T40;
  assign T40 = {20'h0, T7};
  assign T7 = wmask[1'h0:1'h0];
  assign wmask = rst ? 4'hf : io_write_bits_way_en;
  assign rst = rst_cnt < 8'h80;
  assign T41 = reset ? 8'h0 : T8;
  assign T8 = rst ? T9 : rst_cnt;
  assign T9 = rst_cnt + 8'h1;
  assign T10 = 21'h0 - T42;
  assign T42 = {20'h0, T11};
  assign T11 = wmask[1'h1:1'h1];
  assign T12 = {T15, T13};
  assign T13 = 21'h0 - T43;
  assign T43 = {20'h0, T14};
  assign T14 = wmask[2'h2:2'h2];
  assign T15 = 21'h0 - T44;
  assign T44 = {20'h0, T16};
  assign T16 = wmask[2'h3:2'h3];
  assign T17 = {T18, T18};
  assign T18 = {wdata, wdata};
  assign wdata = T19;
  assign T19 = {T22, T20};
  assign T20 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T21;
  assign T21 = 2'h0;
  assign T22 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 19'h0;
  assign T23 = rst | io_write_valid;
  assign T45 = waddr[3'h6:1'h0];
  assign waddr = rst ? rst_cnt : T46;
  assign T46 = {1'h0, io_write_bits_idx};
  assign T25 = io_read_valid ? io_read_bits_idx : R24;
  assign io_resp_0_tag = T26;
  assign T26 = T1[5'h14:2'h2];
  assign io_resp_1_coh_state = T27;
  assign T27 = T28[1'h1:1'h0];
  assign T28 = tags[6'h29:5'h15];
  assign io_resp_1_tag = T29;
  assign T29 = T28[5'h14:2'h2];
  assign io_resp_2_coh_state = T30;
  assign T30 = T31[1'h1:1'h0];
  assign T31 = tags[6'h3e:6'h2a];
  assign io_resp_2_tag = T32;
  assign T32 = T31[5'h14:2'h2];
  assign io_resp_3_coh_state = T33;
  assign T33 = T34[1'h1:1'h0];
  assign T34 = tags[7'h53:6'h3f];
  assign io_resp_3_tag = T35;
  assign T35 = T34[5'h14:2'h2];
  assign io_write_ready = T36;
  assign T36 = rst ^ 1'h1;
  assign io_read_ready = T37;
  assign T37 = T39 & T38;
  assign T38 = io_write_valid ^ 1'h1;
  assign T39 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 8'h0;
    end else if(rst) begin
      rst_cnt <= T9;
    end
    if(io_read_valid) begin
      R24 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [6:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [6:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [6:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[6:0] T5;
  wire[6:0] T6;
  wire[6:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T5;
  assign T5 = T13 ? io_in_4_bits_idx : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_valid = T14;
  assign T14 = T21 ? io_in_4_valid : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26 ^ 1'h1;
  assign T26 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T30 | io_in_2_valid;
  assign T30 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T34 | io_in_3_valid;
  assign T34 = T35 | io_in_2_valid;
  assign T35 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input [3:0] io_read_bits_way_en,
    input [12:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input [3:0] io_write_bits_way_en,
    input [12:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_3,
    output[127:0] io_resp_2,
    output[127:0] io_resp_1,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[127:0] T4;
  wire[127:0] T5;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire[8:0] raddr;
  wire[127:0] T7;
  wire[127:0] T8;
  wire[127:0] T9;
  wire[63:0] T10;
  wire[63:0] T116;
  wire T11;
  wire[1:0] T12;
  wire[63:0] T13;
  wire[63:0] T117;
  wire T14;
  wire[127:0] T15;
  wire[63:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[8:0] waddr;
  reg [8:0] R21;
  wire[8:0] T22;
  wire T26;
  wire T27;
  reg [12:0] R28;
  wire[12:0] T29;
  wire[63:0] T30;
  wire[127:0] T31;
  wire[127:0] T32;
  wire T49;
  wire T50;
  wire[127:0] T34;
  wire[127:0] T35;
  wire[127:0] T36;
  wire[63:0] T37;
  wire[63:0] T118;
  wire T38;
  wire[63:0] T39;
  wire[63:0] T119;
  wire T40;
  wire[127:0] T41;
  wire[63:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg [8:0] R47;
  wire[8:0] T48;
  wire[127:0] T51;
  wire[127:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire T55;
  wire T56;
  wire[63:0] T57;
  wire[127:0] T58;
  wire[127:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[127:0] T62;
  wire[127:0] T63;
  wire T81;
  wire T82;
  wire[1:0] T83;
  wire[127:0] T65;
  wire[127:0] T66;
  wire[127:0] T67;
  wire[63:0] T68;
  wire[63:0] T120;
  wire T69;
  wire[1:0] T70;
  wire[63:0] T71;
  wire[63:0] T121;
  wire T72;
  wire[127:0] T73;
  wire[63:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [8:0] R79;
  wire[8:0] T80;
  wire T84;
  wire T85;
  reg [12:0] R86;
  wire[12:0] T87;
  wire[63:0] T88;
  wire[127:0] T89;
  wire[127:0] T90;
  wire T107;
  wire T108;
  wire[127:0] T92;
  wire[127:0] T93;
  wire[127:0] T94;
  wire[63:0] T95;
  wire[63:0] T122;
  wire T96;
  wire[63:0] T97;
  wire[63:0] T123;
  wire T98;
  wire[127:0] T99;
  wire[63:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg [8:0] R105;
  wire[8:0] T106;
  wire[127:0] T109;
  wire[127:0] T110;
  wire[63:0] T111;
  wire[63:0] T112;
  wire T113;
  wire T114;
  wire[63:0] T115;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R21 = {1{$random}};
    R28 = {1{$random}};
    R47 = {1{$random}};
    R79 = {1{$random}};
    R86 = {1{$random}};
    R105 = {1{$random}};
  end
`endif

  assign io_resp_0 = T0;
  assign T0 = T1;
  assign T1 = {T30, T2};
  assign T2 = T26 ? T30 : T3;
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = T5;
  assign T23 = T24 & io_read_valid;
  assign T24 = T25 != 2'h0;
  assign T25 = io_read_bits_way_en[1'h1:1'h0];
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T6 T6 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T17),
    .W0I(T15),
    .W0M(T8),
    .R1A(raddr),
    .R1E(T23),
    .R1O(T5)
  );
  assign T8 = T9;
  assign T9 = {T13, T10};
  assign T10 = 64'h0 - T116;
  assign T116 = {63'h0, T11};
  assign T11 = T12[1'h0:1'h0];
  assign T12 = io_write_bits_way_en[1'h1:1'h0];
  assign T13 = 64'h0 - T117;
  assign T117 = {63'h0, T14};
  assign T14 = T12[1'h1:1'h1];
  assign T15 = {T16, T16};
  assign T16 = io_write_bits_data[6'h3f:1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_write_bits_wmask[1'h0:1'h0];
  assign T19 = T20 & io_write_valid;
  assign T20 = T12 != 2'h0;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T22 = T23 ? raddr : R21;
  assign T26 = T27;
  assign T27 = R28[2'h3:2'h3];
  assign T29 = io_read_valid ? io_read_bits_addr : R28;
  assign T30 = T31[6'h3f:1'h0];
  assign T31 = T32;
  assign T49 = T50 & io_read_valid;
  assign T50 = T25 != 2'h0;
  DataArray_T6 T33 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T43),
    .W0I(T41),
    .W0M(T35),
    .R1A(raddr),
    .R1E(T49),
    .R1O(T32)
  );
  assign T35 = T36;
  assign T36 = {T39, T37};
  assign T37 = 64'h0 - T118;
  assign T118 = {63'h0, T38};
  assign T38 = T12[1'h0:1'h0];
  assign T39 = 64'h0 - T119;
  assign T119 = {63'h0, T40};
  assign T40 = T12[1'h1:1'h1];
  assign T41 = {T42, T42};
  assign T42 = io_write_bits_data[7'h7f:7'h40];
  assign T43 = T45 & T44;
  assign T44 = io_write_bits_wmask[1'h1:1'h1];
  assign T45 = T46 & io_write_valid;
  assign T46 = T12 != 2'h0;
  assign T48 = T49 ? raddr : R47;
  assign io_resp_1 = T51;
  assign T51 = T52;
  assign T52 = {T57, T53};
  assign T53 = T55 ? T57 : T54;
  assign T54 = T4[7'h7f:7'h40];
  assign T55 = T56;
  assign T56 = R28[2'h3:2'h3];
  assign T57 = T31[7'h7f:7'h40];
  assign io_resp_2 = T58;
  assign T58 = T59;
  assign T59 = {T88, T60};
  assign T60 = T84 ? T88 : T61;
  assign T61 = T62[6'h3f:1'h0];
  assign T62 = T63;
  assign T81 = T82 & io_read_valid;
  assign T82 = T83 != 2'h0;
  assign T83 = io_read_bits_way_en[2'h3:2'h2];
  DataArray_T6 T64 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T75),
    .W0I(T73),
    .W0M(T66),
    .R1A(raddr),
    .R1E(T81),
    .R1O(T63)
  );
  assign T66 = T67;
  assign T67 = {T71, T68};
  assign T68 = 64'h0 - T120;
  assign T120 = {63'h0, T69};
  assign T69 = T70[1'h0:1'h0];
  assign T70 = io_write_bits_way_en[2'h3:2'h2];
  assign T71 = 64'h0 - T121;
  assign T121 = {63'h0, T72};
  assign T72 = T70[1'h1:1'h1];
  assign T73 = {T74, T74};
  assign T74 = io_write_bits_data[6'h3f:1'h0];
  assign T75 = T77 & T76;
  assign T76 = io_write_bits_wmask[1'h0:1'h0];
  assign T77 = T78 & io_write_valid;
  assign T78 = T70 != 2'h0;
  assign T80 = T81 ? raddr : R79;
  assign T84 = T85;
  assign T85 = R86[2'h3:2'h3];
  assign T87 = io_read_valid ? io_read_bits_addr : R86;
  assign T88 = T89[6'h3f:1'h0];
  assign T89 = T90;
  assign T107 = T108 & io_read_valid;
  assign T108 = T83 != 2'h0;
  DataArray_T6 T91 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T101),
    .W0I(T99),
    .W0M(T93),
    .R1A(raddr),
    .R1E(T107),
    .R1O(T90)
  );
  assign T93 = T94;
  assign T94 = {T97, T95};
  assign T95 = 64'h0 - T122;
  assign T122 = {63'h0, T96};
  assign T96 = T70[1'h0:1'h0];
  assign T97 = 64'h0 - T123;
  assign T123 = {63'h0, T98};
  assign T98 = T70[1'h1:1'h1];
  assign T99 = {T100, T100};
  assign T100 = io_write_bits_data[7'h7f:7'h40];
  assign T101 = T103 & T102;
  assign T102 = io_write_bits_wmask[1'h1:1'h1];
  assign T103 = T104 & io_write_valid;
  assign T104 = T70 != 2'h0;
  assign T106 = T107 ? raddr : R105;
  assign io_resp_3 = T109;
  assign T109 = T110;
  assign T110 = {T115, T111};
  assign T111 = T113 ? T115 : T112;
  assign T112 = T62[7'h7f:7'h40];
  assign T113 = T114;
  assign T114 = R86[2'h3:2'h3];
  assign T115 = T89[7'h7f:7'h40];
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T23) begin
      R21 <= raddr;
    end
    if(io_read_valid) begin
      R28 <= io_read_bits_addr;
    end
    if(T49) begin
      R47 <= raddr;
    end
    if(T81) begin
      R79 <= raddr;
    end
    if(io_read_valid) begin
      R86 <= io_read_bits_addr;
    end
    if(T107) begin
      R105 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input [3:0] io_in_3_bits_way_en,
    input [12:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [3:0] io_in_2_bits_way_en,
    input [12:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [12:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [12:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[12:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[12:0] T4;
  wire[12:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[12:0] T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[3:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : T3;
  assign T3 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = T0;
  assign T8 = T9 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign io_out_bits_way_en = T11;
  assign T11 = T16 ? T14 : T12;
  assign T12 = T13 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T13 = T7[1'h0:1'h0];
  assign T14 = T15 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T7[1'h1:1'h1];
  assign io_out_valid = T17;
  assign T17 = T22 ? T20 : T18;
  assign T18 = T19 ? io_in_1_valid : io_in_0_valid;
  assign T19 = T7[1'h0:1'h0];
  assign T20 = T21 ? io_in_3_valid : io_in_2_valid;
  assign T21 = T7[1'h0:1'h0];
  assign T22 = T7[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_2_valid;
  assign T31 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [12:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [12:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[12:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[127:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[12:0] T5;
  wire[3:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T2;
  assign T2 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T3 = T0;
  assign io_out_bits_wmask = T4;
  assign T4 = T3 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T5;
  assign T5 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [3:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T118;
  wire[87:0] T0;
  wire[87:0] T1;
  wire[87:0] T119;
  wire[87:0] T2;
  wire[87:0] wmask;
  wire[87:0] T3;
  wire[47:0] T4;
  wire[23:0] T5;
  wire[15:0] T6;
  wire[7:0] T7;
  wire[7:0] T120;
  wire T8;
  wire[10:0] T9;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[10:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[10:0] T121;
  wire[8:0] T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[10:0] T122;
  wire[7:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T123;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T124;
  wire T32;
  wire[23:0] T33;
  wire[15:0] T34;
  wire[7:0] T35;
  wire[7:0] T125;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T126;
  wire T38;
  wire[7:0] T39;
  wire[7:0] T127;
  wire T40;
  wire[39:0] T41;
  wire[23:0] T42;
  wire[15:0] T43;
  wire[7:0] T44;
  wire[7:0] T128;
  wire T45;
  wire[7:0] T46;
  wire[7:0] T129;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T130;
  wire T49;
  wire[15:0] T50;
  wire[7:0] T51;
  wire[7:0] T131;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T132;
  wire T54;
  wire[87:0] T55;
  wire[87:0] T133;
  wire[63:0] out;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] rhs;
  wire[63:0] T62;
  wire[31:0] T63;
  wire[63:0] T64;
  wire[31:0] T65;
  wire[15:0] T66;
  wire[63:0] T67;
  wire[31:0] T68;
  wire[15:0] T69;
  wire[7:0] T70;
  wire T71;
  wire max;
  wire T72;
  wire[4:0] T134;
  wire T73;
  wire[4:0] T135;
  wire min;
  wire T74;
  wire[4:0] T136;
  wire T75;
  wire[4:0] T137;
  wire less;
  wire T76;
  wire cmp_rhs;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire word;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire cmp_lhs;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire sgned;
  wire T93;
  wire[4:0] T138;
  wire T94;
  wire[4:0] T139;
  wire lt;
  wire T95;
  wire T96;
  wire lt_lo;
  wire[31:0] T97;
  wire[31:0] T98;
  wire eq_hi;
  wire[31:0] T99;
  wire[31:0] T100;
  wire lt_hi;
  wire[31:0] T101;
  wire[31:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[63:0] T106;
  wire T107;
  wire[4:0] T140;
  wire[63:0] T108;
  wire T109;
  wire[4:0] T141;
  wire[63:0] T110;
  wire T111;
  wire[4:0] T142;
  wire[63:0] adder_out;
  wire[63:0] T112;
  wire[63:0] mask;
  wire[63:0] T143;
  wire[31:0] T113;
  wire T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire T117;
  wire[4:0] T144;


  assign io_out = T118;
  assign T118 = T0[6'h3f:1'h0];
  assign T0 = T55 | T1;
  assign T1 = T2 & T119;
  assign T119 = {24'h0, io_lhs};
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T41, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = {T29, T7};
  assign T7 = 8'h0 - T120;
  assign T120 = {7'h0, T8};
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T26 ? T122 : T10;
  assign T10 = T21 ? T121 : T11;
  assign T11 = T15 ? T12 : 11'hff;
  assign T12 = 4'hf << T13;
  assign T13 = {T14, 2'h0};
  assign T14 = io_addr[2'h2:2'h2];
  assign T15 = T17 | T16;
  assign T16 = io_typ == 3'h6;
  assign T17 = io_typ == 3'h2;
  assign T121 = {2'h0, T18};
  assign T18 = 2'h3 << T19;
  assign T19 = {T20, 1'h0};
  assign T20 = io_addr[2'h2:1'h1];
  assign T21 = T23 | T22;
  assign T22 = io_typ == 3'h5;
  assign T23 = io_typ == 3'h1;
  assign T122 = {3'h0, T24};
  assign T24 = 1'h1 << T25;
  assign T25 = io_addr[2'h2:1'h0];
  assign T26 = T28 | T27;
  assign T27 = io_typ == 3'h4;
  assign T28 = io_typ == 3'h0;
  assign T29 = 8'h0 - T123;
  assign T123 = {7'h0, T30};
  assign T30 = T9[1'h1:1'h1];
  assign T31 = 8'h0 - T124;
  assign T124 = {7'h0, T32};
  assign T32 = T9[2'h2:2'h2];
  assign T33 = {T39, T34};
  assign T34 = {T37, T35};
  assign T35 = 8'h0 - T125;
  assign T125 = {7'h0, T36};
  assign T36 = T9[2'h3:2'h3];
  assign T37 = 8'h0 - T126;
  assign T126 = {7'h0, T38};
  assign T38 = T9[3'h4:3'h4];
  assign T39 = 8'h0 - T127;
  assign T127 = {7'h0, T40};
  assign T40 = T9[3'h5:3'h5];
  assign T41 = {T50, T42};
  assign T42 = {T48, T43};
  assign T43 = {T46, T44};
  assign T44 = 8'h0 - T128;
  assign T128 = {7'h0, T45};
  assign T45 = T9[3'h6:3'h6];
  assign T46 = 8'h0 - T129;
  assign T129 = {7'h0, T47};
  assign T47 = T9[3'h7:3'h7];
  assign T48 = 8'h0 - T130;
  assign T130 = {7'h0, T49};
  assign T49 = T9[4'h8:4'h8];
  assign T50 = {T53, T51};
  assign T51 = 8'h0 - T131;
  assign T131 = {7'h0, T52};
  assign T52 = T9[4'h9:4'h9];
  assign T53 = 8'h0 - T132;
  assign T132 = {7'h0, T54};
  assign T54 = T9[4'ha:4'ha];
  assign T55 = wmask & T133;
  assign T133 = {24'h0, out};
  assign out = T117 ? adder_out : T56;
  assign T56 = T111 ? T110 : T57;
  assign T57 = T109 ? T108 : T58;
  assign T58 = T107 ? T106 : T59;
  assign T59 = T71 ? io_lhs : T60;
  assign T60 = T26 ? T67 : T61;
  assign T61 = T21 ? T64 : rhs;
  assign rhs = T15 ? T62 : io_rhs;
  assign T62 = {T63, T63};
  assign T63 = io_rhs[5'h1f:1'h0];
  assign T64 = {T65, T65};
  assign T65 = {T66, T66};
  assign T66 = io_rhs[4'hf:1'h0];
  assign T67 = {T68, T68};
  assign T68 = {T69, T69};
  assign T69 = {T70, T70};
  assign T70 = io_rhs[3'h7:1'h0];
  assign T71 = less ? min : max;
  assign max = T73 | T72;
  assign T72 = T134 == 5'hf;
  assign T134 = {1'h0, io_cmd};
  assign T73 = T135 == 5'hd;
  assign T135 = {1'h0, io_cmd};
  assign min = T75 | T74;
  assign T74 = T136 == 5'he;
  assign T136 = {1'h0, io_cmd};
  assign T75 = T137 == 5'hc;
  assign T137 = {1'h0, io_cmd};
  assign less = T105 ? lt : T76;
  assign T76 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T79 ? T78 : T77;
  assign T77 = rhs[6'h3f:6'h3f];
  assign T78 = rhs[5'h1f:5'h1f];
  assign T79 = word & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_addr[2'h2:2'h2];
  assign word = T83 | T82;
  assign T82 = io_typ == 3'h4;
  assign T83 = T85 | T84;
  assign T84 = io_typ == 3'h0;
  assign T85 = T87 | T86;
  assign T86 = io_typ == 3'h6;
  assign T87 = io_typ == 3'h2;
  assign cmp_lhs = T90 ? T89 : T88;
  assign T88 = io_lhs[6'h3f:6'h3f];
  assign T89 = io_lhs[5'h1f:5'h1f];
  assign T90 = word & T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = io_addr[2'h2:2'h2];
  assign sgned = T94 | T93;
  assign T93 = T138 == 5'hd;
  assign T138 = {1'h0, io_cmd};
  assign T94 = T139 == 5'hc;
  assign T139 = {1'h0, io_cmd};
  assign lt = word ? T103 : T95;
  assign T95 = lt_hi | T96;
  assign T96 = eq_hi & lt_lo;
  assign lt_lo = T98 < T97;
  assign T97 = rhs[5'h1f:1'h0];
  assign T98 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T100 == T99;
  assign T99 = rhs[6'h3f:6'h20];
  assign T100 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T102 < T101;
  assign T101 = rhs[6'h3f:6'h20];
  assign T102 = io_lhs[6'h3f:6'h20];
  assign T103 = T104 ? lt_hi : lt_lo;
  assign T104 = io_addr[2'h2:2'h2];
  assign T105 = cmp_lhs == cmp_rhs;
  assign T106 = io_lhs ^ rhs;
  assign T107 = T140 == 5'h9;
  assign T140 = {1'h0, io_cmd};
  assign T108 = io_lhs | rhs;
  assign T109 = T141 == 5'ha;
  assign T141 = {1'h0, io_cmd};
  assign T110 = io_lhs & rhs;
  assign T111 = T142 == 5'hb;
  assign T142 = {1'h0, io_cmd};
  assign adder_out = T115 + T112;
  assign T112 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T143;
  assign T143 = {32'h0, T113};
  assign T113 = T114 << 5'h1f;
  assign T114 = io_addr[2'h2:2'h2];
  assign T115 = T116;
  assign T116 = io_lhs & mask;
  assign T117 = T144 == 5'h8;
  assign T144 = {1'h0, io_cmd};
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_master_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_master_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_master_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[511:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire[25:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_data = T4;
  assign T4 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_master_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module FlowThroughSerializer_0(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  active;
  wire T46;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T47;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T48;
  wire[1:0] T18;
  wire T19;
  wire[3:0] T20;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T49;
  wire[3:0] T21;
  wire[2:0] T22;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T50;
  wire[2:0] T23;
  wire[1:0] T24;
  reg [1:0] rbits_payload_client_xact_id;
  wire[1:0] T51;
  wire[1:0] T25;
  wire[511:0] T26;
  wire[511:0] T27;
  reg [511:0] rbits_payload_data;
  wire[511:0] T52;
  wire[511:0] T28;
  wire[511:0] T53;
  wire[127:0] T29;
  wire[127:0] T30;
  wire[127:0] shifter_0;
  wire[127:0] T31;
  wire[127:0] shifter_1;
  wire[127:0] T32;
  wire T33;
  wire[1:0] T34;
  wire[127:0] T35;
  wire[127:0] shifter_2;
  wire[127:0] T36;
  wire[127:0] shifter_3;
  wire[127:0] T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  reg [1:0] rbits_header_dst;
  wire[1:0] T54;
  wire[1:0] T41;
  wire[1:0] T42;
  reg [1:0] rbits_header_src;
  wire[1:0] T55;
  wire[1:0] T43;
  wire T44;
  wire T45;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    active = {1{$random}};
    cnt = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T14 ? 1'h1 : T1;
  assign T1 = T6 ? T2 : 1'h0;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 | T4;
  assign T4 = io_in_bits_payload_g_type == 4'h2;
  assign T5 = io_in_bits_payload_g_type == 4'h1;
  assign T6 = T7 & io_in_valid;
  assign T7 = active ^ 1'h1;
  assign T46 = reset ? 1'h0 : T8;
  assign T8 = T14 ? 1'h0 : T9;
  assign T9 = T10 ? 1'h1 : active;
  assign T10 = T6 & T11;
  assign T11 = T13 | T12;
  assign T12 = io_in_bits_payload_g_type == 4'h2;
  assign T13 = io_in_bits_payload_g_type == 4'h1;
  assign T14 = T19 & wrap;
  assign wrap = cnt == 2'h3;
  assign T47 = reset ? 2'h0 : T15;
  assign T15 = T14 ? 2'h0 : T16;
  assign T16 = T19 ? T18 : T17;
  assign T17 = T10 ? T48 : cnt;
  assign T48 = {1'h0, io_out_ready};
  assign T18 = cnt + 2'h1;
  assign T19 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T20;
  assign T20 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T49 = reset ? io_in_bits_payload_g_type : T21;
  assign T21 = T10 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T22;
  assign T22 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T50 = reset ? io_in_bits_payload_master_xact_id : T23;
  assign T23 = T10 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T24;
  assign T24 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T51 = reset ? io_in_bits_payload_client_xact_id : T25;
  assign T25 = T10 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T26;
  assign T26 = active ? T53 : T27;
  assign T27 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T52 = reset ? io_in_bits_payload_data : T28;
  assign T28 = T10 ? io_in_bits_payload_data : rbits_payload_data;
  assign T53 = {384'h0, T29};
  assign T29 = T39 ? T35 : T30;
  assign T30 = T33 ? shifter_1 : shifter_0;
  assign shifter_0 = T31;
  assign T31 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T32;
  assign T32 = rbits_payload_data[8'hff:8'h80];
  assign T33 = T34[1'h0:1'h0];
  assign T34 = cnt;
  assign T35 = T38 ? shifter_3 : shifter_2;
  assign shifter_2 = T36;
  assign T36 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T37;
  assign T37 = rbits_payload_data[9'h1ff:9'h180];
  assign T38 = T34[1'h0:1'h0];
  assign T39 = T34[1'h1:1'h1];
  assign io_out_bits_header_dst = T40;
  assign T40 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T54 = reset ? io_in_bits_header_dst : T41;
  assign T41 = T10 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T42;
  assign T42 = active ? rbits_header_src : io_in_bits_header_src;
  assign T55 = reset ? io_in_bits_header_src : T43;
  assign T43 = T10 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T44;
  assign T44 = active | io_in_valid;
  assign io_in_ready = T45;
  assign T45 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else if(T14) begin
      active <= 1'h0;
    end else if(T10) begin
      active <= 1'h1;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T14) begin
      cnt <= 2'h0;
    end else if(T19) begin
      cnt <= T18;
    end else if(T10) begin
      cnt <= T48;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T10) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T10) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T10) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T10) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T10) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T10) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input  io_cpu_req_bits_kill,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_phys,
    input [43:0] io_cpu_req_bits_addr,
    input [63:0] io_cpu_req_bits_data,
    input [7:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    output io_cpu_resp_valid,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output[2:0] io_cpu_resp_bits_typ,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[7:0] io_cpu_resp_bits_tag,
    output[3:0] io_cpu_resp_bits_cmd,
    output[43:0] io_cpu_resp_bits_addr,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[7:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    output io_cpu_ordered,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [2:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_header_src,
    output[1:0] io_mem_release_bits_header_dst,
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[2:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type
);

  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  reg [63:0] s2_req_data;
  wire[63:0] T196;
  wire[63:0] T197;
  wire[63:0] T198;
  reg  s1_replay;
  wire T424;
  wire T26;
  wire T199;
  wire s1_write;
  wire T154;
  wire T155;
  reg [4:0] s1_req_cmd;
  wire[4:0] T19;
  wire[4:0] T20;
  wire[4:0] T21;
  reg [4:0] s2_req_cmd;
  wire[4:0] T18;
  wire s2_recycle;
  wire T22;
  reg  s2_recycle_next;
  wire T423;
  wire T23;
  wire T24;
  wire T25;
  reg  s1_valid;
  wire T425;
  wire T27;
  wire T28;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire[1:0] T29;
  wire T30;
  wire s2_hit;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  reg [1:0] R45;
  wire[1:0] T46;
  wire T47;
  reg [3:0] s2_tag_match_way;
  wire[3:0] T48;
  wire[3:0] s1_tag_match_way;
  wire[3:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire[3:0] s1_tag_eq_way;
  wire[3:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[18:0] T57;
  wire[31:0] s1_addr;
  wire[12:0] T58;
  reg [43:0] s1_req_addr;
  wire[43:0] T59;
  wire[43:0] T60;
  wire[43:0] T61;
  wire[43:0] T62;
  wire[43:0] T63;
  wire[43:0] T426;
  wire[31:0] T64;
  wire[25:0] T65;
  wire[43:0] T427;
  wire[31:0] T66;
  wire[25:0] T67;
  reg [43:0] s2_req_addr;
  wire[43:0] T68;
  wire[43:0] T428;
  wire T69;
  wire[18:0] T70;
  wire[1:0] T71;
  wire T72;
  wire[18:0] T73;
  wire T74;
  wire[18:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire[1:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  reg [1:0] R89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T92;
  wire[1:0] T93;
  wire[1:0] T94;
  reg [1:0] R95;
  wire[1:0] T96;
  wire T97;
  wire[1:0] T98;
  wire[1:0] T99;
  reg [1:0] R100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire s2_tag_match;
  wire T120;
  wire s2_replay;
  wire T121;
  reg  R122;
  wire T429;
  reg  s2_valid;
  wire T430;
  wire s1_valid_masked;
  wire T123;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  wire T203;
  reg  s1_recycled;
  wire T204;
  wire[63:0] T460;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T221;
  wire[63:0] T222;
  wire[127:0] s2_data_muxed;
  wire[127:0] T223;
  wire[127:0] s2_data_3;
  wire[127:0] T224;
  wire[127:0] T225;
  reg [63:0] R226;
  wire[63:0] T433;
  wire[127:0] T227;
  wire[127:0] T434;
  wire[127:0] T228;
  wire T229;
  wire T230;
  reg [63:0] R231;
  wire[63:0] T232;
  wire[63:0] T233;
  wire T234;
  wire s1_writeback;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire[127:0] T239;
  wire[127:0] T240;
  wire[127:0] s2_data_2;
  wire[127:0] T241;
  wire[127:0] T242;
  reg [63:0] R243;
  wire[63:0] T435;
  wire[127:0] T244;
  wire[127:0] T436;
  wire[127:0] T245;
  wire T246;
  wire T247;
  reg [63:0] R248;
  wire[63:0] T249;
  wire[63:0] T250;
  wire T251;
  wire T252;
  wire[127:0] T253;
  wire[127:0] T254;
  wire[127:0] s2_data_1;
  wire[127:0] T255;
  wire[127:0] T256;
  reg [63:0] R257;
  wire[63:0] T437;
  wire[127:0] T258;
  wire[127:0] T438;
  wire[127:0] T259;
  wire T260;
  wire T261;
  reg [63:0] R262;
  wire[63:0] T263;
  wire[63:0] T264;
  wire T265;
  wire T266;
  wire[127:0] T267;
  wire[127:0] s2_data_0;
  wire[127:0] T268;
  wire[127:0] T269;
  reg [63:0] R270;
  wire[63:0] T439;
  wire[127:0] T271;
  wire[127:0] T440;
  wire[127:0] T272;
  wire T273;
  wire T274;
  reg [63:0] R275;
  wire[63:0] T276;
  wire[63:0] T277;
  wire T278;
  wire T279;
  wire[63:0] T280;
  wire[127:0] T441;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T281;
  wire[63:0] T282;
  wire[63:0] T283;
  reg [63:0] s4_req_data;
  wire[63:0] T284;
  wire T285;
  reg  s3_valid;
  wire T442;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire s2_sc_fail;
  wire T206;
  wire s2_lrsc_addr_match;
  wire T207;
  wire[37:0] T208;
  reg [37:0] lrsc_addr;
  wire[37:0] T209;
  wire[37:0] T210;
  wire T17;
  wire s2_lr;
  wire T124;
  wire T125;
  wire s2_valid_masked;
  wire T126;
  wire T127;
  wire s2_nack;
  wire s2_nack_miss;
  wire T128;
  wire T129;
  wire T130;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T131;
  wire s1_nack;
  wire T132;
  wire T133;
  wire T134;
  wire[6:0] T135;
  wire T136;
  wire T137;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T422;
  wire[4:0] T10;
  wire[4:0] T11;
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire T15;
  wire T16;
  wire T138;
  wire s2_sc;
  wire T296;
  wire T297;
  reg [63:0] s3_req_data;
  wire[63:0] T443;
  wire[127:0] T298;
  wire[127:0] T444;
  wire[63:0] T299;
  wire[127:0] T300;
  wire[127:0] T445;
  wire[127:0] s2_data_corrected;
  wire[127:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  reg [4:0] s3_req_cmd;
  wire[4:0] T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire[40:0] T323;
  reg [43:0] s3_req_addr;
  wire[43:0] T324;
  wire[40:0] T446;
  wire[28:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire[40:0] T336;
  wire[40:0] T447;
  wire[28:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  reg [4:0] s4_req_cmd;
  wire[4:0] T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[40:0] T354;
  reg [43:0] s4_req_addr;
  wire[43:0] T355;
  wire[40:0] T448;
  wire[28:0] T356;
  reg  s4_valid;
  wire T449;
  wire T357;
  reg  s2_store_bypass;
  wire T358;
  wire T359;
  reg [2:0] s2_req_typ;
  wire[2:0] T175;
  reg [2:0] s1_req_typ;
  wire[2:0] T172;
  wire[2:0] T173;
  wire[2:0] T174;
  wire[3:0] T461;
  wire[5:0] T462;
  wire[127:0] T463;
  wire[1:0] T464;
  wire T465;
  wire T466;
  wire[12:0] T467;
  reg [3:0] s3_way;
  wire[3:0] T468;
  wire[127:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[12:0] T476;
  wire[12:0] T477;
  wire[12:0] T478;
  wire[127:0] T479;
  wire[127:0] T480;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[6:0] T481;
  wire[37:0] T482;
  wire[6:0] T483;
  wire[37:0] T484;
  reg  s1_req_phys;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  reg  s2_req_phys;
  wire T490;
  wire[30:0] T491;
  wire T492;
  wire T493;
  wire T494;
  wire s1_readwrite;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire s1_read;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T499;
  wire T500;
  wire[3:0] T501;
  wire[3:0] s2_replaced_way_en;
  reg [1:0] R502;
  wire[1:0] T503;
  wire[1:0] T504;
  reg [15:0] R505;
  wire[15:0] T506;
  wire[15:0] T507;
  wire[15:0] T508;
  wire[14:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire[1:0] T519;
  wire[1:0] T520;
  wire[20:0] T521;
  wire[20:0] T522;
  wire[20:0] T523;
  wire[20:0] T524;
  reg [1:0] R525;
  wire[1:0] T526;
  wire T527;
  wire T528;
  wire[3:0] s1_replaced_way_en;
  wire[1:0] T529;
  reg [18:0] R530;
  wire[18:0] T531;
  wire T532;
  wire[20:0] T533;
  wire[20:0] T534;
  wire[20:0] T535;
  wire[20:0] T536;
  reg [1:0] R537;
  wire[1:0] T538;
  wire T539;
  wire T540;
  reg [18:0] R541;
  wire[18:0] T542;
  wire T543;
  wire[20:0] T544;
  wire[20:0] T545;
  wire[20:0] T546;
  wire[20:0] T547;
  reg [1:0] R548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  reg [18:0] R552;
  wire[18:0] T553;
  wire T554;
  wire[20:0] T555;
  wire[20:0] T556;
  wire[20:0] T557;
  reg [1:0] R558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  reg [18:0] R562;
  wire[18:0] T563;
  wire T564;
  wire[1:0] T565;
  wire[18:0] T566;
  wire[18:0] T567;
  wire[18:0] T568;
  reg [7:0] s2_req_tag;
  wire[7:0] T193;
  reg [7:0] s1_req_tag;
  wire[7:0] T190;
  wire[7:0] T191;
  wire[7:0] T192;
  reg  s2_req_kill;
  wire T569;
  reg  s1_req_kill;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] probe_bits_p_type;
  wire[2:0] probe_bits_master_xact_id;
  wire[25:0] probe_bits_addr;
  wire T596;
  wire T597;
  wire probe_valid;
  wire[2:0] T0;
  wire[511:0] T1;
  wire[2:0] T2;
  wire[1:0] T3;
  wire[25:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire probe_ready;
  wire T8;
  wire T9;
  wire[3:0] T139;
  wire[2:0] T140;
  wire[5:0] T141;
  wire[2:0] T142;
  wire[511:0] T143;
  wire[1:0] T144;
  wire[25:0] T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T160;
  wire T167;
  wire misaligned;
  wire T168;
  wire T169;
  wire[2:0] T170;
  wire T171;
  wire T176;
  wire T177;
  wire T178;
  wire[1:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T194;
  wire T195;
  wire s1_sc;
  wire[3:0] T431;
  wire[63:0] T205;
  wire[63:0] T432;
  wire[63:0] T211;
  wire[7:0] T212;
  wire[7:0] T213;
  wire[7:0] T214;
  wire[63:0] T215;
  wire[15:0] T216;
  wire[15:0] T217;
  wire[63:0] T218;
  wire[31:0] T219;
  wire[31:0] T220;
  wire[31:0] T360;
  wire T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire[31:0] T364;
  wire[31:0] T450;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire[15:0] T377;
  wire T378;
  wire[47:0] T379;
  wire[47:0] T380;
  wire[47:0] T381;
  wire[47:0] T451;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire[7:0] T387;
  wire T388;
  wire[55:0] T389;
  wire[55:0] T390;
  wire[55:0] T391;
  wire[55:0] T452;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  reg  block_miss;
  wire T453;
  wire T420;
  wire T421;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[6:0] wb_io_meta_read_bits_idx;
  wire[18:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire[3:0] wb_io_data_req_bits_way_en;
  wire[12:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[25:0] wb_io_release_bits_addr;
  wire[1:0] wb_io_release_bits_client_xact_id;
  wire[2:0] wb_io_release_bits_master_xact_id;
  wire[511:0] wb_io_release_bits_data;
  wire[2:0] wb_io_release_bits_r_type;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[25:0] prober_io_rep_bits_addr;
  wire[1:0] prober_io_rep_bits_client_xact_id;
  wire[2:0] prober_io_rep_bits_master_xact_id;
  wire[511:0] prober_io_rep_bits_data;
  wire[2:0] prober_io_rep_bits_r_type;
  wire prober_io_meta_read_valid;
  wire[6:0] prober_io_meta_read_bits_idx;
  wire[18:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[6:0] prober_io_meta_write_bits_idx;
  wire[3:0] prober_io_meta_write_bits_way_en;
  wire[18:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[18:0] prober_io_wb_req_bits_tag;
  wire[6:0] prober_io_wb_req_bits_idx;
  wire[3:0] prober_io_wb_req_bits_way_en;
  wire[1:0] prober_io_wb_req_bits_client_xact_id;
  wire[2:0] prober_io_wb_req_bits_master_xact_id;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[18:0] meta_io_resp_3_tag;
  wire[1:0] meta_io_resp_3_coh_state;
  wire[18:0] meta_io_resp_2_tag;
  wire[1:0] meta_io_resp_2_coh_state;
  wire[18:0] meta_io_resp_1_tag;
  wire[1:0] meta_io_resp_1_coh_state;
  wire[18:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[6:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[6:0] metaWriteArb_io_out_bits_idx;
  wire[3:0] metaWriteArb_io_out_bits_way_en;
  wire[18:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_3;
  wire[127:0] data_io_resp_2;
  wire[127:0] data_io_resp_1;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire[3:0] readArb_io_out_bits_way_en;
  wire[12:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire[3:0] writeArb_io_out_bits_way_en;
  wire[12:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[25:0] releaseArb_io_out_bits_addr;
  wire[1:0] releaseArb_io_out_bits_client_xact_id;
  wire[2:0] releaseArb_io_out_bits_master_xact_id;
  wire[511:0] releaseArb_io_out_bits_data;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire FlowThroughSerializer_0_io_in_ready;
  wire FlowThroughSerializer_0_io_out_valid;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_header_src;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_header_dst;
  wire[511:0] FlowThroughSerializer_0_io_out_bits_payload_data;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_payload_client_xact_id;
  wire[2:0] FlowThroughSerializer_0_io_out_bits_payload_master_xact_id;
  wire[3:0] FlowThroughSerializer_0_io_out_bits_payload_g_type;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[18:0] wbArb_io_out_bits_tag;
  wire[6:0] wbArb_io_out_bits_idx;
  wire[3:0] wbArb_io_out_bits_way_en;
  wire[1:0] wbArb_io_out_bits_client_xact_id;
  wire[2:0] wbArb_io_out_bits_master_xact_id;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[18:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[29:0] dtlb_io_ptw_req_bits;
  wire mshrs_io_req_ready;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr;
  wire[1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[511:0] mshrs_io_mem_req_bits_data;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[5:0] mshrs_io_mem_req_bits_write_mask;
  wire[2:0] mshrs_io_mem_req_bits_subword_addr;
  wire[3:0] mshrs_io_mem_req_bits_atomic_opcode;
  wire[3:0] mshrs_io_mem_resp_way_en;
  wire[12:0] mshrs_io_mem_resp_addr;
  wire mshrs_io_meta_read_valid;
  wire[6:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[6:0] mshrs_io_meta_write_bits_idx;
  wire[3:0] mshrs_io_meta_write_bits_way_en;
  wire[18:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire mshrs_io_replay_bits_kill;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_phys;
  wire[43:0] mshrs_io_replay_bits_addr;
  wire[63:0] mshrs_io_replay_bits_data;
  wire[7:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire mshrs_io_mem_finish_valid;
  wire[1:0] mshrs_io_mem_finish_bits_header_src;
  wire[1:0] mshrs_io_mem_finish_bits_header_dst;
  wire[2:0] mshrs_io_mem_finish_bits_payload_master_xact_id;
  wire mshrs_io_wb_req_valid;
  wire[18:0] mshrs_io_wb_req_bits_tag;
  wire[6:0] mshrs_io_wb_req_bits_idx;
  wire[3:0] mshrs_io_wb_req_bits_way_en;
  wire[1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_master_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    R45 = {1{$random}};
    s2_tag_match_way = {1{$random}};
    s1_req_addr = {2{$random}};
    s2_req_addr = {2{$random}};
    R89 = {1{$random}};
    R95 = {1{$random}};
    R100 = {1{$random}};
    R122 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R226 = {2{$random}};
    R231 = {2{$random}};
    R243 = {2{$random}};
    R248 = {2{$random}};
    R257 = {2{$random}};
    R262 = {2{$random}};
    R270 = {2{$random}};
    R275 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R502 = {1{$random}};
    R505 = {1{$random}};
    R525 = {1{$random}};
    R530 = {1{$random}};
    R537 = {1{$random}};
    R541 = {1{$random}};
    R548 = {1{$random}};
    R552 = {1{$random}};
    R558 = {1{$random}};
    R562 = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    block_miss = {1{$random}};
  end
`endif

  assign T454 = writeArb_io_in_1_ready | T455;
  assign T455 = T456 ^ 1'h1;
  assign T456 = T458 | T457;
  assign T457 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h2;
  assign T458 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h1;
  assign T459 = io_mem_release_ready;
  assign T196 = T203 ? s1_req_data : T197;
  assign T197 = T199 ? T198 : s2_req_data;
  assign T198 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T424 = reset ? 1'h0 : T26;
  assign T26 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T199 = s1_clk_en & s1_write;
  assign s1_write = T157 | T154;
  assign T154 = T156 | T155;
  assign T155 = s1_req_cmd == 5'h4;
  assign T19 = s2_recycle ? s2_req_cmd : T20;
  assign T20 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T21;
  assign T21 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T18 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T22;
  assign T22 = s2_recycle_ecc | s2_recycle_next;
  assign T423 = reset ? 1'h0 : T23;
  assign T23 = T28 ? T24 : s2_recycle_next;
  assign T24 = T25 & s2_recycle_ecc;
  assign T25 = s1_valid | s1_replay;
  assign T425 = reset ? 1'h0 : T27;
  assign T27 = io_cpu_req_ready & io_cpu_req_valid;
  assign T28 = s1_valid | s1_replay;
  assign s2_recycle_ecc = T30 & s2_data_correctable;
  assign s2_data_correctable = T29[1'h0:1'h0];
  assign T29 = 2'h0;
  assign T30 = T120 & s2_hit;
  assign s2_hit = T103 & T31;
  assign T31 = T41 == T32;
  assign T32 = T33;
  assign T33 = T34 ? 2'h2 : T41;
  assign T34 = T38 | T35;
  assign T35 = T37 | T36;
  assign T36 = s2_req_cmd == 5'h4;
  assign T37 = s2_req_cmd[2'h3:2'h3];
  assign T38 = T40 | T39;
  assign T39 = s2_req_cmd == 5'h7;
  assign T40 = s2_req_cmd == 5'h1;
  assign T41 = T42[1'h1:1'h0];
  assign T42 = T86 | T43;
  assign T43 = T47 ? T44 : 2'h0;
  assign T44 = R45;
  assign T46 = s1_clk_en ? meta_io_resp_3_coh_state : R45;
  assign T47 = s2_tag_match_way[2'h3:2'h3];
  assign T48 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T49;
  assign T49 = {T79, T50};
  assign T50 = {T76, T51};
  assign T51 = T53 & T52;
  assign T52 = meta_io_resp_0_coh_state != 2'h0;
  assign T53 = s1_tag_eq_way[1'h0:1'h0];
  assign s1_tag_eq_way = T54;
  assign T54 = {T71, T55};
  assign T55 = {T69, T56};
  assign T56 = meta_io_resp_0_tag == T57;
  assign T57 = s1_addr >> 4'hd;
  assign s1_addr = {dtlb_io_resp_ppn, T58};
  assign T58 = s1_req_addr[4'hc:1'h0];
  assign T59 = s2_recycle ? s2_req_addr : T60;
  assign T60 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T61;
  assign T61 = prober_io_meta_read_valid ? T427 : T62;
  assign T62 = wb_io_meta_read_valid ? T426 : T63;
  assign T63 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T426 = {12'h0, T64};
  assign T64 = T65 << 3'h6;
  assign T65 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T427 = {12'h0, T66};
  assign T66 = T67 << 3'h6;
  assign T67 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T68 = s1_clk_en ? T428 : s2_req_addr;
  assign T428 = {12'h0, s1_addr};
  assign T69 = meta_io_resp_1_tag == T70;
  assign T70 = s1_addr >> 4'hd;
  assign T71 = {T74, T72};
  assign T72 = meta_io_resp_2_tag == T73;
  assign T73 = s1_addr >> 4'hd;
  assign T74 = meta_io_resp_3_tag == T75;
  assign T75 = s1_addr >> 4'hd;
  assign T76 = T78 & T77;
  assign T77 = meta_io_resp_1_coh_state != 2'h0;
  assign T78 = s1_tag_eq_way[1'h1:1'h1];
  assign T79 = {T83, T80};
  assign T80 = T82 & T81;
  assign T81 = meta_io_resp_2_coh_state != 2'h0;
  assign T82 = s1_tag_eq_way[2'h2:2'h2];
  assign T83 = T85 & T84;
  assign T84 = meta_io_resp_3_coh_state != 2'h0;
  assign T85 = s1_tag_eq_way[2'h3:2'h3];
  assign T86 = T92 | T87;
  assign T87 = T91 ? T88 : 2'h0;
  assign T88 = R89;
  assign T90 = s1_clk_en ? meta_io_resp_2_coh_state : R89;
  assign T91 = s2_tag_match_way[2'h2:2'h2];
  assign T92 = T98 | T93;
  assign T93 = T97 ? T94 : 2'h0;
  assign T94 = R95;
  assign T96 = s1_clk_en ? meta_io_resp_1_coh_state : R95;
  assign T97 = s2_tag_match_way[1'h1:1'h1];
  assign T98 = T102 ? T99 : 2'h0;
  assign T99 = R100;
  assign T101 = s1_clk_en ? meta_io_resp_0_coh_state : R100;
  assign T102 = s2_tag_match_way[1'h0:1'h0];
  assign T103 = s2_tag_match & T104;
  assign T104 = T109 ? T108 : T105;
  assign T105 = T107 | T106;
  assign T106 = T41 == 2'h2;
  assign T107 = T41 == 2'h1;
  assign T108 = T41 == 2'h2;
  assign T109 = T111 | T110;
  assign T110 = s2_req_cmd == 5'h6;
  assign T111 = T113 | T112;
  assign T112 = s2_req_cmd == 5'h3;
  assign T113 = T117 | T114;
  assign T114 = T116 | T115;
  assign T115 = s2_req_cmd == 5'h4;
  assign T116 = s2_req_cmd[2'h3:2'h3];
  assign T117 = T119 | T118;
  assign T118 = s2_req_cmd == 5'h7;
  assign T119 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 4'h0;
  assign T120 = s2_valid | s2_replay;
  assign s2_replay = R122 & T121;
  assign T121 = s2_req_cmd != 5'h5;
  assign T429 = reset ? 1'h0 : s1_replay;
  assign T430 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T123;
  assign T123 = io_cpu_req_bits_kill ^ 1'h1;
  assign T156 = s1_req_cmd[2'h3:2'h3];
  assign T157 = T159 | T158;
  assign T158 = s1_req_cmd == 5'h7;
  assign T159 = s1_req_cmd == 5'h1;
  assign T200 = s2_recycle ? s2_req_data : T201;
  assign T201 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T202;
  assign T202 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T203 = s1_clk_en & s1_recycled;
  assign T204 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T460 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T441 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> 7'h0;
  assign s2_data_uncorrected = T221;
  assign T221 = {T280, T222};
  assign T222 = s2_data_muxed[6'h3f:1'h0];
  assign s2_data_muxed = T239 | T223;
  assign T223 = T238 ? s2_data_3 : 128'h0;
  assign s2_data_3 = T224;
  assign T224 = T225;
  assign T225 = {R231, R226};
  assign T433 = T227[6'h3f:1'h0];
  assign T227 = T229 ? T228 : T434;
  assign T434 = {64'h0, R226};
  assign T228 = data_io_resp_3 >> 1'h0;
  assign T229 = s1_clk_en & T230;
  assign T230 = s1_tag_eq_way[2'h3:2'h3];
  assign T232 = T234 ? T233 : R231;
  assign T233 = data_io_resp_3 >> 7'h40;
  assign T234 = T229 & s1_writeback;
  assign s1_writeback = T236 & T235;
  assign T235 = s1_replay ^ 1'h1;
  assign T236 = s1_clk_en & T237;
  assign T237 = s1_valid ^ 1'h1;
  assign T238 = s2_tag_match_way[2'h3:2'h3];
  assign T239 = T253 | T240;
  assign T240 = T252 ? s2_data_2 : 128'h0;
  assign s2_data_2 = T241;
  assign T241 = T242;
  assign T242 = {R248, R243};
  assign T435 = T244[6'h3f:1'h0];
  assign T244 = T246 ? T245 : T436;
  assign T436 = {64'h0, R243};
  assign T245 = data_io_resp_2 >> 1'h0;
  assign T246 = s1_clk_en & T247;
  assign T247 = s1_tag_eq_way[2'h2:2'h2];
  assign T249 = T251 ? T250 : R248;
  assign T250 = data_io_resp_2 >> 7'h40;
  assign T251 = T246 & s1_writeback;
  assign T252 = s2_tag_match_way[2'h2:2'h2];
  assign T253 = T267 | T254;
  assign T254 = T266 ? s2_data_1 : 128'h0;
  assign s2_data_1 = T255;
  assign T255 = T256;
  assign T256 = {R262, R257};
  assign T437 = T258[6'h3f:1'h0];
  assign T258 = T260 ? T259 : T438;
  assign T438 = {64'h0, R257};
  assign T259 = data_io_resp_1 >> 1'h0;
  assign T260 = s1_clk_en & T261;
  assign T261 = s1_tag_eq_way[1'h1:1'h1];
  assign T263 = T265 ? T264 : R262;
  assign T264 = data_io_resp_1 >> 7'h40;
  assign T265 = T260 & s1_writeback;
  assign T266 = s2_tag_match_way[1'h1:1'h1];
  assign T267 = T279 ? s2_data_0 : 128'h0;
  assign s2_data_0 = T268;
  assign T268 = T269;
  assign T269 = {R275, R270};
  assign T439 = T271[6'h3f:1'h0];
  assign T271 = T273 ? T272 : T440;
  assign T440 = {64'h0, R270};
  assign T272 = data_io_resp_0 >> 1'h0;
  assign T273 = s1_clk_en & T274;
  assign T274 = s1_tag_eq_way[1'h0:1'h0];
  assign T276 = T278 ? T277 : R275;
  assign T277 = data_io_resp_0 >> 7'h40;
  assign T278 = T273 & s1_writeback;
  assign T279 = s2_tag_match_way[1'h0:1'h0];
  assign T280 = s2_data_muxed[7'h7f:7'h40];
  assign T441 = {64'h0, s2_store_bypass_data};
  assign T281 = T341 ? T282 : s2_store_bypass_data;
  assign T282 = T326 ? amoalu_io_out : T283;
  assign T283 = T312 ? s3_req_data : s4_req_data;
  assign T284 = T285 ? s3_req_data : s4_req_data;
  assign T285 = s3_valid & metaReadArb_io_out_valid;
  assign T442 = reset ? 1'h0 : T286;
  assign T286 = T294 & T287;
  assign T287 = T291 | T288;
  assign T288 = T290 | T289;
  assign T289 = s2_req_cmd == 5'h4;
  assign T290 = s2_req_cmd[2'h3:2'h3];
  assign T291 = T293 | T292;
  assign T292 = s2_req_cmd == 5'h7;
  assign T293 = s2_req_cmd == 5'h1;
  assign T294 = T296 & T295;
  assign T295 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T206;
  assign T206 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T207;
  assign T207 = lrsc_addr == T208;
  assign T208 = s2_req_addr >> 3'h6;
  assign T209 = T17 ? T210 : lrsc_addr;
  assign T210 = s2_req_addr >> 3'h6;
  assign T17 = T124 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T124 = T125 | s2_replay;
  assign T125 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T126;
  assign T126 = s2_valid & T127;
  assign T127 = s2_nack ^ 1'h1;
  assign s2_nack = T130 | s2_nack_miss;
  assign s2_nack_miss = T129 & T128;
  assign T128 = mshrs_io_req_ready ^ 1'h1;
  assign T129 = s2_hit ^ 1'h1;
  assign T130 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T131 = T137 ? s1_nack : s2_nack_hit;
  assign s1_nack = T136 | T132;
  assign T132 = T134 & T133;
  assign T133 = prober_io_req_ready ^ 1'h1;
  assign T134 = T135 == prober_io_meta_write_bits_idx;
  assign T135 = s1_req_addr[4'hc:3'h6];
  assign T136 = T492 & dtlb_io_resp_miss;
  assign T137 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T422 = reset ? 5'h0 : T10;
  assign T10 = io_cpu_ptw_sret ? 5'h0 : T11;
  assign T11 = T138 ? 5'h0 : T12;
  assign T12 = T15 ? 5'h1f : T13;
  assign T13 = lrsc_valid ? T14 : lrsc_count;
  assign T14 = lrsc_count - 5'h1;
  assign T15 = T17 & T16;
  assign T16 = lrsc_valid ^ 1'h1;
  assign T138 = T124 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T296 = T297 | s2_replay;
  assign T297 = s2_valid_masked & s2_hit;
  assign T443 = T298[6'h3f:1'h0];
  assign T298 = T302 ? T300 : T444;
  assign T444 = {64'h0, T299};
  assign T299 = T302 ? s2_req_data : s3_req_data;
  assign T300 = s2_data_correctable ? s2_data_corrected : T445;
  assign T445 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T301;
  assign T301 = {T280, T222};
  assign T302 = T311 & T303;
  assign T303 = T304 | s2_data_correctable;
  assign T304 = T308 | T305;
  assign T305 = T307 | T306;
  assign T306 = s2_req_cmd == 5'h4;
  assign T307 = s2_req_cmd[2'h3:2'h3];
  assign T308 = T310 | T309;
  assign T309 = s2_req_cmd == 5'h7;
  assign T310 = s2_req_cmd == 5'h1;
  assign T311 = s2_valid | s2_replay;
  assign T312 = T321 & T313;
  assign T313 = T318 | T314;
  assign T314 = T317 | T315;
  assign T315 = s3_req_cmd == 5'h4;
  assign T316 = T302 ? s2_req_cmd : s3_req_cmd;
  assign T317 = s3_req_cmd[2'h3:2'h3];
  assign T318 = T320 | T319;
  assign T319 = s3_req_cmd == 5'h7;
  assign T320 = s3_req_cmd == 5'h1;
  assign T321 = s3_valid & T322;
  assign T322 = T446 == T323;
  assign T323 = s3_req_addr >> 2'h3;
  assign T324 = T302 ? s2_req_addr : s3_req_addr;
  assign T446 = {12'h0, T325};
  assign T325 = s1_addr >> 2'h3;
  assign T326 = T334 & T327;
  assign T327 = T331 | T328;
  assign T328 = T330 | T329;
  assign T329 = s2_req_cmd == 5'h4;
  assign T330 = s2_req_cmd[2'h3:2'h3];
  assign T331 = T333 | T332;
  assign T332 = s2_req_cmd == 5'h7;
  assign T333 = s2_req_cmd == 5'h1;
  assign T334 = T338 & T335;
  assign T335 = T447 == T336;
  assign T336 = s2_req_addr >> 2'h3;
  assign T447 = {12'h0, T337};
  assign T337 = s1_addr >> 2'h3;
  assign T338 = T340 & T339;
  assign T339 = s2_sc_fail ^ 1'h1;
  assign T340 = s2_valid_masked | s2_replay;
  assign T341 = s1_clk_en & T342;
  assign T342 = T357 | T343;
  assign T343 = T352 & T344;
  assign T344 = T349 | T345;
  assign T345 = T348 | T346;
  assign T346 = s4_req_cmd == 5'h4;
  assign T347 = T285 ? s3_req_cmd : s4_req_cmd;
  assign T348 = s4_req_cmd[2'h3:2'h3];
  assign T349 = T351 | T350;
  assign T350 = s4_req_cmd == 5'h7;
  assign T351 = s4_req_cmd == 5'h1;
  assign T352 = s4_valid & T353;
  assign T353 = T448 == T354;
  assign T354 = s4_req_addr >> 2'h3;
  assign T355 = T285 ? s3_req_addr : s4_req_addr;
  assign T448 = {12'h0, T356};
  assign T356 = s1_addr >> 2'h3;
  assign T449 = reset ? 1'h0 : s3_valid;
  assign T357 = T326 | T312;
  assign T358 = T341 ? 1'h1 : T359;
  assign T359 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T175 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T172 = s2_recycle ? s2_req_typ : T173;
  assign T173 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T174;
  assign T174 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T461 = s2_req_cmd[2'h3:1'h0];
  assign T462 = s2_req_addr[3'h5:1'h0];
  assign T463 = {s3_req_data, s3_req_data};
  assign T464 = 1'h1 << T465;
  assign T465 = T466;
  assign T466 = s3_req_addr[2'h3:2'h3];
  assign T467 = s3_req_addr[4'hc:1'h0];
  assign T468 = T302 ? s2_tag_match_way : s3_way;
  assign T469 = FlowThroughSerializer_0_io_out_bits_payload_data[7'h7f:1'h0];
  assign T470 = FlowThroughSerializer_0_io_out_valid & T471;
  assign T471 = T473 | T472;
  assign T472 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h2;
  assign T473 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h1;
  assign T474 = T475 | T454;
  assign T475 = FlowThroughSerializer_0_io_out_valid ^ 1'h1;
  assign T476 = s2_req_addr[4'hc:1'h0];
  assign T477 = mshrs_io_replay_bits_addr[4'hc:1'h0];
  assign T478 = io_cpu_req_bits_addr[4'hc:1'h0];
  assign T479 = T480;
  assign T480 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T481 = T482[3'h6:1'h0];
  assign T482 = s2_req_addr >> 3'h6;
  assign T483 = T484[3'h6:1'h0];
  assign T484 = io_cpu_req_bits_addr >> 3'h6;
  assign T485 = s2_recycle ? s2_req_phys : T486;
  assign T486 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T487;
  assign T487 = prober_io_meta_read_valid ? 1'h1 : T488;
  assign T488 = wb_io_meta_read_valid ? 1'h1 : T489;
  assign T489 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T490 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T491 = s1_req_addr >> 4'hd;
  assign T492 = T494 & T493;
  assign T493 = s1_req_phys ^ 1'h1;
  assign T494 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T498 | T495;
  assign T495 = T497 | T496;
  assign T496 = s1_req_cmd == 5'h3;
  assign T497 = s1_req_cmd == 5'h2;
  assign T498 = s1_read | s1_write;
  assign s1_read = T164 | T161;
  assign T161 = T163 | T162;
  assign T162 = s1_req_cmd == 5'h4;
  assign T163 = s1_req_cmd[2'h3:2'h3];
  assign T164 = T166 | T165;
  assign T165 = s1_req_cmd == 5'h6;
  assign T166 = s1_req_cmd == 5'h0;
  assign T499 = T454 & FlowThroughSerializer_0_io_out_valid;
  assign T500 = io_mem_acquire_ready;
  assign T501 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R502;
  assign T503 = s1_clk_en ? T504 : R502;
  assign T504 = R505[1'h1:1'h0];
  assign T506 = reset ? 16'h1 : T507;
  assign T507 = T517 ? T508 : R505;
  assign T508 = {T510, T509};
  assign T509 = R505[4'hf:1'h1];
  assign T510 = T512 ^ T511;
  assign T511 = R505[3'h5:3'h5];
  assign T512 = T514 ^ T513;
  assign T513 = R505[2'h3:2'h3];
  assign T514 = T516 ^ T515;
  assign T515 = R505[2'h2:2'h2];
  assign T516 = R505[1'h0:1'h0];
  assign T517 = T518;
  assign T518 = mshrs_io_req_ready & T573;
  assign T519 = s2_tag_match ? T565 : T520;
  assign T520 = T521[1'h1:1'h0];
  assign T521 = T533 | T522;
  assign T522 = T532 ? T523 : 21'h0;
  assign T523 = T524;
  assign T524 = {R530, R525};
  assign T526 = T527 ? meta_io_resp_3_coh_state : R525;
  assign T527 = s1_clk_en & T528;
  assign T528 = s1_replaced_way_en[2'h3:2'h3];
  assign s1_replaced_way_en = 1'h1 << T529;
  assign T529 = R505[1'h1:1'h0];
  assign T531 = T527 ? meta_io_resp_3_tag : R530;
  assign T532 = s2_replaced_way_en[2'h3:2'h3];
  assign T533 = T544 | T534;
  assign T534 = T543 ? T535 : 21'h0;
  assign T535 = T536;
  assign T536 = {R541, R537};
  assign T538 = T539 ? meta_io_resp_2_coh_state : R537;
  assign T539 = s1_clk_en & T540;
  assign T540 = s1_replaced_way_en[2'h2:2'h2];
  assign T542 = T539 ? meta_io_resp_2_tag : R541;
  assign T543 = s2_replaced_way_en[2'h2:2'h2];
  assign T544 = T555 | T545;
  assign T545 = T554 ? T546 : 21'h0;
  assign T546 = T547;
  assign T547 = {R552, R548};
  assign T549 = T550 ? meta_io_resp_1_coh_state : R548;
  assign T550 = s1_clk_en & T551;
  assign T551 = s1_replaced_way_en[1'h1:1'h1];
  assign T553 = T550 ? meta_io_resp_1_tag : R552;
  assign T554 = s2_replaced_way_en[1'h1:1'h1];
  assign T555 = T564 ? T556 : 21'h0;
  assign T556 = T557;
  assign T557 = {R562, R558};
  assign T559 = T560 ? meta_io_resp_0_coh_state : R558;
  assign T560 = s1_clk_en & T561;
  assign T561 = s1_replaced_way_en[1'h0:1'h0];
  assign T563 = T560 ? meta_io_resp_0_tag : R562;
  assign T564 = s2_replaced_way_en[1'h0:1'h0];
  assign T565 = T41;
  assign T566 = s2_tag_match ? T568 : T567;
  assign T567 = T521[5'h14:2'h2];
  assign T568 = T567;
  assign T193 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T190 = s2_recycle ? s2_req_tag : T191;
  assign T191 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T192;
  assign T192 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T569 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T570 = s2_recycle ? s2_req_kill : T571;
  assign T571 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T572;
  assign T572 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T573 = s2_nack_hit ? 1'h0 : T574;
  assign T574 = T594 & T575;
  assign T575 = T583 | T576;
  assign T576 = T580 | T577;
  assign T577 = T579 | T578;
  assign T578 = s2_req_cmd == 5'h4;
  assign T579 = s2_req_cmd[2'h3:2'h3];
  assign T580 = T582 | T581;
  assign T581 = s2_req_cmd == 5'h7;
  assign T582 = s2_req_cmd == 5'h1;
  assign T583 = T591 | T584;
  assign T584 = T588 | T585;
  assign T585 = T587 | T586;
  assign T586 = s2_req_cmd == 5'h4;
  assign T587 = s2_req_cmd[2'h3:2'h3];
  assign T588 = T590 | T589;
  assign T589 = s2_req_cmd == 5'h6;
  assign T590 = s2_req_cmd == 5'h0;
  assign T591 = T593 | T592;
  assign T592 = s2_req_cmd == 5'h3;
  assign T593 = s2_req_cmd == 5'h2;
  assign T594 = s2_valid_masked & T595;
  assign T595 = s2_hit ^ 1'h1;
  assign probe_bits_p_type = io_mem_probe_bits_payload_p_type;
  assign probe_bits_master_xact_id = io_mem_probe_bits_payload_master_xact_id;
  assign probe_bits_addr = io_mem_probe_bits_payload_addr;
  assign T596 = probe_valid & T597;
  assign T597 = lrsc_valid ^ 1'h1;
  assign probe_valid = io_mem_probe_valid;
  assign io_mem_release_bits_payload_r_type = T0;
  assign T0 = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_payload_data = T1;
  assign T1 = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_payload_master_xact_id = T2;
  assign T2 = releaseArb_io_out_bits_master_xact_id;
  assign io_mem_release_bits_payload_client_xact_id = T3;
  assign T3 = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_payload_addr = T4;
  assign T4 = releaseArb_io_out_bits_addr;
  assign io_mem_release_bits_header_dst = T5;
  assign T5 = 2'h0;
  assign io_mem_release_bits_header_src = T6;
  assign T6 = 2'h0;
  assign io_mem_release_valid = T7;
  assign T7 = releaseArb_io_out_valid;
  assign io_mem_probe_ready = probe_ready;
  assign probe_ready = T8;
  assign T8 = prober_io_req_ready & T9;
  assign T9 = lrsc_valid ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = mshrs_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mshrs_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = mshrs_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_0_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T139;
  assign T139 = mshrs_io_mem_req_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = T140;
  assign T140 = mshrs_io_mem_req_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = T141;
  assign T141 = mshrs_io_mem_req_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = T142;
  assign T142 = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_payload_data = T143;
  assign T143 = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_payload_client_xact_id = T144;
  assign T144 = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = T145;
  assign T145 = mshrs_io_mem_req_bits_addr;
  assign io_mem_acquire_bits_header_dst = T146;
  assign T146 = 2'h0;
  assign io_mem_acquire_bits_header_src = T147;
  assign T147 = 2'h0;
  assign io_mem_acquire_valid = T148;
  assign T148 = mshrs_io_mem_req_valid;
  assign io_cpu_ordered = T149;
  assign T149 = T151 & T150;
  assign T150 = s2_valid ^ 1'h1;
  assign T151 = mshrs_io_fence_rdy & T152;
  assign T152 = s1_valid ^ 1'h1;
  assign io_cpu_ptw_req_bits = dtlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_xcpt_pf_st = T153;
  assign T153 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T160;
  assign T160 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T167;
  assign T167 = s1_write & misaligned;
  assign misaligned = T176 | T168;
  assign T168 = T171 & T169;
  assign T169 = T170 != 3'h0;
  assign T170 = s1_req_addr[2'h2:1'h0];
  assign T171 = s1_req_typ == 3'h3;
  assign T176 = T183 | T177;
  assign T177 = T180 & T178;
  assign T178 = T179 != 2'h0;
  assign T179 = s1_req_addr[1'h1:1'h0];
  assign T180 = T182 | T181;
  assign T181 = s1_req_typ == 3'h6;
  assign T182 = s1_req_typ == 3'h2;
  assign T183 = T186 & T184;
  assign T184 = T185 != 1'h0;
  assign T185 = s1_req_addr[1'h0:1'h0];
  assign T186 = T188 | T187;
  assign T187 = s1_req_typ == 3'h5;
  assign T188 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T189;
  assign T189 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T194;
  assign T194 = s1_replay & T195;
  assign T195 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_cmd = T431;
  assign T431 = s2_req_cmd[2'h3:1'h0];
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data_subword = T205;
  assign T205 = T211 | T432;
  assign T432 = {63'h0, s2_sc_fail};
  assign T211 = {T389, T212};
  assign T212 = s2_sc ? 8'h0 : T213;
  assign T213 = T388 ? T387 : T214;
  assign T214 = T215[3'h7:1'h0];
  assign T215 = {T379, T216};
  assign T216 = T378 ? T377 : T217;
  assign T217 = T218[4'hf:1'h0];
  assign T218 = {T362, T219};
  assign T219 = T361 ? T360 : T220;
  assign T220 = s2_data_word[5'h1f:1'h0];
  assign T360 = s2_data_word[6'h3f:6'h20];
  assign T361 = s2_req_addr[2'h2:2'h2];
  assign T362 = T374 ? T364 : T363;
  assign T363 = s2_data_word[6'h3f:6'h20];
  assign T364 = 32'h0 - T450;
  assign T450 = {31'h0, T365};
  assign T365 = T367 & T366;
  assign T366 = T219[5'h1f:5'h1f];
  assign T367 = T369 | T368;
  assign T368 = s2_req_typ == 3'h3;
  assign T369 = T371 | T370;
  assign T370 = s2_req_typ == 3'h2;
  assign T371 = T373 | T372;
  assign T372 = s2_req_typ == 3'h1;
  assign T373 = s2_req_typ == 3'h0;
  assign T374 = T376 | T375;
  assign T375 = s2_req_typ == 3'h6;
  assign T376 = s2_req_typ == 3'h2;
  assign T377 = T218[5'h1f:5'h10];
  assign T378 = s2_req_addr[1'h1:1'h1];
  assign T379 = T384 ? T381 : T380;
  assign T380 = T218[6'h3f:5'h10];
  assign T381 = 48'h0 - T451;
  assign T451 = {47'h0, T382};
  assign T382 = T367 & T383;
  assign T383 = T216[4'hf:4'hf];
  assign T384 = T386 | T385;
  assign T385 = s2_req_typ == 3'h5;
  assign T386 = s2_req_typ == 3'h1;
  assign T387 = T215[4'hf:4'h8];
  assign T388 = s2_req_addr[1'h0:1'h0];
  assign T389 = T394 ? T391 : T390;
  assign T390 = T215[6'h3f:4'h8];
  assign T391 = 56'h0 - T452;
  assign T452 = {55'h0, T392};
  assign T392 = T367 & T393;
  assign T393 = T212[3'h7:3'h7];
  assign T394 = s2_sc | T395;
  assign T395 = T397 | T396;
  assign T396 = s2_req_typ == 3'h4;
  assign T397 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_data = T218;
  assign io_cpu_resp_bits_has_data = T398;
  assign T398 = T399 | s2_sc;
  assign T399 = T403 | T400;
  assign T400 = T402 | T401;
  assign T401 = s2_req_cmd == 5'h4;
  assign T402 = s2_req_cmd[2'h3:2'h3];
  assign T403 = T405 | T404;
  assign T404 = s2_req_cmd == 5'h6;
  assign T405 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T406;
  assign T406 = s2_valid & s2_nack;
  assign io_cpu_resp_valid = T407;
  assign T407 = T409 & T408;
  assign T408 = s2_data_correctable ^ 1'h1;
  assign T409 = s2_replay | T410;
  assign T410 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T411;
  assign T411 = block_miss ? 1'h0 : T412;
  assign T412 = T419 ? 1'h0 : T413;
  assign T413 = T418 ? 1'h0 : T414;
  assign T414 = T415 == 1'h0;
  assign T415 = T417 & T416;
  assign T416 = io_cpu_req_bits_phys ^ 1'h1;
  assign T417 = dtlb_io_req_ready ^ 1'h1;
  assign T418 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T419 = readArb_io_in_3_ready ^ 1'h1;
  assign T453 = reset ? 1'h0 : T420;
  assign T420 = T421 & s2_nack_miss;
  assign T421 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_tag( wbArb_io_out_bits_tag ),
       .io_req_bits_idx( wbArb_io_out_bits_idx ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr( wb_io_release_bits_addr ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T596 ),
       .io_req_bits_addr( probe_bits_addr ),
       .io_req_bits_master_xact_id( probe_bits_master_xact_id ),
       .io_req_bits_p_type( probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr( prober_io_rep_bits_addr ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_tag( prober_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( prober_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_line_state_state( T41 )
  );
  `ifndef SYNTHESIS
    assign prober.io_req_bits_client_xact_id = {1{$random}};
  `endif
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T573 ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T566 ),
       .io_req_bits_old_meta_coh_state( T519 ),
       .io_req_bits_way_en( T501 ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( T500 ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr( mshrs_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_write_mask( mshrs_io_mem_req_bits_write_mask ),
       .io_mem_req_bits_subword_addr( mshrs_io_mem_req_bits_subword_addr ),
       .io_mem_req_bits_atomic_opcode( mshrs_io_mem_req_bits_atomic_opcode ),
       .io_mem_resp_way_en( mshrs_io_mem_resp_way_en ),
       .io_mem_resp_addr( mshrs_io_mem_resp_addr ),
       //.io_mem_resp_wmask(  )
       //.io_mem_resp_data(  )
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       //.io_replay_bits_sdq_id(  )
       .io_mem_grant_valid( T499 ),
       .io_mem_grant_bits_header_src( FlowThroughSerializer_0_io_out_bits_header_src ),
       .io_mem_grant_bits_header_dst( FlowThroughSerializer_0_io_out_bits_header_dst ),
       .io_mem_grant_bits_payload_data( FlowThroughSerializer_0_io_out_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( FlowThroughSerializer_0_io_out_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( FlowThroughSerializer_0_io_out_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( FlowThroughSerializer_0_io_out_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( mshrs_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( mshrs_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( mshrs_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( mshrs_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T492 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T491 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_resp_miss( dtlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits( dtlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_3_tag( meta_io_resp_3_tag ),
       .io_resp_3_coh_state( meta_io_resp_3_coh_state ),
       .io_resp_2_tag( meta_io_resp_2_tag ),
       .io_resp_2_coh_state( meta_io_resp_2_coh_state ),
       .io_resp_1_tag( meta_io_resp_1_tag ),
       .io_resp_1_coh_state( meta_io_resp_1_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T483 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T481 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T479 ),
       .io_resp_3( data_io_resp_3 ),
       .io_resp_2( data_io_resp_2 ),
       .io_resp_1( data_io_resp_1 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 4'hf ),
       .io_in_3_bits_addr( T478 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 4'hf ),
       .io_in_1_bits_addr( T477 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 4'hf ),
       .io_in_0_bits_addr( T476 ),
       .io_out_ready( T474 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T470 ),
       .io_in_1_bits_way_en( mshrs_io_mem_resp_way_en ),
       .io_in_1_bits_addr( mshrs_io_mem_resp_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( T469 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T467 ),
       .io_in_0_bits_wmask( T464 ),
       .io_in_0_bits_data( T463 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T462 ),
       .io_cmd( T461 ),
       .io_typ( s2_req_typ ),
       .io_lhs( T460 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  Arbiter_4 releaseArb(
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr( prober_io_rep_bits_addr ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr( wb_io_release_bits_addr ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_out_ready( T459 ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr( releaseArb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( releaseArb_io_out_bits_master_xact_id ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  FlowThroughSerializer_0 FlowThroughSerializer_0(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_0_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( T454 ),
       .io_out_valid( FlowThroughSerializer_0_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( FlowThroughSerializer_0_io_out_bits_header_dst ),
       .io_out_bits_payload_data( FlowThroughSerializer_0_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( FlowThroughSerializer_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_0_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_5 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_tag( prober_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( prober_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_tag( wbArb_io_out_bits_tag ),
       .io_out_bits_idx( wbArb_io_out_bits_idx ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(T203) begin
      s2_req_data <= s1_req_data;
    end else if(T199) begin
      s2_req_data <= T198;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T26;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T28) begin
      s2_recycle_next <= T24;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T27;
    end
    if(s1_clk_en) begin
      R45 <= meta_io_resp_3_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T427;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T426;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T428;
    end
    if(s1_clk_en) begin
      R89 <= meta_io_resp_2_coh_state;
    end
    if(s1_clk_en) begin
      R95 <= meta_io_resp_1_coh_state;
    end
    if(s1_clk_en) begin
      R100 <= meta_io_resp_0_coh_state;
    end
    if(reset) begin
      R122 <= 1'h0;
    end else begin
      R122 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R226 <= T433;
    if(T234) begin
      R231 <= T233;
    end
    R243 <= T435;
    if(T251) begin
      R248 <= T250;
    end
    R257 <= T437;
    if(T265) begin
      R262 <= T264;
    end
    R270 <= T439;
    if(T278) begin
      R275 <= T277;
    end
    if(T341) begin
      s2_store_bypass_data <= T282;
    end
    if(T285) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T286;
    end
    if(T17) begin
      lrsc_addr <= T210;
    end
    if(T137) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_ptw_sret) begin
      lrsc_count <= 5'h0;
    end else if(T138) begin
      lrsc_count <= 5'h0;
    end else if(T15) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T14;
    end
    s3_req_data <= T443;
    if(T302) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T302) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T285) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T285) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T341) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T302) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R502 <= T504;
    end
    if(reset) begin
      R505 <= 16'h1;
    end else if(T517) begin
      R505 <= T508;
    end
    if(T527) begin
      R525 <= meta_io_resp_3_coh_state;
    end
    if(T527) begin
      R530 <= meta_io_resp_3_tag;
    end
    if(T539) begin
      R537 <= meta_io_resp_2_coh_state;
    end
    if(T539) begin
      R541 <= meta_io_resp_2_tag;
    end
    if(T550) begin
      R548 <= meta_io_resp_1_coh_state;
    end
    if(T550) begin
      R552 <= meta_io_resp_1_tag;
    end
    if(T560) begin
      R558 <= meta_io_resp_0_coh_state;
    end
    if(T560) begin
      R562 <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T420;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [29:0] io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [29:0] io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output[29:0] io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T28;
  wire T6;
  wire T7;
  wire[29:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T28 = reset ? 1'h0 : T6;
  assign T6 = T7 ? T0 : R5;
  assign T7 = io_out_ready & io_out_valid;
  assign io_out_bits = T8;
  assign T8 = T9 ? io_in_1_bits : io_in_0_bits;
  assign T9 = T0;
  assign io_out_valid = T10;
  assign T10 = T9 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T19 | T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T17 | T15;
  assign T15 = io_in_1_valid & T16;
  assign T16 = R5 < 1'h1;
  assign T17 = io_in_0_valid & T18;
  assign T18 = R5 < 1'h0;
  assign T19 = R5 < 1'h0;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T25 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T24 | io_in_0_valid;
  assign T24 = T17 | T15;
  assign T25 = T27 & T26;
  assign T26 = R5 < 1'h1;
  assign T27 = T17 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T7) begin
      R5 <= T0;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [29:0] io_requestor_1_req_bits,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[18:0] io_requestor_1_resp_bits_ppn,
    output[5:0] io_requestor_1_resp_bits_perm,
    output[7:0] io_requestor_1_status_ip,
    output[7:0] io_requestor_1_status_im,
    output[6:0] io_requestor_1_status_zero,
    output io_requestor_1_status_er,
    output io_requestor_1_status_vm,
    output io_requestor_1_status_s64,
    output io_requestor_1_status_u64,
    output io_requestor_1_status_ef,
    output io_requestor_1_status_pei,
    output io_requestor_1_status_ei,
    output io_requestor_1_status_ps,
    output io_requestor_1_status_s,
    output io_requestor_1_invalidate,
    output io_requestor_1_sret,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [29:0] io_requestor_0_req_bits,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[18:0] io_requestor_0_resp_bits_ppn,
    output[5:0] io_requestor_0_resp_bits_perm,
    output[7:0] io_requestor_0_status_ip,
    output[7:0] io_requestor_0_status_im,
    output[6:0] io_requestor_0_status_zero,
    output io_requestor_0_status_er,
    output io_requestor_0_status_vm,
    output io_requestor_0_status_s64,
    output io_requestor_0_status_u64,
    output io_requestor_0_status_ef,
    output io_requestor_0_status_pei,
    output io_requestor_0_status_ei,
    output io_requestor_0_status_ps,
    output io_requestor_0_status_s,
    output io_requestor_0_invalidate,
    output io_requestor_0_sret,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    //output[63:0] io_mem_req_bits_data
    //output[7:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    //input  io_mem_ptw_req_valid
    //input [29:0] io_mem_ptw_req_bits
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_sret,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s
);

  wire T79;
  reg [2:0] state;
  wire[2:0] T75;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T14;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T37;
  wire T38;
  wire T39;
  reg [1:0] count;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T36;
  wire T40;
  wire T34;
  wire T35;
  wire[43:0] T74;
  wire[31:0] T0;
  wire[28:0] T1;
  wire[28:0] T2;
  wire[9:0] vpn_idx;
  wire[9:0] T3;
  wire[9:0] T4;
  wire[9:0] T5;
  reg [29:0] r_req_vpn;
  wire[29:0] T6;
  wire T7;
  wire[9:0] T8;
  wire[19:0] T9;
  wire T10;
  wire[1:0] T11;
  wire[9:0] T41;
  wire[29:0] T42;
  wire T43;
  wire[18:0] T44;
  reg [63:0] r_pte;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] T76;
  wire[31:0] T47;
  wire[12:0] T48;
  wire[18:0] T49;
  wire T50;
  wire[5:0] T51;
  wire[18:0] T77;
  wire[30:0] T52;
  wire[30:0] resp_ppn;
  wire[30:0] T53;
  wire[30:0] T54;
  wire[19:0] T55;
  wire[10:0] T56;
  wire[30:0] T57;
  wire[9:0] T58;
  wire[20:0] T59;
  wire T60;
  wire[1:0] T61;
  wire[30:0] r_resp_ppn;
  wire T62;
  wire resp_err;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  reg  r_req_dest;
  wire T67;
  wire resp_val;
  wire T68;
  wire T69;
  wire[5:0] T70;
  wire[18:0] T78;
  wire[30:0] T71;
  wire T72;
  wire T73;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[29:0] arb_io_out_bits;
  wire arb_io_chosen;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    r_req_vpn = {1{$random}};
    r_pte = {2{$random}};
    r_req_dest = {1{$random}};
  end
`endif

  assign T79 = state == 3'h0;
  assign T75 = reset ? 3'h0 : T15;
  assign T15 = T35 ? 3'h0 : T16;
  assign T16 = T34 ? 3'h0 : T17;
  assign T17 = T37 ? 3'h1 : T18;
  assign T18 = T29 ? 3'h3 : T19;
  assign T19 = T28 ? 3'h4 : T20;
  assign T20 = T26 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h1 : state;
  assign T23 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T24 = T25 & io_mem_req_ready;
  assign T25 = 3'h1 == state;
  assign T26 = T27 & io_mem_resp_bits_nack;
  assign T27 = 3'h2 == state;
  assign T28 = T27 & io_mem_resp_valid;
  assign T29 = T32 & T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_mem_resp_bits_data[1'h1:1'h1];
  assign T32 = T28 & T33;
  assign T33 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T37 = T32 & T38;
  assign T38 = T40 & T39;
  assign T39 = count < 2'h2;
  assign T12 = T37 ? T36 : T13;
  assign T13 = T14 ? 2'h0 : count;
  assign T36 = count + 2'h1;
  assign T40 = T30 ^ 1'h1;
  assign T34 = 3'h3 == state;
  assign T35 = 3'h4 == state;
  assign io_mem_req_bits_cmd = 5'h0;
  assign io_mem_req_bits_addr = T74;
  assign T74 = {12'h0, T0};
  assign T0 = T1 << 2'h3;
  assign T1 = T2;
  assign T2 = {T44, vpn_idx};
  assign vpn_idx = T43 ? T41 : T3;
  assign T3 = T10 ? T8 : T4;
  assign T4 = T5[4'h9:1'h0];
  assign T5 = r_req_vpn >> 5'h14;
  assign T6 = T7 ? arb_io_out_bits : r_req_vpn;
  assign T7 = T79 & arb_io_out_valid;
  assign T8 = T9[4'h9:1'h0];
  assign T9 = r_req_vpn >> 4'ha;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = count;
  assign T41 = T42[4'h9:1'h0];
  assign T42 = r_req_vpn >> 1'h0;
  assign T43 = T11[1'h1:1'h1];
  assign T44 = r_pte[5'h1f:4'hd];
  assign T45 = io_mem_resp_valid ? io_mem_resp_bits_data : T46;
  assign T46 = T7 ? T76 : r_pte;
  assign T76 = {32'h0, T47};
  assign T47 = {T49, T48};
  assign T48 = io_mem_resp_bits_data[4'hc:1'h0];
  assign T49 = io_dpath_ptbr[5'h1f:4'hd];
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T50;
  assign T50 = state == 3'h1;
  assign io_requestor_0_sret = io_dpath_sret;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_s = io_dpath_status_s;
  assign io_requestor_0_status_ps = io_dpath_status_ps;
  assign io_requestor_0_status_ei = io_dpath_status_ei;
  assign io_requestor_0_status_pei = io_dpath_status_pei;
  assign io_requestor_0_status_ef = io_dpath_status_ef;
  assign io_requestor_0_status_u64 = io_dpath_status_u64;
  assign io_requestor_0_status_s64 = io_dpath_status_s64;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_er = io_dpath_status_er;
  assign io_requestor_0_status_zero = io_dpath_status_zero;
  assign io_requestor_0_status_im = io_dpath_status_im;
  assign io_requestor_0_status_ip = io_dpath_status_ip;
  assign io_requestor_0_resp_bits_perm = T51;
  assign T51 = r_pte[4'h8:2'h3];
  assign io_requestor_0_resp_bits_ppn = T77;
  assign T77 = T52[5'h12:1'h0];
  assign T52 = resp_ppn;
  assign resp_ppn = T62 ? r_resp_ppn : T53;
  assign T53 = T60 ? T57 : T54;
  assign T54 = {T56, T55};
  assign T55 = r_req_vpn[5'h13:1'h0];
  assign T56 = r_resp_ppn >> 5'h14;
  assign T57 = {T59, T58};
  assign T58 = r_req_vpn[4'h9:1'h0];
  assign T59 = r_resp_ppn >> 4'ha;
  assign T60 = T61[1'h0:1'h0];
  assign T61 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hd;
  assign T62 = T61[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = T64 | T63;
  assign T63 = state == 3'h2;
  assign T64 = state == 3'h4;
  assign io_requestor_0_resp_valid = T65;
  assign T65 = resp_val & T66;
  assign T66 = r_req_dest == 1'h0;
  assign T67 = T7 ? arb_io_chosen : r_req_dest;
  assign resp_val = T69 | T68;
  assign T68 = state == 3'h4;
  assign T69 = state == 3'h3;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_sret = io_dpath_sret;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_s = io_dpath_status_s;
  assign io_requestor_1_status_ps = io_dpath_status_ps;
  assign io_requestor_1_status_ei = io_dpath_status_ei;
  assign io_requestor_1_status_pei = io_dpath_status_pei;
  assign io_requestor_1_status_ef = io_dpath_status_ef;
  assign io_requestor_1_status_u64 = io_dpath_status_u64;
  assign io_requestor_1_status_s64 = io_dpath_status_s64;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_er = io_dpath_status_er;
  assign io_requestor_1_status_zero = io_dpath_status_zero;
  assign io_requestor_1_status_im = io_dpath_status_im;
  assign io_requestor_1_status_ip = io_dpath_status_ip;
  assign io_requestor_1_resp_bits_perm = T70;
  assign T70 = r_pte[4'h8:2'h3];
  assign io_requestor_1_resp_bits_ppn = T78;
  assign T78 = T71[5'h12:1'h0];
  assign T71 = resp_ppn;
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T72;
  assign T72 = resp_val & T73;
  assign T73 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits( io_requestor_1_req_bits ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits( io_requestor_0_req_bits ),
       .io_out_ready( T79 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits( arb_io_out_bits ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h0;
    end else if(T37) begin
      state <= 3'h1;
    end else if(T29) begin
      state <= 3'h3;
    end else if(T28) begin
      state <= 3'h4;
    end else if(T26) begin
      state <= 3'h1;
    end else if(T24) begin
      state <= 3'h2;
    end else if(T23) begin
      state <= 3'h1;
    end
    if(T37) begin
      count <= T36;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T7) begin
      r_req_vpn <= arb_io_out_bits;
    end
    if(io_mem_resp_valid) begin
      r_pte <= io_mem_resp_bits_data;
    end else if(T7) begin
      r_pte <= T76;
    end
    if(T7) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module Control(input clk, input reset,
    output[2:0] io_dpath_sel_pc,
    output io_dpath_killd,
    output io_dpath_ren_1,
    output io_dpath_ren_0,
    output[2:0] io_dpath_sel_alu2,
    output[1:0] io_dpath_sel_alu1,
    output[2:0] io_dpath_sel_imm,
    output io_dpath_fn_dw,
    output[3:0] io_dpath_fn_alu,
    output io_dpath_div_mul_val,
    output io_dpath_div_mul_kill,
    //output io_dpath_div_val
    //output io_dpath_div_kill
    output[2:0] io_dpath_csr,
    output io_dpath_sret,
    output io_dpath_mem_load,
    output io_dpath_wb_load,
    output io_dpath_ex_fp_val,
    output io_dpath_mem_fp_val,
    output io_dpath_ex_wen,
    output io_dpath_ex_valid,
    output io_dpath_mem_jalr,
    output io_dpath_mem_branch,
    output io_dpath_mem_wen,
    output io_dpath_wb_wen,
    output[2:0] io_dpath_ex_mem_type,
    output io_dpath_ex_rs2_val,
    output io_dpath_ex_rocc_val,
    output io_dpath_mem_rocc_val,
    output io_dpath_bypass_1,
    output io_dpath_bypass_0,
    output[1:0] io_dpath_bypass_src_1,
    output[1:0] io_dpath_bypass_src_0,
    output io_dpath_ll_ready,
    output io_dpath_retire,
    output io_dpath_exception,
    output[63:0] io_dpath_cause,
    output io_dpath_badvaddr_wen,
    input [31:0] io_dpath_inst,
    //input  io_dpath_jalr_eq
    input  io_dpath_mem_br_taken,
    input  io_dpath_mem_misprediction,
    input  io_dpath_div_mul_rdy,
    input  io_dpath_ll_wen,
    input [4:0] io_dpath_ll_waddr,
    input [4:0] io_dpath_ex_waddr,
    input  io_dpath_mem_rs1_ra,
    input [4:0] io_dpath_mem_waddr,
    input [4:0] io_dpath_wb_waddr,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s,
    input  io_dpath_fp_sboard_clr,
    input [4:0] io_dpath_fp_sboard_clra,
    input  io_dpath_csr_replay,
    output io_imem_req_valid,
    //output[43:0] io_imem_req_bits_pc
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_btb_update_bits_pc
    //output[42:0] io_imem_btb_update_bits_target
    //output[42:0] io_imem_btb_update_bits_returnAddr
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_mispredict,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    //output[43:0] io_dmem_req_bits_addr
    //output[63:0] io_dmem_req_bits_data
    //output[7:0] io_dmem_req_bits_tag
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output io_fpu_valid,
    input  io_fpu_fcsr_rdy,
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    input [4:0] io_fpu_dec_cmd,
    input  io_fpu_dec_ldst,
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    input  io_fpu_dec_swap23,
    input  io_fpu_dec_single,
    input  io_fpu_dec_fromint,
    input  io_fpu_dec_toint,
    input  io_fpu_dec_fastpipe,
    input  io_fpu_dec_fma,
    input  io_fpu_dec_round,
    input  io_fpu_sboard_set,
    input  io_fpu_sboard_clr,
    input [4:0] io_fpu_sboard_clra,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire T0;
  reg  wb_reg_xcpt;
  wire T1;
  wire T2;
  wire take_pc_wb;
  wire T3;
  reg  wb_reg_sret;
  wire T4;
  wire T5;
  wire T6;
  reg  mem_reg_replay;
  wire T7;
  wire replay_ex;
  wire replay_ex_other;
  reg  mem_reg_replay_next;
  wire T8;
  reg  ex_reg_replay_next;
  wire T9;
  wire T10;
  wire id_csr_flush;
  wire T11;
  wire T12;
  wire T13;
  wire[11:0] T14;
  wire[11:0] id_csr_addr;
  wire T15;
  wire[11:0] T16;
  wire T17;
  wire id_csr_wen;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] id_csr;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[4:0] id_raddr1;
  wire id_csr_en;
  wire id_replay_next;
  wire[31:0] T27;
  wire ctrl_killd;
  wire T28;
  wire ctrl_draind;
  wire id_interrupt;
  wire id_interrupt_unmasked;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire ctrl_stalld;
  wire id_do_fence;
  wire T60;
  wire T61;
  wire T62;
  wire id_mem_val;
  wire T63;
  wire[31:0] T64;
  wire T65;
  wire T66;
  wire[31:0] T67;
  wire T68;
  wire T69;
  wire[31:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T76;
  wire T77;
  wire T78;
  wire[31:0] T79;
  wire T80;
  wire[31:0] T81;
  reg  id_reg_fence;
  wire T793;
  wire T82;
  wire T83;
  wire id_fence_next;
  wire T84;
  wire id_amo_rl;
  wire id_amo;
  wire[31:0] T85;
  wire id_fence;
  wire[31:0] T86;
  wire T87;
  wire id_fence_i;
  wire[31:0] T88;
  wire T89;
  wire id_amo_aq;
  wire id_mem_busy;
  reg  ex_reg_mem_val;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire id_stall_fpu;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[4:0] T102;
  wire[4:0] T103;
  wire[4:0] id_waddr;
  wire T104;
  reg [31:0] R105;
  wire[31:0] T794;
  wire[31:0] T106;
  wire[31:0] T107;
  wire[31:0] T108;
  wire[31:0] T109;
  wire[31:0] T110;
  wire[31:0] T111;
  wire T112;
  wire T113;
  wire replay_wb;
  wire T114;
  wire T115;
  reg  wb_reg_rocc_val;
  wire T116;
  reg  mem_reg_rocc_val;
  wire T117;
  reg  ex_reg_rocc_val;
  wire T118;
  wire T119;
  wire replay_wb_common;
  wire T120;
  reg  wb_reg_replay;
  wire T121;
  wire T122;
  wire replay_mem;
  wire fpu_kill_mem;
  reg  mem_reg_fp_val;
  wire T123;
  reg  ex_reg_fp_val;
  wire T124;
  wire T125;
  wire dcache_kill_mem;
  reg  mem_reg_wen;
  wire T126;
  reg  ex_reg_wen;
  wire T127;
  wire id_wen;
  wire T128;
  wire[31:0] T129;
  wire T130;
  wire T131;
  wire[31:0] T132;
  wire T133;
  wire T134;
  wire[31:0] T135;
  wire T136;
  wire T137;
  wire[31:0] T138;
  wire T139;
  wire T140;
  wire[31:0] T141;
  wire T142;
  wire T143;
  wire[31:0] T144;
  wire T145;
  wire[31:0] T146;
  wire T147;
  wire T148;
  reg  wb_reg_fp_wen;
  wire T149;
  reg  mem_reg_fp_wen;
  wire T150;
  reg  ex_reg_fp_wen;
  wire T151;
  wire T152;
  wire wb_dcache_miss;
  wire T153;
  reg  wb_reg_mem_val;
  wire T154;
  reg  mem_reg_mem_val;
  wire T155;
  wire[31:0] T156;
  wire[31:0] T157;
  wire[31:0] T158;
  wire[31:0] T159;
  wire T160;
  wire[31:0] T161;
  wire[31:0] T162;
  wire[31:0] T163;
  wire[31:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire[4:0] T171;
  wire[4:0] T172;
  wire[4:0] id_raddr3;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire[4:0] T180;
  wire[4:0] id_raddr2;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[4:0] T187;
  wire[4:0] T188;
  wire T189;
  wire T190;
  wire T191;
  wire id_fp_val;
  wire T192;
  wire[31:0] T193;
  wire T194;
  wire[31:0] T195;
  wire T196;
  wire id_sboard_hazard;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire[4:0] T201;
  wire[4:0] T202;
  wire T203;
  wire[31:0] T204;
  wire[31:0] T205;
  wire[31:0] T206;
  wire[31:0] T207;
  reg [31:0] R208;
  wire[31:0] T795;
  wire[31:0] T209;
  wire[31:0] T210;
  wire[31:0] T211;
  wire[31:0] T212;
  wire[31:0] T213;
  wire T214;
  wire wb_set_sboard;
  wire T215;
  reg  wb_reg_div_mul_val;
  wire T216;
  reg  mem_reg_div_mul_val;
  wire T217;
  reg  ex_reg_div_mul_val;
  wire T218;
  wire T219;
  wire id_div_val;
  wire[31:0] T220;
  wire id_mul_val;
  wire[31:0] T221;
  wire T222;
  wire id_wen_not0;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire[4:0] T229;
  wire[4:0] T230;
  wire T231;
  wire id_renx2_not0;
  wire T232;
  wire id_renx2;
  wire T233;
  wire[31:0] T234;
  wire T235;
  wire T236;
  wire[31:0] T237;
  wire T238;
  wire[31:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[4:0] T244;
  wire[4:0] T245;
  wire T246;
  wire id_renx1_not0;
  wire T247;
  wire id_renx1;
  wire T248;
  wire[31:0] T249;
  wire T250;
  wire T251;
  wire[31:0] T252;
  wire T253;
  wire T254;
  wire[31:0] T255;
  wire T256;
  wire T257;
  wire[31:0] T258;
  wire T259;
  wire T260;
  wire[31:0] T261;
  wire T262;
  wire[31:0] T263;
  wire T264;
  wire id_wb_hazard;
  wire T265;
  wire T266;
  reg  wb_reg_fp_val;
  wire T267;
  wire fp_data_hazard_wb;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire data_hazard_wb;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  reg  wb_reg_wen;
  wire T288;
  wire T289;
  wire id_mem_hazard;
  wire T290;
  wire fp_data_hazard_mem;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  reg  mem_mem_cmd_bh;
  wire T308;
  wire ex_slow_bypass;
  wire T309;
  wire T310;
  reg [2:0] ex_reg_mem_type;
  wire[2:0] T311;
  wire[2:0] T312;
  wire[2:0] id_mem_type;
  wire[1:0] T313;
  wire T314;
  wire[31:0] T315;
  wire T316;
  wire[31:0] T317;
  wire T318;
  wire[31:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  reg [4:0] ex_reg_mem_cmd;
  wire[4:0] T327;
  wire[4:0] id_mem_cmd;
  wire[3:0] T328;
  wire[2:0] T329;
  wire[1:0] T330;
  wire T331;
  wire T332;
  wire[31:0] T333;
  wire T334;
  wire T335;
  wire[31:0] T336;
  wire T337;
  wire[31:0] T338;
  wire T339;
  wire T340;
  wire[31:0] T341;
  wire T342;
  wire[31:0] T343;
  wire T344;
  wire T345;
  wire[31:0] T346;
  wire T347;
  wire T348;
  wire[31:0] T349;
  wire T350;
  wire[31:0] T351;
  wire T352;
  wire T353;
  reg [1:0] mem_reg_csr;
  wire[1:0] T354;
  reg [1:0] ex_reg_csr;
  wire[1:0] T355;
  wire data_hazard_mem;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire id_ex_hazard;
  wire T364;
  wire T365;
  wire fp_data_hazard_ex;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  reg  ex_reg_jalr;
  wire T383;
  wire id_jalr;
  wire[31:0] T384;
  wire T385;
  wire data_hazard_ex;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire take_pc;
  wire take_pc_mem;
  wire T395;
  reg  mem_reg_jal;
  wire T396;
  reg  ex_reg_jal;
  wire T397;
  wire id_jal;
  wire[31:0] T398;
  wire T399;
  reg  mem_reg_jalr;
  wire T400;
  reg  mem_reg_branch;
  wire T401;
  reg  ex_reg_branch;
  wire T402;
  wire id_branch;
  wire[31:0] T403;
  wire T404;
  wire ctrl_killx;
  wire T405;
  wire T406;
  reg  ex_reg_load_use;
  wire T407;
  wire id_load_use;
  wire T408;
  wire T409;
  wire replay_ex_structural;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  reg  mem_reg_sret;
  wire T415;
  reg  ex_reg_sret;
  wire T416;
  wire id_sret;
  wire[31:0] T417;
  wire ctrl_killm;
  wire T418;
  wire T419;
  wire killm_common;
  wire T420;
  reg  mem_reg_valid;
  wire T421;
  reg  ex_reg_valid;
  wire T422;
  wire T423;
  reg  mem_reg_xcpt;
  wire T424;
  wire ex_xcpt;
  wire T425;
  wire T426;
  reg  ex_reg_xcpt;
  wire T427;
  wire id_xcpt;
  wire id_syscall;
  wire[31:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire id_csr_fp;
  wire T433;
  wire[11:0] T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire id_csr_privileged;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire T445;
  wire T446;
  wire[1:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire T453;
  wire T454;
  wire[1:0] T455;
  wire T456;
  wire T457;
  wire[1:0] T458;
  wire T459;
  wire T460;
  wire id_csr_invalid;
  wire T461;
  reg  T462;
  wire T464;
  wire id_int_val;
  wire T465;
  wire[31:0] T466;
  wire T467;
  wire T468;
  wire[31:0] T469;
  wire T470;
  wire T471;
  wire[31:0] T472;
  wire T473;
  wire T474;
  wire[31:0] T475;
  wire T476;
  wire T477;
  wire[31:0] T478;
  wire T479;
  wire T480;
  wire[31:0] T481;
  wire T482;
  wire T483;
  wire[31:0] T484;
  wire T485;
  wire T486;
  wire[31:0] T487;
  wire T488;
  wire T489;
  wire[31:0] T490;
  wire T491;
  wire T492;
  wire[31:0] T493;
  wire T494;
  wire T495;
  wire[31:0] T496;
  wire T497;
  wire T498;
  wire[31:0] T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire[31:0] T504;
  wire T505;
  wire T506;
  wire[31:0] T507;
  wire T508;
  wire T509;
  wire[31:0] T510;
  wire T511;
  wire T512;
  wire[31:0] T513;
  wire T514;
  wire T515;
  wire[31:0] T516;
  wire T517;
  wire T518;
  wire T519;
  wire[31:0] T520;
  wire T521;
  wire T522;
  wire T523;
  wire[31:0] T524;
  wire T525;
  wire T526;
  wire[31:0] T527;
  wire T528;
  wire T529;
  wire[31:0] T530;
  wire T531;
  wire T532;
  wire[31:0] T533;
  wire T534;
  wire T535;
  wire[31:0] T536;
  wire T537;
  wire T538;
  wire[31:0] T539;
  wire T540;
  wire T541;
  wire[31:0] T542;
  wire T543;
  wire T544;
  wire[31:0] T545;
  wire T546;
  wire T547;
  wire[31:0] T548;
  wire T549;
  wire T550;
  wire[31:0] T551;
  wire T552;
  wire T553;
  wire[31:0] T554;
  wire T555;
  wire T556;
  wire[31:0] T557;
  wire T558;
  wire T559;
  wire[31:0] T560;
  wire T561;
  wire T562;
  wire[31:0] T563;
  wire T564;
  wire T565;
  reg  ex_reg_xcpt_interrupt;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire mem_xcpt;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  reg  mem_reg_xcpt_interrupt;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire wb_rocc_val;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  reg  wb_reg_flush_inst;
  wire T587;
  reg  mem_reg_flush_inst;
  wire T588;
  reg  ex_reg_flush_inst;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T596;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T597;
  wire T598;
  wire T599;
  reg  ex_reg_btb_hit;
  wire T600;
  reg [6:0] mem_reg_btb_resp_bht_history;
  wire[6:0] T601;
  reg [6:0] ex_reg_btb_resp_bht_history;
  wire[6:0] T602;
  reg [5:0] mem_reg_btb_resp_entry;
  wire[5:0] T603;
  reg [5:0] ex_reg_btb_resp_entry;
  wire[5:0] T604;
  reg [42:0] mem_reg_btb_resp_target;
  wire[42:0] T605;
  reg [42:0] ex_reg_btb_resp_target;
  wire[42:0] T606;
  reg  mem_reg_btb_resp_taken;
  wire T607;
  reg  ex_reg_btb_resp_taken;
  wire T608;
  reg  mem_reg_btb_hit;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  reg [63:0] wb_reg_cause;
  wire[63:0] T615;
  wire[63:0] mem_cause;
  wire[63:0] T796;
  wire[3:0] T616;
  wire[3:0] T617;
  wire[3:0] T618;
  reg [63:0] mem_reg_cause;
  wire[63:0] T619;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T620;
  wire[63:0] id_cause;
  wire[63:0] T797;
  wire[3:0] T621;
  wire[3:0] T622;
  wire[3:0] T623;
  wire[3:0] T624;
  wire[3:0] T625;
  wire[3:0] T626;
  wire[3:0] T627;
  wire[63:0] id_interrupt_cause;
  wire[63:0] T628;
  wire[63:0] T629;
  wire[63:0] T630;
  wire[63:0] T631;
  wire[63:0] T632;
  wire[63:0] T633;
  wire T634;
  wire T635;
  reg  wb_reg_valid;
  wire T636;
  wire T637;
  wire[1:0] T638;
  wire[1:0] T639;
  wire[1:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire[1:0] T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire[2:0] T798;
  reg [1:0] wb_reg_csr;
  wire[1:0] T679;
  wire T680;
  wire[3:0] T681;
  wire[3:0] id_fn_alu;
  wire[2:0] T682;
  wire[1:0] T683;
  wire T684;
  wire T685;
  wire[31:0] T686;
  wire T687;
  wire T688;
  wire[31:0] T689;
  wire T690;
  wire[31:0] T691;
  wire T692;
  wire T693;
  wire[31:0] T694;
  wire T695;
  wire T696;
  wire[31:0] T697;
  wire T698;
  wire T699;
  wire[31:0] T700;
  wire T701;
  wire T702;
  wire[31:0] T703;
  wire T704;
  wire[31:0] T705;
  wire T706;
  wire T707;
  wire[31:0] T708;
  wire T709;
  wire T710;
  wire[31:0] T711;
  wire T712;
  wire T713;
  wire[31:0] T714;
  wire T715;
  wire[31:0] T716;
  wire T717;
  wire T718;
  wire[31:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire[31:0] T723;
  wire T724;
  wire[31:0] T725;
  wire T726;
  wire id_fn_dw;
  wire T727;
  wire[31:0] T728;
  wire T729;
  wire[31:0] T730;
  wire[2:0] T731;
  wire[2:0] id_sel_imm;
  wire[1:0] T732;
  wire T733;
  wire T734;
  wire[31:0] T735;
  wire T736;
  wire[31:0] T737;
  wire T738;
  wire T739;
  wire[31:0] T740;
  wire T741;
  wire T742;
  wire[31:0] T743;
  wire T744;
  wire T745;
  wire[31:0] T746;
  wire T747;
  wire[31:0] T748;
  wire[1:0] T749;
  wire[1:0] id_sel_alu1;
  wire T750;
  wire T751;
  wire[31:0] T752;
  wire T753;
  wire T754;
  wire[31:0] T755;
  wire T756;
  wire T757;
  wire T758;
  wire[31:0] T759;
  wire T760;
  wire[31:0] T761;
  wire T762;
  wire T763;
  wire[31:0] T764;
  wire T765;
  wire[31:0] T766;
  wire[2:0] T799;
  wire[1:0] T767;
  wire[1:0] id_sel_alu2;
  wire T768;
  wire T769;
  wire[31:0] T770;
  wire T771;
  wire T772;
  wire T773;
  wire[31:0] T774;
  wire T775;
  wire T776;
  wire[31:0] T777;
  wire T778;
  wire[31:0] T779;
  wire T780;
  wire T781;
  wire[31:0] T782;
  wire T783;
  wire T784;
  wire T785;
  wire[31:0] T786;
  wire T787;
  wire T788;
  wire T789;
  wire[2:0] T800;
  wire[1:0] T790;
  wire[1:0] T791;
  wire[1:0] T792;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_xcpt = {1{$random}};
    wb_reg_sret = {1{$random}};
    mem_reg_replay = {1{$random}};
    mem_reg_replay_next = {1{$random}};
    ex_reg_replay_next = {1{$random}};
    id_reg_fence = {1{$random}};
    ex_reg_mem_val = {1{$random}};
    R105 = {1{$random}};
    wb_reg_rocc_val = {1{$random}};
    mem_reg_rocc_val = {1{$random}};
    ex_reg_rocc_val = {1{$random}};
    wb_reg_replay = {1{$random}};
    mem_reg_fp_val = {1{$random}};
    ex_reg_fp_val = {1{$random}};
    mem_reg_wen = {1{$random}};
    ex_reg_wen = {1{$random}};
    wb_reg_fp_wen = {1{$random}};
    mem_reg_fp_wen = {1{$random}};
    ex_reg_fp_wen = {1{$random}};
    wb_reg_mem_val = {1{$random}};
    mem_reg_mem_val = {1{$random}};
    R208 = {1{$random}};
    wb_reg_div_mul_val = {1{$random}};
    mem_reg_div_mul_val = {1{$random}};
    ex_reg_div_mul_val = {1{$random}};
    wb_reg_fp_val = {1{$random}};
    wb_reg_wen = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_reg_mem_type = {1{$random}};
    ex_reg_mem_cmd = {1{$random}};
    mem_reg_csr = {1{$random}};
    ex_reg_csr = {1{$random}};
    ex_reg_jalr = {1{$random}};
    mem_reg_jal = {1{$random}};
    ex_reg_jal = {1{$random}};
    mem_reg_jalr = {1{$random}};
    mem_reg_branch = {1{$random}};
    ex_reg_branch = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_reg_sret = {1{$random}};
    ex_reg_sret = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    wb_reg_flush_inst = {1{$random}};
    mem_reg_flush_inst = {1{$random}};
    ex_reg_flush_inst = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_valid = {1{$random}};
    wb_reg_csr = {1{$random}};
  end
`endif

  assign io_rocc_exception = T0;
  assign T0 = wb_reg_xcpt & io_dpath_status_er;
  assign T1 = mem_xcpt & T2;
  assign T2 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T3;
  assign T3 = T570 | wb_reg_sret;
  assign T4 = ctrl_killm ? 1'h0 : T5;
  assign T5 = mem_reg_sret & T6;
  assign T6 = mem_reg_replay ^ 1'h1;
  assign T7 = T414 & replay_ex;
  assign replay_ex = replay_ex_structural | replay_ex_other;
  assign replay_ex_other = T406 | mem_reg_replay_next;
  assign T8 = ctrl_killx ? 1'h0 : ex_reg_replay_next;
  assign T9 = ctrl_killd ? 1'h0 : T10;
  assign T10 = id_replay_next | id_csr_flush;
  assign id_csr_flush = T17 & T11;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T15 | T13;
  assign T13 = T14 == 12'h400;
  assign T14 = id_csr_addr & 12'hc2d;
  assign id_csr_addr = io_dpath_inst[5'h1f:5'h14];
  assign T15 = T16 == 12'h400;
  assign T16 = id_csr_addr & 12'hc2e;
  assign T17 = id_csr_en & id_csr_wen;
  assign id_csr_wen = T26 | T18;
  assign T18 = T19 ^ 1'h1;
  assign T19 = T25 | T20;
  assign T20 = 2'h3 == id_csr;
  assign id_csr = {T23, T21};
  assign T21 = T22 == 32'h1070;
  assign T22 = io_dpath_inst & 32'h1070;
  assign T23 = T24 == 32'h2070;
  assign T24 = io_dpath_inst & 32'h2070;
  assign T25 = 2'h2 == id_csr;
  assign T26 = id_raddr1 != 5'h0;
  assign id_raddr1 = io_dpath_inst[5'h13:4'hf];
  assign id_csr_en = id_csr != 2'h0;
  assign id_replay_next = T27 == 32'h1008;
  assign T27 = io_dpath_inst & 32'h3058;
  assign ctrl_killd = T28;
  assign T28 = T59 | ctrl_draind;
  assign ctrl_draind = id_interrupt | ex_reg_replay_next;
  assign id_interrupt = io_dpath_status_ei & id_interrupt_unmasked;
  assign id_interrupt_unmasked = T32 | T29;
  assign T29 = T31 & T30;
  assign T30 = io_dpath_status_ip[3'h7:3'h7];
  assign T31 = io_dpath_status_im[3'h7:3'h7];
  assign T32 = T36 | T33;
  assign T33 = T35 & T34;
  assign T34 = io_dpath_status_ip[3'h6:3'h6];
  assign T35 = io_dpath_status_im[3'h6:3'h6];
  assign T36 = T40 | T37;
  assign T37 = T39 & T38;
  assign T38 = io_dpath_status_ip[3'h5:3'h5];
  assign T39 = io_dpath_status_im[3'h5:3'h5];
  assign T40 = T44 | T41;
  assign T41 = T43 & T42;
  assign T42 = io_dpath_status_ip[3'h4:3'h4];
  assign T43 = io_dpath_status_im[3'h4:3'h4];
  assign T44 = T48 | T45;
  assign T45 = T47 & T46;
  assign T46 = io_dpath_status_ip[2'h3:2'h3];
  assign T47 = io_dpath_status_im[2'h3:2'h3];
  assign T48 = T52 | T49;
  assign T49 = T51 & T50;
  assign T50 = io_dpath_status_ip[2'h2:2'h2];
  assign T51 = io_dpath_status_im[2'h2:2'h2];
  assign T52 = T56 | T53;
  assign T53 = T55 & T54;
  assign T54 = io_dpath_status_ip[1'h1:1'h1];
  assign T55 = io_dpath_status_im[1'h1:1'h1];
  assign T56 = T58 & T57;
  assign T57 = io_dpath_status_ip[1'h0:1'h0];
  assign T58 = io_dpath_status_im[1'h0:1'h0];
  assign T59 = T394 | ctrl_stalld;
  assign ctrl_stalld = T93 | id_do_fence;
  assign id_do_fence = id_mem_busy & T60;
  assign T60 = T61 | id_csr_flush;
  assign T61 = T87 | T62;
  assign T62 = id_reg_fence & id_mem_val;
  assign id_mem_val = T65 | T63;
  assign T63 = T64 == 32'h1000202f;
  assign T64 = io_dpath_inst & 32'hf9f0607f;
  assign T65 = T68 | T66;
  assign T66 = T67 == 32'h800202f;
  assign T67 = io_dpath_inst & 32'he800607f;
  assign T68 = T71 | T69;
  assign T69 = T70 == 32'h202f;
  assign T70 = io_dpath_inst & 32'h1800607f;
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h2003;
  assign T73 = io_dpath_inst & 32'h605b;
  assign T74 = T77 | T75;
  assign T75 = T76 == 32'h3;
  assign T76 = io_dpath_inst & 32'h107f;
  assign T77 = T80 | T78;
  assign T78 = T79 == 32'h3;
  assign T79 = io_dpath_inst & 32'h207f;
  assign T80 = T81 == 32'h3;
  assign T81 = io_dpath_inst & 32'h405f;
  assign T793 = reset ? 1'h0 : T82;
  assign T82 = id_fence_next | T83;
  assign T83 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_fence | T84;
  assign T84 = id_amo & id_amo_rl;
  assign id_amo_rl = io_dpath_inst[5'h19:5'h19];
  assign id_amo = T85 == 32'h2008;
  assign T85 = io_dpath_inst & 32'h6048;
  assign id_fence = T86 == 32'h8;
  assign T86 = io_dpath_inst & 32'h3058;
  assign T87 = T89 | id_fence_i;
  assign id_fence_i = T88 == 32'h100f;
  assign T88 = io_dpath_inst & 32'h707f;
  assign T89 = id_amo & id_amo_aq;
  assign id_amo_aq = io_dpath_inst[5'h1a:5'h1a];
  assign id_mem_busy = T92 | ex_reg_mem_val;
  assign T90 = ctrl_killd ? 1'h0 : T91;
  assign T91 = id_mem_val;
  assign T92 = io_dmem_ordered ^ 1'h1;
  assign T93 = T96 | T94;
  assign T94 = id_mem_val & T95;
  assign T95 = io_dmem_req_ready ^ 1'h1;
  assign T96 = T196 | T97;
  assign T97 = id_fp_val & id_stall_fpu;
  assign id_stall_fpu = T166 | T98;
  assign T98 = io_fpu_dec_wen & T99;
  assign T99 = T104 & T100;
  assign T100 = T101 - 1'h1;
  assign T101 = 1'h1 << T102;
  assign T102 = T103 + 5'h1;
  assign T103 = id_waddr - id_waddr;
  assign id_waddr = io_dpath_inst[4'hb:3'h7];
  assign T104 = R105 >> id_waddr;
  assign T794 = reset ? 32'h0 : T106;
  assign T106 = T165 ? T161 : T107;
  assign T107 = T160 ? T156 : T108;
  assign T108 = T112 ? T109 : R105;
  assign T109 = R105 | T110;
  assign T110 = T112 ? T111 : 32'h0;
  assign T111 = 1'h1 << io_dpath_wb_waddr;
  assign T112 = T147 & T113;
  assign T113 = replay_wb ^ 1'h1;
  assign replay_wb = replay_wb_common | T114;
  assign T114 = wb_reg_rocc_val & T115;
  assign T115 = io_rocc_cmd_ready ^ 1'h1;
  assign T116 = ctrl_killm ? 1'h0 : mem_reg_rocc_val;
  assign T117 = ctrl_killx ? 1'h0 : ex_reg_rocc_val;
  assign T118 = ctrl_killd ? 1'h0 : T119;
  assign T119 = 1'h0;
  assign replay_wb_common = T120 | io_dpath_csr_replay;
  assign T120 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T121 = replay_mem & T122;
  assign T122 = take_pc_wb ^ 1'h1;
  assign replay_mem = T125 | fpu_kill_mem;
  assign fpu_kill_mem = mem_reg_fp_val & io_fpu_nack_mem;
  assign T123 = ctrl_killx ? 1'h0 : ex_reg_fp_val;
  assign T124 = ctrl_killd ? 1'h0 : id_fp_val;
  assign T125 = dcache_kill_mem | mem_reg_replay;
  assign dcache_kill_mem = mem_reg_wen & io_dmem_replay_next_valid;
  assign T126 = ctrl_killx ? 1'h0 : ex_reg_wen;
  assign T127 = ctrl_killd ? 1'h0 : id_wen;
  assign id_wen = T130 | T128;
  assign T128 = T129 == 32'h80000010;
  assign T129 = io_dpath_inst & 32'h90000030;
  assign T130 = T133 | T131;
  assign T131 = T132 == 32'h2030;
  assign T132 = io_dpath_inst & 32'h2030;
  assign T133 = T136 | T134;
  assign T134 = T135 == 32'h1030;
  assign T135 = io_dpath_inst & 32'h1030;
  assign T136 = T139 | T137;
  assign T137 = T138 == 32'h28;
  assign T138 = io_dpath_inst & 32'h28;
  assign T139 = T142 | T140;
  assign T140 = T141 == 32'h24;
  assign T141 = io_dpath_inst & 32'h2024;
  assign T142 = T145 | T143;
  assign T143 = T144 == 32'h10;
  assign T144 = io_dpath_inst & 32'h50;
  assign T145 = T146 == 32'h0;
  assign T146 = io_dpath_inst & 32'h64;
  assign T147 = T148 | io_fpu_sboard_set;
  assign T148 = wb_dcache_miss & wb_reg_fp_wen;
  assign T149 = ctrl_killm ? 1'h0 : mem_reg_fp_wen;
  assign T150 = ctrl_killx ? 1'h0 : ex_reg_fp_wen;
  assign T151 = ctrl_killd ? 1'h0 : T152;
  assign T152 = id_fp_val & io_fpu_dec_wen;
  assign wb_dcache_miss = wb_reg_mem_val & T153;
  assign T153 = io_dmem_resp_valid ^ 1'h1;
  assign T154 = ctrl_killm ? 1'h0 : mem_reg_mem_val;
  assign T155 = ctrl_killx ? 1'h0 : ex_reg_mem_val;
  assign T156 = T109 & T157;
  assign T157 = ~ T158;
  assign T158 = io_dpath_fp_sboard_clr ? T159 : 32'h0;
  assign T159 = 1'h1 << io_dpath_fp_sboard_clra;
  assign T160 = T112 | io_dpath_fp_sboard_clr;
  assign T161 = T156 & T162;
  assign T162 = ~ T163;
  assign T163 = io_fpu_sboard_clr ? T164 : 32'h0;
  assign T164 = 1'h1 << io_fpu_sboard_clra;
  assign T165 = T160 | io_fpu_sboard_clr;
  assign T166 = T174 | T167;
  assign T167 = io_fpu_dec_ren3 & T168;
  assign T168 = T173 & T169;
  assign T169 = T170 - 1'h1;
  assign T170 = 1'h1 << T171;
  assign T171 = T172 + 5'h1;
  assign T172 = id_raddr3 - id_raddr3;
  assign id_raddr3 = io_dpath_inst[5'h1f:5'h1b];
  assign T173 = R105 >> id_raddr3;
  assign T174 = T182 | T175;
  assign T175 = io_fpu_dec_ren2 & T176;
  assign T176 = T181 & T177;
  assign T177 = T178 - 1'h1;
  assign T178 = 1'h1 << T179;
  assign T179 = T180 + 5'h1;
  assign T180 = id_raddr2 - id_raddr2;
  assign id_raddr2 = io_dpath_inst[5'h18:5'h14];
  assign T181 = R105 >> id_raddr2;
  assign T182 = T190 | T183;
  assign T183 = io_fpu_dec_ren1 & T184;
  assign T184 = T189 & T185;
  assign T185 = T186 - 1'h1;
  assign T186 = 1'h1 << T187;
  assign T187 = T188 + 5'h1;
  assign T188 = id_raddr1 - id_raddr1;
  assign T189 = R105 >> id_raddr1;
  assign T190 = id_csr_en & T191;
  assign T191 = io_fpu_fcsr_rdy ^ 1'h1;
  assign id_fp_val = T194 | T192;
  assign T192 = T193 == 32'h40;
  assign T193 = io_dpath_inst & 32'h60;
  assign T194 = T195 == 32'h4;
  assign T195 = io_dpath_inst & 32'h5c;
  assign T196 = T264 | id_sboard_hazard;
  assign id_sboard_hazard = T224 | T197;
  assign T197 = id_wen_not0 & T198;
  assign T198 = T203 & T199;
  assign T199 = T200 - 1'h1;
  assign T200 = 1'h1 << T201;
  assign T201 = T202 + 5'h1;
  assign T202 = id_waddr - id_waddr;
  assign T203 = T204 >> id_waddr;
  assign T204 = R208 & T205;
  assign T205 = ~ T206;
  assign T206 = io_dpath_ll_wen ? T207 : 32'h0;
  assign T207 = 1'h1 << io_dpath_ll_waddr;
  assign T795 = reset ? 32'h0 : T209;
  assign T209 = T222 ? T211 : T210;
  assign T210 = io_dpath_ll_wen ? T204 : R208;
  assign T211 = T204 | T212;
  assign T212 = T214 ? T213 : 32'h0;
  assign T213 = 1'h1 << io_dpath_wb_waddr;
  assign T214 = wb_set_sboard & io_dpath_wb_wen;
  assign wb_set_sboard = T215 | wb_reg_rocc_val;
  assign T215 = wb_reg_div_mul_val | wb_dcache_miss;
  assign T216 = ctrl_killm ? 1'h0 : mem_reg_div_mul_val;
  assign T217 = ex_reg_div_mul_val & io_dpath_div_mul_rdy;
  assign T218 = ctrl_killd ? 1'h0 : T219;
  assign T219 = id_mul_val | id_div_val;
  assign id_div_val = T220 == 32'h2004020;
  assign T220 = io_dpath_inst & 32'h2004064;
  assign id_mul_val = T221 == 32'h2000030;
  assign T221 = io_dpath_inst & 32'h2004074;
  assign T222 = io_dpath_ll_wen | T214;
  assign id_wen_not0 = id_wen & T223;
  assign T223 = id_waddr != 5'h0;
  assign T224 = T240 | T225;
  assign T225 = id_renx2_not0 & T226;
  assign T226 = T231 & T227;
  assign T227 = T228 - 1'h1;
  assign T228 = 1'h1 << T229;
  assign T229 = T230 + 5'h1;
  assign T230 = id_raddr2 - id_raddr2;
  assign T231 = T204 >> id_raddr2;
  assign id_renx2_not0 = id_renx2 & T232;
  assign T232 = id_raddr2 != 5'h0;
  assign id_renx2 = T235 | T233;
  assign T233 = T234 == 32'h2008;
  assign T234 = io_dpath_inst & 32'h2048;
  assign T235 = T238 | T236;
  assign T236 = T237 == 32'h20;
  assign T237 = io_dpath_inst & 32'h34;
  assign T238 = T239 == 32'h20;
  assign T239 = io_dpath_inst & 32'h64;
  assign T240 = id_renx1_not0 & T241;
  assign T241 = T246 & T242;
  assign T242 = T243 - 1'h1;
  assign T243 = 1'h1 << T244;
  assign T244 = T245 + 5'h1;
  assign T245 = id_raddr1 - id_raddr1;
  assign T246 = T204 >> id_raddr1;
  assign id_renx1_not0 = id_renx1 & T247;
  assign T247 = id_raddr1 != 5'h0;
  assign id_renx1 = T250 | T248;
  assign T248 = T249 == 32'h90000010;
  assign T249 = io_dpath_inst & 32'h90000034;
  assign T250 = T253 | T251;
  assign T251 = T252 == 32'h2020;
  assign T252 = io_dpath_inst & 32'h6024;
  assign T253 = T256 | T254;
  assign T254 = T255 == 32'h2000;
  assign T255 = io_dpath_inst & 32'h2050;
  assign T256 = T259 | T257;
  assign T257 = T258 == 32'h1020;
  assign T258 = io_dpath_inst & 32'h5024;
  assign T259 = T262 | T260;
  assign T260 = T261 == 32'h20;
  assign T261 = io_dpath_inst & 32'h38;
  assign T262 = T263 == 32'h0;
  assign T263 = io_dpath_inst & 32'h44;
  assign T264 = T289 | id_wb_hazard;
  assign id_wb_hazard = T279 | T265;
  assign T265 = fp_data_hazard_wb & T266;
  assign T266 = wb_dcache_miss | wb_reg_fp_val;
  assign T267 = ctrl_killm ? 1'h0 : mem_reg_fp_val;
  assign fp_data_hazard_wb = wb_reg_fp_wen & T268;
  assign T268 = T271 | T269;
  assign T269 = io_fpu_dec_wen & T270;
  assign T270 = id_waddr == io_dpath_wb_waddr;
  assign T271 = T274 | T272;
  assign T272 = io_fpu_dec_ren3 & T273;
  assign T273 = id_raddr3 == io_dpath_wb_waddr;
  assign T274 = T277 | T275;
  assign T275 = io_fpu_dec_ren2 & T276;
  assign T276 = id_raddr2 == io_dpath_wb_waddr;
  assign T277 = io_fpu_dec_ren1 & T278;
  assign T278 = id_raddr1 == io_dpath_wb_waddr;
  assign T279 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_reg_wen & T280;
  assign T280 = T283 | T281;
  assign T281 = id_wen_not0 & T282;
  assign T282 = id_waddr == io_dpath_wb_waddr;
  assign T283 = T286 | T284;
  assign T284 = id_renx2_not0 & T285;
  assign T285 = id_raddr2 == io_dpath_wb_waddr;
  assign T286 = id_renx1_not0 & T287;
  assign T287 = id_raddr1 == io_dpath_wb_waddr;
  assign T288 = ctrl_killm ? 1'h0 : mem_reg_wen;
  assign T289 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = T302 | T290;
  assign T290 = fp_data_hazard_mem & mem_reg_fp_val;
  assign fp_data_hazard_mem = mem_reg_fp_wen & T291;
  assign T291 = T294 | T292;
  assign T292 = io_fpu_dec_wen & T293;
  assign T293 = id_waddr == io_dpath_mem_waddr;
  assign T294 = T297 | T295;
  assign T295 = io_fpu_dec_ren3 & T296;
  assign T296 = id_raddr3 == io_dpath_mem_waddr;
  assign T297 = T300 | T298;
  assign T298 = io_fpu_dec_ren2 & T299;
  assign T299 = id_raddr2 == io_dpath_mem_waddr;
  assign T300 = io_fpu_dec_ren1 & T301;
  assign T301 = id_raddr1 == io_dpath_mem_waddr;
  assign T302 = data_hazard_mem & T303;
  assign T303 = T304 | mem_reg_rocc_val;
  assign T304 = T305 | mem_reg_fp_val;
  assign T305 = T306 | mem_reg_div_mul_val;
  assign T306 = T353 | T307;
  assign T307 = mem_reg_mem_val & mem_mem_cmd_bh;
  assign T308 = T352 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T326 | T309;
  assign T309 = T321 | T310;
  assign T310 = 3'h5 == ex_reg_mem_type;
  assign T311 = T320 ? T312 : ex_reg_mem_type;
  assign T312 = id_mem_type;
  assign id_mem_type = {T318, T313};
  assign T313 = {T316, T314};
  assign T314 = T315 == 32'h1000;
  assign T315 = io_dpath_inst & 32'h1000;
  assign T316 = T317 == 32'h2000;
  assign T317 = io_dpath_inst & 32'h2000;
  assign T318 = T319 == 32'h4000;
  assign T319 = io_dpath_inst & 32'h4000;
  assign T320 = ctrl_killd ^ 1'h1;
  assign T321 = T323 | T322;
  assign T322 = 3'h1 == ex_reg_mem_type;
  assign T323 = T325 | T324;
  assign T324 = 3'h4 == ex_reg_mem_type;
  assign T325 = 3'h0 == ex_reg_mem_type;
  assign T326 = ex_reg_mem_cmd == 5'h7;
  assign T327 = T320 ? id_mem_cmd : ex_reg_mem_cmd;
  assign id_mem_cmd = {1'h0, T328};
  assign T328 = {T350, T329};
  assign T329 = {T344, T330};
  assign T330 = {T339, T331};
  assign T331 = T334 | T332;
  assign T332 = T333 == 32'h20000020;
  assign T333 = io_dpath_inst & 32'h20000020;
  assign T334 = T337 | T335;
  assign T335 = T336 == 32'h18000020;
  assign T336 = io_dpath_inst & 32'h18000020;
  assign T337 = T338 == 32'h20;
  assign T338 = io_dpath_inst & 32'h28;
  assign T339 = T342 | T340;
  assign T340 = T341 == 32'h40000008;
  assign T341 = io_dpath_inst & 32'h40000008;
  assign T342 = T343 == 32'h10000008;
  assign T343 = io_dpath_inst & 32'h10000008;
  assign T344 = T347 | T345;
  assign T345 = T346 == 32'h80000008;
  assign T346 = io_dpath_inst & 32'h80000008;
  assign T347 = T348 | T342;
  assign T348 = T349 == 32'h8000008;
  assign T349 = io_dpath_inst & 32'h8000008;
  assign T350 = T351 == 32'h8;
  assign T351 = io_dpath_inst & 32'h18000008;
  assign T352 = ctrl_killx ^ 1'h1;
  assign T353 = mem_reg_csr != 2'h0;
  assign T354 = ctrl_killx ? 2'h0 : ex_reg_csr;
  assign T355 = ctrl_killd ? 2'h0 : id_csr;
  assign data_hazard_mem = mem_reg_wen & T356;
  assign T356 = T359 | T357;
  assign T357 = id_wen_not0 & T358;
  assign T358 = id_waddr == io_dpath_mem_waddr;
  assign T359 = T362 | T360;
  assign T360 = id_renx2_not0 & T361;
  assign T361 = id_raddr2 == io_dpath_mem_waddr;
  assign T362 = id_renx1_not0 & T363;
  assign T363 = id_raddr1 == io_dpath_mem_waddr;
  assign id_ex_hazard = T377 | T364;
  assign T364 = fp_data_hazard_ex & T365;
  assign T365 = ex_reg_mem_val | ex_reg_fp_val;
  assign fp_data_hazard_ex = ex_reg_fp_wen & T366;
  assign T366 = T369 | T367;
  assign T367 = io_fpu_dec_wen & T368;
  assign T368 = id_waddr == io_dpath_ex_waddr;
  assign T369 = T372 | T370;
  assign T370 = io_fpu_dec_ren3 & T371;
  assign T371 = id_raddr3 == io_dpath_ex_waddr;
  assign T372 = T375 | T373;
  assign T373 = io_fpu_dec_ren2 & T374;
  assign T374 = id_raddr2 == io_dpath_ex_waddr;
  assign T375 = io_fpu_dec_ren1 & T376;
  assign T376 = id_raddr1 == io_dpath_ex_waddr;
  assign T377 = data_hazard_ex & T378;
  assign T378 = T379 | ex_reg_rocc_val;
  assign T379 = T380 | ex_reg_fp_val;
  assign T380 = T381 | ex_reg_div_mul_val;
  assign T381 = T382 | ex_reg_mem_val;
  assign T382 = T385 | ex_reg_jalr;
  assign T383 = ctrl_killd ? 1'h0 : id_jalr;
  assign id_jalr = T384 == 32'h24;
  assign T384 = io_dpath_inst & 32'h203c;
  assign T385 = ex_reg_csr != 2'h0;
  assign data_hazard_ex = ex_reg_wen & T386;
  assign T386 = T389 | T387;
  assign T387 = id_wen_not0 & T388;
  assign T388 = id_waddr == io_dpath_ex_waddr;
  assign T389 = T392 | T390;
  assign T390 = id_renx2_not0 & T391;
  assign T391 = id_raddr2 == io_dpath_ex_waddr;
  assign T392 = id_renx1_not0 & T393;
  assign T393 = id_raddr1 == io_dpath_ex_waddr;
  assign T394 = T404 | take_pc;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = io_dpath_mem_misprediction & T395;
  assign T395 = T399 | mem_reg_jal;
  assign T396 = ctrl_killx ? 1'h0 : ex_reg_jal;
  assign T397 = ctrl_killd ? 1'h0 : id_jal;
  assign id_jal = T398 == 32'h68;
  assign T398 = io_dpath_inst & 32'h68;
  assign T399 = mem_reg_branch | mem_reg_jalr;
  assign T400 = ctrl_killx ? 1'h0 : ex_reg_jalr;
  assign T401 = ctrl_killx ? 1'h0 : ex_reg_branch;
  assign T402 = ctrl_killd ? 1'h0 : id_branch;
  assign id_branch = T403 == 32'h60;
  assign T403 = io_dpath_inst & 32'h74;
  assign T404 = io_imem_resp_valid ^ 1'h1;
  assign ctrl_killx = T405;
  assign T405 = take_pc | replay_ex;
  assign T406 = wb_dcache_miss & ex_reg_load_use;
  assign T407 = ctrl_killd ? 1'h0 : id_load_use;
  assign id_load_use = T408;
  assign T408 = mem_reg_mem_val & T409;
  assign T409 = data_hazard_mem | fp_data_hazard_mem;
  assign replay_ex_structural = T412 | T410;
  assign T410 = ex_reg_div_mul_val & T411;
  assign T411 = io_dpath_div_mul_rdy ^ 1'h1;
  assign T412 = ex_reg_mem_val & T413;
  assign T413 = io_dmem_req_ready ^ 1'h1;
  assign T414 = take_pc ^ 1'h1;
  assign T415 = ctrl_killx ? 1'h0 : ex_reg_sret;
  assign T416 = ctrl_killd ? 1'h0 : id_sret;
  assign id_sret = T417 == 32'h80000050;
  assign T417 = io_dpath_inst & 32'he0003050;
  assign ctrl_killm = T418;
  assign T418 = T419 | fpu_kill_mem;
  assign T419 = killm_common | mem_xcpt;
  assign killm_common = T423 | T420;
  assign T420 = mem_reg_valid ^ 1'h1;
  assign T421 = ctrl_killx ? 1'h0 : ex_reg_valid;
  assign T422 = ctrl_killd ? 1'h0 : 1'h1;
  assign T423 = T569 | mem_reg_xcpt;
  assign T424 = ctrl_killx ? 1'h0 : ex_xcpt;
  assign ex_xcpt = T426 | T425;
  assign T425 = ex_reg_fp_val & io_fpu_illegal_rm;
  assign T426 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T427 = ctrl_killd ? 1'h0 : id_xcpt;
  assign id_xcpt = T429 | id_syscall;
  assign id_syscall = T428 == 32'h70;
  assign T428 = io_dpath_inst & 32'h80003070;
  assign T429 = T435 | T430;
  assign T430 = T432 & T431;
  assign T431 = io_dpath_status_ef ^ 1'h1;
  assign T432 = id_fp_val | id_csr_fp;
  assign id_csr_fp = id_csr_en & T433;
  assign T433 = T434 == 12'h0;
  assign T434 = id_csr_addr & 12'h480;
  assign T435 = T438 | T436;
  assign T436 = id_sret & T437;
  assign T437 = io_dpath_status_s ^ 1'h1;
  assign T438 = T459 | id_csr_privileged;
  assign id_csr_privileged = id_csr_en & T439;
  assign T439 = T445 | T440;
  assign T440 = T441 & id_csr_wen;
  assign T441 = T443 & T442;
  assign T442 = io_dpath_status_s ^ 1'h1;
  assign T443 = T444 == 2'h1;
  assign T444 = id_csr_addr[4'h9:4'h8];
  assign T445 = T448 | T446;
  assign T446 = 2'h2 <= T447;
  assign T447 = id_csr_addr[4'h9:4'h8];
  assign T448 = T453 | T449;
  assign T449 = T451 & T450;
  assign T450 = io_dpath_status_s ^ 1'h1;
  assign T451 = T452 == 2'h1;
  assign T452 = id_csr_addr[4'hb:4'ha];
  assign T453 = T456 | T454;
  assign T454 = T455 == 2'h2;
  assign T455 = id_csr_addr[4'hb:4'ha];
  assign T456 = T457 & id_csr_wen;
  assign T457 = T458 == 2'h3;
  assign T458 = id_csr_addr[4'hb:4'ha];
  assign T459 = T564 | T460;
  assign T460 = T464 | id_csr_invalid;
  assign id_csr_invalid = id_csr_en & T461;
  assign T461 = T462 ^ 1'h1;
  always @(*) case (id_csr_addr)
    0: T462 = 1'h0;
    1: T462 = 1'h1;
    2: T462 = 1'h1;
    3: T462 = 1'h1;
    4: T462 = 1'h0;
    5: T462 = 1'h0;
    6: T462 = 1'h0;
    7: T462 = 1'h0;
    8: T462 = 1'h0;
    9: T462 = 1'h0;
    10: T462 = 1'h0;
    11: T462 = 1'h0;
    12: T462 = 1'h0;
    13: T462 = 1'h0;
    14: T462 = 1'h0;
    15: T462 = 1'h0;
    16: T462 = 1'h0;
    17: T462 = 1'h0;
    18: T462 = 1'h0;
    19: T462 = 1'h0;
    20: T462 = 1'h0;
    21: T462 = 1'h0;
    22: T462 = 1'h0;
    23: T462 = 1'h0;
    24: T462 = 1'h0;
    25: T462 = 1'h0;
    26: T462 = 1'h0;
    27: T462 = 1'h0;
    28: T462 = 1'h0;
    29: T462 = 1'h0;
    30: T462 = 1'h0;
    31: T462 = 1'h0;
    32: T462 = 1'h0;
    33: T462 = 1'h0;
    34: T462 = 1'h0;
    35: T462 = 1'h0;
    36: T462 = 1'h0;
    37: T462 = 1'h0;
    38: T462 = 1'h0;
    39: T462 = 1'h0;
    40: T462 = 1'h0;
    41: T462 = 1'h0;
    42: T462 = 1'h0;
    43: T462 = 1'h0;
    44: T462 = 1'h0;
    45: T462 = 1'h0;
    46: T462 = 1'h0;
    47: T462 = 1'h0;
    48: T462 = 1'h0;
    49: T462 = 1'h0;
    50: T462 = 1'h0;
    51: T462 = 1'h0;
    52: T462 = 1'h0;
    53: T462 = 1'h0;
    54: T462 = 1'h0;
    55: T462 = 1'h0;
    56: T462 = 1'h0;
    57: T462 = 1'h0;
    58: T462 = 1'h0;
    59: T462 = 1'h0;
    60: T462 = 1'h0;
    61: T462 = 1'h0;
    62: T462 = 1'h0;
    63: T462 = 1'h0;
    64: T462 = 1'h0;
    65: T462 = 1'h0;
    66: T462 = 1'h0;
    67: T462 = 1'h0;
    68: T462 = 1'h0;
    69: T462 = 1'h0;
    70: T462 = 1'h0;
    71: T462 = 1'h0;
    72: T462 = 1'h0;
    73: T462 = 1'h0;
    74: T462 = 1'h0;
    75: T462 = 1'h0;
    76: T462 = 1'h0;
    77: T462 = 1'h0;
    78: T462 = 1'h0;
    79: T462 = 1'h0;
    80: T462 = 1'h0;
    81: T462 = 1'h0;
    82: T462 = 1'h0;
    83: T462 = 1'h0;
    84: T462 = 1'h0;
    85: T462 = 1'h0;
    86: T462 = 1'h0;
    87: T462 = 1'h0;
    88: T462 = 1'h0;
    89: T462 = 1'h0;
    90: T462 = 1'h0;
    91: T462 = 1'h0;
    92: T462 = 1'h0;
    93: T462 = 1'h0;
    94: T462 = 1'h0;
    95: T462 = 1'h0;
    96: T462 = 1'h0;
    97: T462 = 1'h0;
    98: T462 = 1'h0;
    99: T462 = 1'h0;
    100: T462 = 1'h0;
    101: T462 = 1'h0;
    102: T462 = 1'h0;
    103: T462 = 1'h0;
    104: T462 = 1'h0;
    105: T462 = 1'h0;
    106: T462 = 1'h0;
    107: T462 = 1'h0;
    108: T462 = 1'h0;
    109: T462 = 1'h0;
    110: T462 = 1'h0;
    111: T462 = 1'h0;
    112: T462 = 1'h0;
    113: T462 = 1'h0;
    114: T462 = 1'h0;
    115: T462 = 1'h0;
    116: T462 = 1'h0;
    117: T462 = 1'h0;
    118: T462 = 1'h0;
    119: T462 = 1'h0;
    120: T462 = 1'h0;
    121: T462 = 1'h0;
    122: T462 = 1'h0;
    123: T462 = 1'h0;
    124: T462 = 1'h0;
    125: T462 = 1'h0;
    126: T462 = 1'h0;
    127: T462 = 1'h0;
    128: T462 = 1'h0;
    129: T462 = 1'h0;
    130: T462 = 1'h0;
    131: T462 = 1'h0;
    132: T462 = 1'h0;
    133: T462 = 1'h0;
    134: T462 = 1'h0;
    135: T462 = 1'h0;
    136: T462 = 1'h0;
    137: T462 = 1'h0;
    138: T462 = 1'h0;
    139: T462 = 1'h0;
    140: T462 = 1'h0;
    141: T462 = 1'h0;
    142: T462 = 1'h0;
    143: T462 = 1'h0;
    144: T462 = 1'h0;
    145: T462 = 1'h0;
    146: T462 = 1'h0;
    147: T462 = 1'h0;
    148: T462 = 1'h0;
    149: T462 = 1'h0;
    150: T462 = 1'h0;
    151: T462 = 1'h0;
    152: T462 = 1'h0;
    153: T462 = 1'h0;
    154: T462 = 1'h0;
    155: T462 = 1'h0;
    156: T462 = 1'h0;
    157: T462 = 1'h0;
    158: T462 = 1'h0;
    159: T462 = 1'h0;
    160: T462 = 1'h0;
    161: T462 = 1'h0;
    162: T462 = 1'h0;
    163: T462 = 1'h0;
    164: T462 = 1'h0;
    165: T462 = 1'h0;
    166: T462 = 1'h0;
    167: T462 = 1'h0;
    168: T462 = 1'h0;
    169: T462 = 1'h0;
    170: T462 = 1'h0;
    171: T462 = 1'h0;
    172: T462 = 1'h0;
    173: T462 = 1'h0;
    174: T462 = 1'h0;
    175: T462 = 1'h0;
    176: T462 = 1'h0;
    177: T462 = 1'h0;
    178: T462 = 1'h0;
    179: T462 = 1'h0;
    180: T462 = 1'h0;
    181: T462 = 1'h0;
    182: T462 = 1'h0;
    183: T462 = 1'h0;
    184: T462 = 1'h0;
    185: T462 = 1'h0;
    186: T462 = 1'h0;
    187: T462 = 1'h0;
    188: T462 = 1'h0;
    189: T462 = 1'h0;
    190: T462 = 1'h0;
    191: T462 = 1'h0;
    192: T462 = 1'h1;
    193: T462 = 1'h0;
    194: T462 = 1'h0;
    195: T462 = 1'h0;
    196: T462 = 1'h0;
    197: T462 = 1'h0;
    198: T462 = 1'h0;
    199: T462 = 1'h0;
    200: T462 = 1'h0;
    201: T462 = 1'h0;
    202: T462 = 1'h0;
    203: T462 = 1'h0;
    204: T462 = 1'h0;
    205: T462 = 1'h0;
    206: T462 = 1'h0;
    207: T462 = 1'h0;
    208: T462 = 1'h0;
    209: T462 = 1'h0;
    210: T462 = 1'h0;
    211: T462 = 1'h0;
    212: T462 = 1'h0;
    213: T462 = 1'h0;
    214: T462 = 1'h0;
    215: T462 = 1'h0;
    216: T462 = 1'h0;
    217: T462 = 1'h0;
    218: T462 = 1'h0;
    219: T462 = 1'h0;
    220: T462 = 1'h0;
    221: T462 = 1'h0;
    222: T462 = 1'h0;
    223: T462 = 1'h0;
    224: T462 = 1'h0;
    225: T462 = 1'h0;
    226: T462 = 1'h0;
    227: T462 = 1'h0;
    228: T462 = 1'h0;
    229: T462 = 1'h0;
    230: T462 = 1'h0;
    231: T462 = 1'h0;
    232: T462 = 1'h0;
    233: T462 = 1'h0;
    234: T462 = 1'h0;
    235: T462 = 1'h0;
    236: T462 = 1'h0;
    237: T462 = 1'h0;
    238: T462 = 1'h0;
    239: T462 = 1'h0;
    240: T462 = 1'h0;
    241: T462 = 1'h0;
    242: T462 = 1'h0;
    243: T462 = 1'h0;
    244: T462 = 1'h0;
    245: T462 = 1'h0;
    246: T462 = 1'h0;
    247: T462 = 1'h0;
    248: T462 = 1'h0;
    249: T462 = 1'h0;
    250: T462 = 1'h0;
    251: T462 = 1'h0;
    252: T462 = 1'h0;
    253: T462 = 1'h0;
    254: T462 = 1'h0;
    255: T462 = 1'h0;
    256: T462 = 1'h0;
    257: T462 = 1'h0;
    258: T462 = 1'h0;
    259: T462 = 1'h0;
    260: T462 = 1'h0;
    261: T462 = 1'h0;
    262: T462 = 1'h0;
    263: T462 = 1'h0;
    264: T462 = 1'h0;
    265: T462 = 1'h0;
    266: T462 = 1'h0;
    267: T462 = 1'h0;
    268: T462 = 1'h0;
    269: T462 = 1'h0;
    270: T462 = 1'h0;
    271: T462 = 1'h0;
    272: T462 = 1'h0;
    273: T462 = 1'h0;
    274: T462 = 1'h0;
    275: T462 = 1'h0;
    276: T462 = 1'h0;
    277: T462 = 1'h0;
    278: T462 = 1'h0;
    279: T462 = 1'h0;
    280: T462 = 1'h0;
    281: T462 = 1'h0;
    282: T462 = 1'h0;
    283: T462 = 1'h0;
    284: T462 = 1'h0;
    285: T462 = 1'h0;
    286: T462 = 1'h0;
    287: T462 = 1'h0;
    288: T462 = 1'h0;
    289: T462 = 1'h0;
    290: T462 = 1'h0;
    291: T462 = 1'h0;
    292: T462 = 1'h0;
    293: T462 = 1'h0;
    294: T462 = 1'h0;
    295: T462 = 1'h0;
    296: T462 = 1'h0;
    297: T462 = 1'h0;
    298: T462 = 1'h0;
    299: T462 = 1'h0;
    300: T462 = 1'h0;
    301: T462 = 1'h0;
    302: T462 = 1'h0;
    303: T462 = 1'h0;
    304: T462 = 1'h0;
    305: T462 = 1'h0;
    306: T462 = 1'h0;
    307: T462 = 1'h0;
    308: T462 = 1'h0;
    309: T462 = 1'h0;
    310: T462 = 1'h0;
    311: T462 = 1'h0;
    312: T462 = 1'h0;
    313: T462 = 1'h0;
    314: T462 = 1'h0;
    315: T462 = 1'h0;
    316: T462 = 1'h0;
    317: T462 = 1'h0;
    318: T462 = 1'h0;
    319: T462 = 1'h0;
    320: T462 = 1'h0;
    321: T462 = 1'h0;
    322: T462 = 1'h0;
    323: T462 = 1'h0;
    324: T462 = 1'h0;
    325: T462 = 1'h0;
    326: T462 = 1'h0;
    327: T462 = 1'h0;
    328: T462 = 1'h0;
    329: T462 = 1'h0;
    330: T462 = 1'h0;
    331: T462 = 1'h0;
    332: T462 = 1'h0;
    333: T462 = 1'h0;
    334: T462 = 1'h0;
    335: T462 = 1'h0;
    336: T462 = 1'h0;
    337: T462 = 1'h0;
    338: T462 = 1'h0;
    339: T462 = 1'h0;
    340: T462 = 1'h0;
    341: T462 = 1'h0;
    342: T462 = 1'h0;
    343: T462 = 1'h0;
    344: T462 = 1'h0;
    345: T462 = 1'h0;
    346: T462 = 1'h0;
    347: T462 = 1'h0;
    348: T462 = 1'h0;
    349: T462 = 1'h0;
    350: T462 = 1'h0;
    351: T462 = 1'h0;
    352: T462 = 1'h0;
    353: T462 = 1'h0;
    354: T462 = 1'h0;
    355: T462 = 1'h0;
    356: T462 = 1'h0;
    357: T462 = 1'h0;
    358: T462 = 1'h0;
    359: T462 = 1'h0;
    360: T462 = 1'h0;
    361: T462 = 1'h0;
    362: T462 = 1'h0;
    363: T462 = 1'h0;
    364: T462 = 1'h0;
    365: T462 = 1'h0;
    366: T462 = 1'h0;
    367: T462 = 1'h0;
    368: T462 = 1'h0;
    369: T462 = 1'h0;
    370: T462 = 1'h0;
    371: T462 = 1'h0;
    372: T462 = 1'h0;
    373: T462 = 1'h0;
    374: T462 = 1'h0;
    375: T462 = 1'h0;
    376: T462 = 1'h0;
    377: T462 = 1'h0;
    378: T462 = 1'h0;
    379: T462 = 1'h0;
    380: T462 = 1'h0;
    381: T462 = 1'h0;
    382: T462 = 1'h0;
    383: T462 = 1'h0;
    384: T462 = 1'h0;
    385: T462 = 1'h0;
    386: T462 = 1'h0;
    387: T462 = 1'h0;
    388: T462 = 1'h0;
    389: T462 = 1'h0;
    390: T462 = 1'h0;
    391: T462 = 1'h0;
    392: T462 = 1'h0;
    393: T462 = 1'h0;
    394: T462 = 1'h0;
    395: T462 = 1'h0;
    396: T462 = 1'h0;
    397: T462 = 1'h0;
    398: T462 = 1'h0;
    399: T462 = 1'h0;
    400: T462 = 1'h0;
    401: T462 = 1'h0;
    402: T462 = 1'h0;
    403: T462 = 1'h0;
    404: T462 = 1'h0;
    405: T462 = 1'h0;
    406: T462 = 1'h0;
    407: T462 = 1'h0;
    408: T462 = 1'h0;
    409: T462 = 1'h0;
    410: T462 = 1'h0;
    411: T462 = 1'h0;
    412: T462 = 1'h0;
    413: T462 = 1'h0;
    414: T462 = 1'h0;
    415: T462 = 1'h0;
    416: T462 = 1'h0;
    417: T462 = 1'h0;
    418: T462 = 1'h0;
    419: T462 = 1'h0;
    420: T462 = 1'h0;
    421: T462 = 1'h0;
    422: T462 = 1'h0;
    423: T462 = 1'h0;
    424: T462 = 1'h0;
    425: T462 = 1'h0;
    426: T462 = 1'h0;
    427: T462 = 1'h0;
    428: T462 = 1'h0;
    429: T462 = 1'h0;
    430: T462 = 1'h0;
    431: T462 = 1'h0;
    432: T462 = 1'h0;
    433: T462 = 1'h0;
    434: T462 = 1'h0;
    435: T462 = 1'h0;
    436: T462 = 1'h0;
    437: T462 = 1'h0;
    438: T462 = 1'h0;
    439: T462 = 1'h0;
    440: T462 = 1'h0;
    441: T462 = 1'h0;
    442: T462 = 1'h0;
    443: T462 = 1'h0;
    444: T462 = 1'h0;
    445: T462 = 1'h0;
    446: T462 = 1'h0;
    447: T462 = 1'h0;
    448: T462 = 1'h0;
    449: T462 = 1'h0;
    450: T462 = 1'h0;
    451: T462 = 1'h0;
    452: T462 = 1'h0;
    453: T462 = 1'h0;
    454: T462 = 1'h0;
    455: T462 = 1'h0;
    456: T462 = 1'h0;
    457: T462 = 1'h0;
    458: T462 = 1'h0;
    459: T462 = 1'h0;
    460: T462 = 1'h0;
    461: T462 = 1'h0;
    462: T462 = 1'h0;
    463: T462 = 1'h0;
    464: T462 = 1'h0;
    465: T462 = 1'h0;
    466: T462 = 1'h0;
    467: T462 = 1'h0;
    468: T462 = 1'h0;
    469: T462 = 1'h0;
    470: T462 = 1'h0;
    471: T462 = 1'h0;
    472: T462 = 1'h0;
    473: T462 = 1'h0;
    474: T462 = 1'h0;
    475: T462 = 1'h0;
    476: T462 = 1'h0;
    477: T462 = 1'h0;
    478: T462 = 1'h0;
    479: T462 = 1'h0;
    480: T462 = 1'h0;
    481: T462 = 1'h0;
    482: T462 = 1'h0;
    483: T462 = 1'h0;
    484: T462 = 1'h0;
    485: T462 = 1'h0;
    486: T462 = 1'h0;
    487: T462 = 1'h0;
    488: T462 = 1'h0;
    489: T462 = 1'h0;
    490: T462 = 1'h0;
    491: T462 = 1'h0;
    492: T462 = 1'h0;
    493: T462 = 1'h0;
    494: T462 = 1'h0;
    495: T462 = 1'h0;
    496: T462 = 1'h0;
    497: T462 = 1'h0;
    498: T462 = 1'h0;
    499: T462 = 1'h0;
    500: T462 = 1'h0;
    501: T462 = 1'h0;
    502: T462 = 1'h0;
    503: T462 = 1'h0;
    504: T462 = 1'h0;
    505: T462 = 1'h0;
    506: T462 = 1'h0;
    507: T462 = 1'h0;
    508: T462 = 1'h0;
    509: T462 = 1'h0;
    510: T462 = 1'h0;
    511: T462 = 1'h0;
    512: T462 = 1'h0;
    513: T462 = 1'h0;
    514: T462 = 1'h0;
    515: T462 = 1'h0;
    516: T462 = 1'h0;
    517: T462 = 1'h0;
    518: T462 = 1'h0;
    519: T462 = 1'h0;
    520: T462 = 1'h0;
    521: T462 = 1'h0;
    522: T462 = 1'h0;
    523: T462 = 1'h0;
    524: T462 = 1'h0;
    525: T462 = 1'h0;
    526: T462 = 1'h0;
    527: T462 = 1'h0;
    528: T462 = 1'h0;
    529: T462 = 1'h0;
    530: T462 = 1'h0;
    531: T462 = 1'h0;
    532: T462 = 1'h0;
    533: T462 = 1'h0;
    534: T462 = 1'h0;
    535: T462 = 1'h0;
    536: T462 = 1'h0;
    537: T462 = 1'h0;
    538: T462 = 1'h0;
    539: T462 = 1'h0;
    540: T462 = 1'h0;
    541: T462 = 1'h0;
    542: T462 = 1'h0;
    543: T462 = 1'h0;
    544: T462 = 1'h0;
    545: T462 = 1'h0;
    546: T462 = 1'h0;
    547: T462 = 1'h0;
    548: T462 = 1'h0;
    549: T462 = 1'h0;
    550: T462 = 1'h0;
    551: T462 = 1'h0;
    552: T462 = 1'h0;
    553: T462 = 1'h0;
    554: T462 = 1'h0;
    555: T462 = 1'h0;
    556: T462 = 1'h0;
    557: T462 = 1'h0;
    558: T462 = 1'h0;
    559: T462 = 1'h0;
    560: T462 = 1'h0;
    561: T462 = 1'h0;
    562: T462 = 1'h0;
    563: T462 = 1'h0;
    564: T462 = 1'h0;
    565: T462 = 1'h0;
    566: T462 = 1'h0;
    567: T462 = 1'h0;
    568: T462 = 1'h0;
    569: T462 = 1'h0;
    570: T462 = 1'h0;
    571: T462 = 1'h0;
    572: T462 = 1'h0;
    573: T462 = 1'h0;
    574: T462 = 1'h0;
    575: T462 = 1'h0;
    576: T462 = 1'h0;
    577: T462 = 1'h0;
    578: T462 = 1'h0;
    579: T462 = 1'h0;
    580: T462 = 1'h0;
    581: T462 = 1'h0;
    582: T462 = 1'h0;
    583: T462 = 1'h0;
    584: T462 = 1'h0;
    585: T462 = 1'h0;
    586: T462 = 1'h0;
    587: T462 = 1'h0;
    588: T462 = 1'h0;
    589: T462 = 1'h0;
    590: T462 = 1'h0;
    591: T462 = 1'h0;
    592: T462 = 1'h0;
    593: T462 = 1'h0;
    594: T462 = 1'h0;
    595: T462 = 1'h0;
    596: T462 = 1'h0;
    597: T462 = 1'h0;
    598: T462 = 1'h0;
    599: T462 = 1'h0;
    600: T462 = 1'h0;
    601: T462 = 1'h0;
    602: T462 = 1'h0;
    603: T462 = 1'h0;
    604: T462 = 1'h0;
    605: T462 = 1'h0;
    606: T462 = 1'h0;
    607: T462 = 1'h0;
    608: T462 = 1'h0;
    609: T462 = 1'h0;
    610: T462 = 1'h0;
    611: T462 = 1'h0;
    612: T462 = 1'h0;
    613: T462 = 1'h0;
    614: T462 = 1'h0;
    615: T462 = 1'h0;
    616: T462 = 1'h0;
    617: T462 = 1'h0;
    618: T462 = 1'h0;
    619: T462 = 1'h0;
    620: T462 = 1'h0;
    621: T462 = 1'h0;
    622: T462 = 1'h0;
    623: T462 = 1'h0;
    624: T462 = 1'h0;
    625: T462 = 1'h0;
    626: T462 = 1'h0;
    627: T462 = 1'h0;
    628: T462 = 1'h0;
    629: T462 = 1'h0;
    630: T462 = 1'h0;
    631: T462 = 1'h0;
    632: T462 = 1'h0;
    633: T462 = 1'h0;
    634: T462 = 1'h0;
    635: T462 = 1'h0;
    636: T462 = 1'h0;
    637: T462 = 1'h0;
    638: T462 = 1'h0;
    639: T462 = 1'h0;
    640: T462 = 1'h0;
    641: T462 = 1'h0;
    642: T462 = 1'h0;
    643: T462 = 1'h0;
    644: T462 = 1'h0;
    645: T462 = 1'h0;
    646: T462 = 1'h0;
    647: T462 = 1'h0;
    648: T462 = 1'h0;
    649: T462 = 1'h0;
    650: T462 = 1'h0;
    651: T462 = 1'h0;
    652: T462 = 1'h0;
    653: T462 = 1'h0;
    654: T462 = 1'h0;
    655: T462 = 1'h0;
    656: T462 = 1'h0;
    657: T462 = 1'h0;
    658: T462 = 1'h0;
    659: T462 = 1'h0;
    660: T462 = 1'h0;
    661: T462 = 1'h0;
    662: T462 = 1'h0;
    663: T462 = 1'h0;
    664: T462 = 1'h0;
    665: T462 = 1'h0;
    666: T462 = 1'h0;
    667: T462 = 1'h0;
    668: T462 = 1'h0;
    669: T462 = 1'h0;
    670: T462 = 1'h0;
    671: T462 = 1'h0;
    672: T462 = 1'h0;
    673: T462 = 1'h0;
    674: T462 = 1'h0;
    675: T462 = 1'h0;
    676: T462 = 1'h0;
    677: T462 = 1'h0;
    678: T462 = 1'h0;
    679: T462 = 1'h0;
    680: T462 = 1'h0;
    681: T462 = 1'h0;
    682: T462 = 1'h0;
    683: T462 = 1'h0;
    684: T462 = 1'h0;
    685: T462 = 1'h0;
    686: T462 = 1'h0;
    687: T462 = 1'h0;
    688: T462 = 1'h0;
    689: T462 = 1'h0;
    690: T462 = 1'h0;
    691: T462 = 1'h0;
    692: T462 = 1'h0;
    693: T462 = 1'h0;
    694: T462 = 1'h0;
    695: T462 = 1'h0;
    696: T462 = 1'h0;
    697: T462 = 1'h0;
    698: T462 = 1'h0;
    699: T462 = 1'h0;
    700: T462 = 1'h0;
    701: T462 = 1'h0;
    702: T462 = 1'h0;
    703: T462 = 1'h0;
    704: T462 = 1'h0;
    705: T462 = 1'h0;
    706: T462 = 1'h0;
    707: T462 = 1'h0;
    708: T462 = 1'h0;
    709: T462 = 1'h0;
    710: T462 = 1'h0;
    711: T462 = 1'h0;
    712: T462 = 1'h0;
    713: T462 = 1'h0;
    714: T462 = 1'h0;
    715: T462 = 1'h0;
    716: T462 = 1'h0;
    717: T462 = 1'h0;
    718: T462 = 1'h0;
    719: T462 = 1'h0;
    720: T462 = 1'h0;
    721: T462 = 1'h0;
    722: T462 = 1'h0;
    723: T462 = 1'h0;
    724: T462 = 1'h0;
    725: T462 = 1'h0;
    726: T462 = 1'h0;
    727: T462 = 1'h0;
    728: T462 = 1'h0;
    729: T462 = 1'h0;
    730: T462 = 1'h0;
    731: T462 = 1'h0;
    732: T462 = 1'h0;
    733: T462 = 1'h0;
    734: T462 = 1'h0;
    735: T462 = 1'h0;
    736: T462 = 1'h0;
    737: T462 = 1'h0;
    738: T462 = 1'h0;
    739: T462 = 1'h0;
    740: T462 = 1'h0;
    741: T462 = 1'h0;
    742: T462 = 1'h0;
    743: T462 = 1'h0;
    744: T462 = 1'h0;
    745: T462 = 1'h0;
    746: T462 = 1'h0;
    747: T462 = 1'h0;
    748: T462 = 1'h0;
    749: T462 = 1'h0;
    750: T462 = 1'h0;
    751: T462 = 1'h0;
    752: T462 = 1'h0;
    753: T462 = 1'h0;
    754: T462 = 1'h0;
    755: T462 = 1'h0;
    756: T462 = 1'h0;
    757: T462 = 1'h0;
    758: T462 = 1'h0;
    759: T462 = 1'h0;
    760: T462 = 1'h0;
    761: T462 = 1'h0;
    762: T462 = 1'h0;
    763: T462 = 1'h0;
    764: T462 = 1'h0;
    765: T462 = 1'h0;
    766: T462 = 1'h0;
    767: T462 = 1'h0;
    768: T462 = 1'h0;
    769: T462 = 1'h0;
    770: T462 = 1'h0;
    771: T462 = 1'h0;
    772: T462 = 1'h0;
    773: T462 = 1'h0;
    774: T462 = 1'h0;
    775: T462 = 1'h0;
    776: T462 = 1'h0;
    777: T462 = 1'h0;
    778: T462 = 1'h0;
    779: T462 = 1'h0;
    780: T462 = 1'h0;
    781: T462 = 1'h0;
    782: T462 = 1'h0;
    783: T462 = 1'h0;
    784: T462 = 1'h0;
    785: T462 = 1'h0;
    786: T462 = 1'h0;
    787: T462 = 1'h0;
    788: T462 = 1'h0;
    789: T462 = 1'h0;
    790: T462 = 1'h0;
    791: T462 = 1'h0;
    792: T462 = 1'h0;
    793: T462 = 1'h0;
    794: T462 = 1'h0;
    795: T462 = 1'h0;
    796: T462 = 1'h0;
    797: T462 = 1'h0;
    798: T462 = 1'h0;
    799: T462 = 1'h0;
    800: T462 = 1'h0;
    801: T462 = 1'h0;
    802: T462 = 1'h0;
    803: T462 = 1'h0;
    804: T462 = 1'h0;
    805: T462 = 1'h0;
    806: T462 = 1'h0;
    807: T462 = 1'h0;
    808: T462 = 1'h0;
    809: T462 = 1'h0;
    810: T462 = 1'h0;
    811: T462 = 1'h0;
    812: T462 = 1'h0;
    813: T462 = 1'h0;
    814: T462 = 1'h0;
    815: T462 = 1'h0;
    816: T462 = 1'h0;
    817: T462 = 1'h0;
    818: T462 = 1'h0;
    819: T462 = 1'h0;
    820: T462 = 1'h0;
    821: T462 = 1'h0;
    822: T462 = 1'h0;
    823: T462 = 1'h0;
    824: T462 = 1'h0;
    825: T462 = 1'h0;
    826: T462 = 1'h0;
    827: T462 = 1'h0;
    828: T462 = 1'h0;
    829: T462 = 1'h0;
    830: T462 = 1'h0;
    831: T462 = 1'h0;
    832: T462 = 1'h0;
    833: T462 = 1'h0;
    834: T462 = 1'h0;
    835: T462 = 1'h0;
    836: T462 = 1'h0;
    837: T462 = 1'h0;
    838: T462 = 1'h0;
    839: T462 = 1'h0;
    840: T462 = 1'h0;
    841: T462 = 1'h0;
    842: T462 = 1'h0;
    843: T462 = 1'h0;
    844: T462 = 1'h0;
    845: T462 = 1'h0;
    846: T462 = 1'h0;
    847: T462 = 1'h0;
    848: T462 = 1'h0;
    849: T462 = 1'h0;
    850: T462 = 1'h0;
    851: T462 = 1'h0;
    852: T462 = 1'h0;
    853: T462 = 1'h0;
    854: T462 = 1'h0;
    855: T462 = 1'h0;
    856: T462 = 1'h0;
    857: T462 = 1'h0;
    858: T462 = 1'h0;
    859: T462 = 1'h0;
    860: T462 = 1'h0;
    861: T462 = 1'h0;
    862: T462 = 1'h0;
    863: T462 = 1'h0;
    864: T462 = 1'h0;
    865: T462 = 1'h0;
    866: T462 = 1'h0;
    867: T462 = 1'h0;
    868: T462 = 1'h0;
    869: T462 = 1'h0;
    870: T462 = 1'h0;
    871: T462 = 1'h0;
    872: T462 = 1'h0;
    873: T462 = 1'h0;
    874: T462 = 1'h0;
    875: T462 = 1'h0;
    876: T462 = 1'h0;
    877: T462 = 1'h0;
    878: T462 = 1'h0;
    879: T462 = 1'h0;
    880: T462 = 1'h0;
    881: T462 = 1'h0;
    882: T462 = 1'h0;
    883: T462 = 1'h0;
    884: T462 = 1'h0;
    885: T462 = 1'h0;
    886: T462 = 1'h0;
    887: T462 = 1'h0;
    888: T462 = 1'h0;
    889: T462 = 1'h0;
    890: T462 = 1'h0;
    891: T462 = 1'h0;
    892: T462 = 1'h0;
    893: T462 = 1'h0;
    894: T462 = 1'h0;
    895: T462 = 1'h0;
    896: T462 = 1'h0;
    897: T462 = 1'h0;
    898: T462 = 1'h0;
    899: T462 = 1'h0;
    900: T462 = 1'h0;
    901: T462 = 1'h0;
    902: T462 = 1'h0;
    903: T462 = 1'h0;
    904: T462 = 1'h0;
    905: T462 = 1'h0;
    906: T462 = 1'h0;
    907: T462 = 1'h0;
    908: T462 = 1'h0;
    909: T462 = 1'h0;
    910: T462 = 1'h0;
    911: T462 = 1'h0;
    912: T462 = 1'h0;
    913: T462 = 1'h0;
    914: T462 = 1'h0;
    915: T462 = 1'h0;
    916: T462 = 1'h0;
    917: T462 = 1'h0;
    918: T462 = 1'h0;
    919: T462 = 1'h0;
    920: T462 = 1'h0;
    921: T462 = 1'h0;
    922: T462 = 1'h0;
    923: T462 = 1'h0;
    924: T462 = 1'h0;
    925: T462 = 1'h0;
    926: T462 = 1'h0;
    927: T462 = 1'h0;
    928: T462 = 1'h0;
    929: T462 = 1'h0;
    930: T462 = 1'h0;
    931: T462 = 1'h0;
    932: T462 = 1'h0;
    933: T462 = 1'h0;
    934: T462 = 1'h0;
    935: T462 = 1'h0;
    936: T462 = 1'h0;
    937: T462 = 1'h0;
    938: T462 = 1'h0;
    939: T462 = 1'h0;
    940: T462 = 1'h0;
    941: T462 = 1'h0;
    942: T462 = 1'h0;
    943: T462 = 1'h0;
    944: T462 = 1'h0;
    945: T462 = 1'h0;
    946: T462 = 1'h0;
    947: T462 = 1'h0;
    948: T462 = 1'h0;
    949: T462 = 1'h0;
    950: T462 = 1'h0;
    951: T462 = 1'h0;
    952: T462 = 1'h0;
    953: T462 = 1'h0;
    954: T462 = 1'h0;
    955: T462 = 1'h0;
    956: T462 = 1'h0;
    957: T462 = 1'h0;
    958: T462 = 1'h0;
    959: T462 = 1'h0;
    960: T462 = 1'h0;
    961: T462 = 1'h0;
    962: T462 = 1'h0;
    963: T462 = 1'h0;
    964: T462 = 1'h0;
    965: T462 = 1'h0;
    966: T462 = 1'h0;
    967: T462 = 1'h0;
    968: T462 = 1'h0;
    969: T462 = 1'h0;
    970: T462 = 1'h0;
    971: T462 = 1'h0;
    972: T462 = 1'h0;
    973: T462 = 1'h0;
    974: T462 = 1'h0;
    975: T462 = 1'h0;
    976: T462 = 1'h0;
    977: T462 = 1'h0;
    978: T462 = 1'h0;
    979: T462 = 1'h0;
    980: T462 = 1'h0;
    981: T462 = 1'h0;
    982: T462 = 1'h0;
    983: T462 = 1'h0;
    984: T462 = 1'h0;
    985: T462 = 1'h0;
    986: T462 = 1'h0;
    987: T462 = 1'h0;
    988: T462 = 1'h0;
    989: T462 = 1'h0;
    990: T462 = 1'h0;
    991: T462 = 1'h0;
    992: T462 = 1'h0;
    993: T462 = 1'h0;
    994: T462 = 1'h0;
    995: T462 = 1'h0;
    996: T462 = 1'h0;
    997: T462 = 1'h0;
    998: T462 = 1'h0;
    999: T462 = 1'h0;
    1000: T462 = 1'h0;
    1001: T462 = 1'h0;
    1002: T462 = 1'h0;
    1003: T462 = 1'h0;
    1004: T462 = 1'h0;
    1005: T462 = 1'h0;
    1006: T462 = 1'h0;
    1007: T462 = 1'h0;
    1008: T462 = 1'h0;
    1009: T462 = 1'h0;
    1010: T462 = 1'h0;
    1011: T462 = 1'h0;
    1012: T462 = 1'h0;
    1013: T462 = 1'h0;
    1014: T462 = 1'h0;
    1015: T462 = 1'h0;
    1016: T462 = 1'h0;
    1017: T462 = 1'h0;
    1018: T462 = 1'h0;
    1019: T462 = 1'h0;
    1020: T462 = 1'h0;
    1021: T462 = 1'h0;
    1022: T462 = 1'h0;
    1023: T462 = 1'h0;
    1024: T462 = 1'h0;
    1025: T462 = 1'h0;
    1026: T462 = 1'h0;
    1027: T462 = 1'h0;
    1028: T462 = 1'h0;
    1029: T462 = 1'h0;
    1030: T462 = 1'h0;
    1031: T462 = 1'h0;
    1032: T462 = 1'h0;
    1033: T462 = 1'h0;
    1034: T462 = 1'h0;
    1035: T462 = 1'h0;
    1036: T462 = 1'h0;
    1037: T462 = 1'h0;
    1038: T462 = 1'h0;
    1039: T462 = 1'h0;
    1040: T462 = 1'h0;
    1041: T462 = 1'h0;
    1042: T462 = 1'h0;
    1043: T462 = 1'h0;
    1044: T462 = 1'h0;
    1045: T462 = 1'h0;
    1046: T462 = 1'h0;
    1047: T462 = 1'h0;
    1048: T462 = 1'h0;
    1049: T462 = 1'h0;
    1050: T462 = 1'h0;
    1051: T462 = 1'h0;
    1052: T462 = 1'h0;
    1053: T462 = 1'h0;
    1054: T462 = 1'h0;
    1055: T462 = 1'h0;
    1056: T462 = 1'h0;
    1057: T462 = 1'h0;
    1058: T462 = 1'h0;
    1059: T462 = 1'h0;
    1060: T462 = 1'h0;
    1061: T462 = 1'h0;
    1062: T462 = 1'h0;
    1063: T462 = 1'h0;
    1064: T462 = 1'h0;
    1065: T462 = 1'h0;
    1066: T462 = 1'h0;
    1067: T462 = 1'h0;
    1068: T462 = 1'h0;
    1069: T462 = 1'h0;
    1070: T462 = 1'h0;
    1071: T462 = 1'h0;
    1072: T462 = 1'h0;
    1073: T462 = 1'h0;
    1074: T462 = 1'h0;
    1075: T462 = 1'h0;
    1076: T462 = 1'h0;
    1077: T462 = 1'h0;
    1078: T462 = 1'h0;
    1079: T462 = 1'h0;
    1080: T462 = 1'h0;
    1081: T462 = 1'h0;
    1082: T462 = 1'h0;
    1083: T462 = 1'h0;
    1084: T462 = 1'h0;
    1085: T462 = 1'h0;
    1086: T462 = 1'h0;
    1087: T462 = 1'h0;
    1088: T462 = 1'h0;
    1089: T462 = 1'h0;
    1090: T462 = 1'h0;
    1091: T462 = 1'h0;
    1092: T462 = 1'h0;
    1093: T462 = 1'h0;
    1094: T462 = 1'h0;
    1095: T462 = 1'h0;
    1096: T462 = 1'h0;
    1097: T462 = 1'h0;
    1098: T462 = 1'h0;
    1099: T462 = 1'h0;
    1100: T462 = 1'h0;
    1101: T462 = 1'h0;
    1102: T462 = 1'h0;
    1103: T462 = 1'h0;
    1104: T462 = 1'h0;
    1105: T462 = 1'h0;
    1106: T462 = 1'h0;
    1107: T462 = 1'h0;
    1108: T462 = 1'h0;
    1109: T462 = 1'h0;
    1110: T462 = 1'h0;
    1111: T462 = 1'h0;
    1112: T462 = 1'h0;
    1113: T462 = 1'h0;
    1114: T462 = 1'h0;
    1115: T462 = 1'h0;
    1116: T462 = 1'h0;
    1117: T462 = 1'h0;
    1118: T462 = 1'h0;
    1119: T462 = 1'h0;
    1120: T462 = 1'h0;
    1121: T462 = 1'h0;
    1122: T462 = 1'h0;
    1123: T462 = 1'h0;
    1124: T462 = 1'h0;
    1125: T462 = 1'h0;
    1126: T462 = 1'h0;
    1127: T462 = 1'h0;
    1128: T462 = 1'h0;
    1129: T462 = 1'h0;
    1130: T462 = 1'h0;
    1131: T462 = 1'h0;
    1132: T462 = 1'h0;
    1133: T462 = 1'h0;
    1134: T462 = 1'h0;
    1135: T462 = 1'h0;
    1136: T462 = 1'h0;
    1137: T462 = 1'h0;
    1138: T462 = 1'h0;
    1139: T462 = 1'h0;
    1140: T462 = 1'h0;
    1141: T462 = 1'h0;
    1142: T462 = 1'h0;
    1143: T462 = 1'h0;
    1144: T462 = 1'h0;
    1145: T462 = 1'h0;
    1146: T462 = 1'h0;
    1147: T462 = 1'h0;
    1148: T462 = 1'h0;
    1149: T462 = 1'h0;
    1150: T462 = 1'h0;
    1151: T462 = 1'h0;
    1152: T462 = 1'h0;
    1153: T462 = 1'h0;
    1154: T462 = 1'h0;
    1155: T462 = 1'h0;
    1156: T462 = 1'h0;
    1157: T462 = 1'h0;
    1158: T462 = 1'h0;
    1159: T462 = 1'h0;
    1160: T462 = 1'h0;
    1161: T462 = 1'h0;
    1162: T462 = 1'h0;
    1163: T462 = 1'h0;
    1164: T462 = 1'h0;
    1165: T462 = 1'h0;
    1166: T462 = 1'h0;
    1167: T462 = 1'h0;
    1168: T462 = 1'h0;
    1169: T462 = 1'h0;
    1170: T462 = 1'h0;
    1171: T462 = 1'h0;
    1172: T462 = 1'h0;
    1173: T462 = 1'h0;
    1174: T462 = 1'h0;
    1175: T462 = 1'h0;
    1176: T462 = 1'h0;
    1177: T462 = 1'h0;
    1178: T462 = 1'h0;
    1179: T462 = 1'h0;
    1180: T462 = 1'h0;
    1181: T462 = 1'h0;
    1182: T462 = 1'h0;
    1183: T462 = 1'h0;
    1184: T462 = 1'h0;
    1185: T462 = 1'h0;
    1186: T462 = 1'h0;
    1187: T462 = 1'h0;
    1188: T462 = 1'h0;
    1189: T462 = 1'h0;
    1190: T462 = 1'h0;
    1191: T462 = 1'h0;
    1192: T462 = 1'h0;
    1193: T462 = 1'h0;
    1194: T462 = 1'h0;
    1195: T462 = 1'h0;
    1196: T462 = 1'h0;
    1197: T462 = 1'h0;
    1198: T462 = 1'h0;
    1199: T462 = 1'h0;
    1200: T462 = 1'h0;
    1201: T462 = 1'h0;
    1202: T462 = 1'h0;
    1203: T462 = 1'h0;
    1204: T462 = 1'h0;
    1205: T462 = 1'h0;
    1206: T462 = 1'h0;
    1207: T462 = 1'h0;
    1208: T462 = 1'h0;
    1209: T462 = 1'h0;
    1210: T462 = 1'h0;
    1211: T462 = 1'h0;
    1212: T462 = 1'h0;
    1213: T462 = 1'h0;
    1214: T462 = 1'h0;
    1215: T462 = 1'h0;
    1216: T462 = 1'h0;
    1217: T462 = 1'h0;
    1218: T462 = 1'h0;
    1219: T462 = 1'h0;
    1220: T462 = 1'h0;
    1221: T462 = 1'h0;
    1222: T462 = 1'h0;
    1223: T462 = 1'h0;
    1224: T462 = 1'h0;
    1225: T462 = 1'h0;
    1226: T462 = 1'h0;
    1227: T462 = 1'h0;
    1228: T462 = 1'h0;
    1229: T462 = 1'h0;
    1230: T462 = 1'h0;
    1231: T462 = 1'h0;
    1232: T462 = 1'h0;
    1233: T462 = 1'h0;
    1234: T462 = 1'h0;
    1235: T462 = 1'h0;
    1236: T462 = 1'h0;
    1237: T462 = 1'h0;
    1238: T462 = 1'h0;
    1239: T462 = 1'h0;
    1240: T462 = 1'h0;
    1241: T462 = 1'h0;
    1242: T462 = 1'h0;
    1243: T462 = 1'h0;
    1244: T462 = 1'h0;
    1245: T462 = 1'h0;
    1246: T462 = 1'h0;
    1247: T462 = 1'h0;
    1248: T462 = 1'h0;
    1249: T462 = 1'h0;
    1250: T462 = 1'h0;
    1251: T462 = 1'h0;
    1252: T462 = 1'h0;
    1253: T462 = 1'h0;
    1254: T462 = 1'h0;
    1255: T462 = 1'h0;
    1256: T462 = 1'h0;
    1257: T462 = 1'h0;
    1258: T462 = 1'h0;
    1259: T462 = 1'h0;
    1260: T462 = 1'h0;
    1261: T462 = 1'h0;
    1262: T462 = 1'h0;
    1263: T462 = 1'h0;
    1264: T462 = 1'h0;
    1265: T462 = 1'h0;
    1266: T462 = 1'h0;
    1267: T462 = 1'h0;
    1268: T462 = 1'h0;
    1269: T462 = 1'h0;
    1270: T462 = 1'h0;
    1271: T462 = 1'h0;
    1272: T462 = 1'h0;
    1273: T462 = 1'h0;
    1274: T462 = 1'h0;
    1275: T462 = 1'h0;
    1276: T462 = 1'h0;
    1277: T462 = 1'h0;
    1278: T462 = 1'h0;
    1279: T462 = 1'h0;
    1280: T462 = 1'h1;
    1281: T462 = 1'h1;
    1282: T462 = 1'h1;
    1283: T462 = 1'h1;
    1284: T462 = 1'h1;
    1285: T462 = 1'h1;
    1286: T462 = 1'h1;
    1287: T462 = 1'h1;
    1288: T462 = 1'h1;
    1289: T462 = 1'h1;
    1290: T462 = 1'h1;
    1291: T462 = 1'h1;
    1292: T462 = 1'h1;
    1293: T462 = 1'h1;
    1294: T462 = 1'h1;
    1295: T462 = 1'h1;
    1296: T462 = 1'h0;
    1297: T462 = 1'h0;
    1298: T462 = 1'h0;
    1299: T462 = 1'h0;
    1300: T462 = 1'h0;
    1301: T462 = 1'h0;
    1302: T462 = 1'h0;
    1303: T462 = 1'h0;
    1304: T462 = 1'h0;
    1305: T462 = 1'h0;
    1306: T462 = 1'h0;
    1307: T462 = 1'h0;
    1308: T462 = 1'h0;
    1309: T462 = 1'h1;
    1310: T462 = 1'h1;
    1311: T462 = 1'h1;
    1312: T462 = 1'h1;
    1313: T462 = 1'h1;
    1314: T462 = 1'h1;
    1315: T462 = 1'h1;
    1316: T462 = 1'h0;
    1317: T462 = 1'h0;
    1318: T462 = 1'h0;
    1319: T462 = 1'h0;
    1320: T462 = 1'h0;
    1321: T462 = 1'h0;
    1322: T462 = 1'h0;
    1323: T462 = 1'h0;
    1324: T462 = 1'h0;
    1325: T462 = 1'h0;
    1326: T462 = 1'h0;
    1327: T462 = 1'h0;
    1328: T462 = 1'h0;
    1329: T462 = 1'h0;
    1330: T462 = 1'h0;
    1331: T462 = 1'h0;
    1332: T462 = 1'h0;
    1333: T462 = 1'h0;
    1334: T462 = 1'h0;
    1335: T462 = 1'h0;
    1336: T462 = 1'h0;
    1337: T462 = 1'h0;
    1338: T462 = 1'h0;
    1339: T462 = 1'h0;
    1340: T462 = 1'h0;
    1341: T462 = 1'h0;
    1342: T462 = 1'h0;
    1343: T462 = 1'h0;
    1344: T462 = 1'h0;
    1345: T462 = 1'h0;
    1346: T462 = 1'h0;
    1347: T462 = 1'h0;
    1348: T462 = 1'h0;
    1349: T462 = 1'h0;
    1350: T462 = 1'h0;
    1351: T462 = 1'h0;
    1352: T462 = 1'h0;
    1353: T462 = 1'h0;
    1354: T462 = 1'h0;
    1355: T462 = 1'h0;
    1356: T462 = 1'h0;
    1357: T462 = 1'h0;
    1358: T462 = 1'h0;
    1359: T462 = 1'h0;
    1360: T462 = 1'h0;
    1361: T462 = 1'h0;
    1362: T462 = 1'h0;
    1363: T462 = 1'h0;
    1364: T462 = 1'h0;
    1365: T462 = 1'h0;
    1366: T462 = 1'h0;
    1367: T462 = 1'h0;
    1368: T462 = 1'h0;
    1369: T462 = 1'h0;
    1370: T462 = 1'h0;
    1371: T462 = 1'h0;
    1372: T462 = 1'h0;
    1373: T462 = 1'h0;
    1374: T462 = 1'h0;
    1375: T462 = 1'h0;
    1376: T462 = 1'h0;
    1377: T462 = 1'h0;
    1378: T462 = 1'h0;
    1379: T462 = 1'h0;
    1380: T462 = 1'h0;
    1381: T462 = 1'h0;
    1382: T462 = 1'h0;
    1383: T462 = 1'h0;
    1384: T462 = 1'h0;
    1385: T462 = 1'h0;
    1386: T462 = 1'h0;
    1387: T462 = 1'h0;
    1388: T462 = 1'h0;
    1389: T462 = 1'h0;
    1390: T462 = 1'h0;
    1391: T462 = 1'h0;
    1392: T462 = 1'h0;
    1393: T462 = 1'h0;
    1394: T462 = 1'h0;
    1395: T462 = 1'h0;
    1396: T462 = 1'h0;
    1397: T462 = 1'h0;
    1398: T462 = 1'h0;
    1399: T462 = 1'h0;
    1400: T462 = 1'h0;
    1401: T462 = 1'h0;
    1402: T462 = 1'h0;
    1403: T462 = 1'h0;
    1404: T462 = 1'h0;
    1405: T462 = 1'h0;
    1406: T462 = 1'h0;
    1407: T462 = 1'h0;
    1408: T462 = 1'h0;
    1409: T462 = 1'h0;
    1410: T462 = 1'h0;
    1411: T462 = 1'h0;
    1412: T462 = 1'h0;
    1413: T462 = 1'h0;
    1414: T462 = 1'h0;
    1415: T462 = 1'h0;
    1416: T462 = 1'h0;
    1417: T462 = 1'h0;
    1418: T462 = 1'h0;
    1419: T462 = 1'h0;
    1420: T462 = 1'h0;
    1421: T462 = 1'h0;
    1422: T462 = 1'h0;
    1423: T462 = 1'h0;
    1424: T462 = 1'h0;
    1425: T462 = 1'h0;
    1426: T462 = 1'h0;
    1427: T462 = 1'h0;
    1428: T462 = 1'h0;
    1429: T462 = 1'h0;
    1430: T462 = 1'h0;
    1431: T462 = 1'h0;
    1432: T462 = 1'h0;
    1433: T462 = 1'h0;
    1434: T462 = 1'h0;
    1435: T462 = 1'h0;
    1436: T462 = 1'h0;
    1437: T462 = 1'h0;
    1438: T462 = 1'h0;
    1439: T462 = 1'h0;
    1440: T462 = 1'h0;
    1441: T462 = 1'h0;
    1442: T462 = 1'h0;
    1443: T462 = 1'h0;
    1444: T462 = 1'h0;
    1445: T462 = 1'h0;
    1446: T462 = 1'h0;
    1447: T462 = 1'h0;
    1448: T462 = 1'h0;
    1449: T462 = 1'h0;
    1450: T462 = 1'h0;
    1451: T462 = 1'h0;
    1452: T462 = 1'h0;
    1453: T462 = 1'h0;
    1454: T462 = 1'h0;
    1455: T462 = 1'h0;
    1456: T462 = 1'h0;
    1457: T462 = 1'h0;
    1458: T462 = 1'h0;
    1459: T462 = 1'h0;
    1460: T462 = 1'h0;
    1461: T462 = 1'h0;
    1462: T462 = 1'h0;
    1463: T462 = 1'h0;
    1464: T462 = 1'h0;
    1465: T462 = 1'h0;
    1466: T462 = 1'h0;
    1467: T462 = 1'h0;
    1468: T462 = 1'h0;
    1469: T462 = 1'h0;
    1470: T462 = 1'h0;
    1471: T462 = 1'h0;
    1472: T462 = 1'h0;
    1473: T462 = 1'h0;
    1474: T462 = 1'h0;
    1475: T462 = 1'h0;
    1476: T462 = 1'h0;
    1477: T462 = 1'h0;
    1478: T462 = 1'h0;
    1479: T462 = 1'h0;
    1480: T462 = 1'h0;
    1481: T462 = 1'h0;
    1482: T462 = 1'h0;
    1483: T462 = 1'h0;
    1484: T462 = 1'h0;
    1485: T462 = 1'h0;
    1486: T462 = 1'h0;
    1487: T462 = 1'h0;
    1488: T462 = 1'h0;
    1489: T462 = 1'h0;
    1490: T462 = 1'h0;
    1491: T462 = 1'h0;
    1492: T462 = 1'h0;
    1493: T462 = 1'h0;
    1494: T462 = 1'h0;
    1495: T462 = 1'h0;
    1496: T462 = 1'h0;
    1497: T462 = 1'h0;
    1498: T462 = 1'h0;
    1499: T462 = 1'h0;
    1500: T462 = 1'h0;
    1501: T462 = 1'h0;
    1502: T462 = 1'h0;
    1503: T462 = 1'h0;
    1504: T462 = 1'h0;
    1505: T462 = 1'h0;
    1506: T462 = 1'h0;
    1507: T462 = 1'h0;
    1508: T462 = 1'h0;
    1509: T462 = 1'h0;
    1510: T462 = 1'h0;
    1511: T462 = 1'h0;
    1512: T462 = 1'h0;
    1513: T462 = 1'h0;
    1514: T462 = 1'h0;
    1515: T462 = 1'h0;
    1516: T462 = 1'h0;
    1517: T462 = 1'h0;
    1518: T462 = 1'h0;
    1519: T462 = 1'h0;
    1520: T462 = 1'h0;
    1521: T462 = 1'h0;
    1522: T462 = 1'h0;
    1523: T462 = 1'h0;
    1524: T462 = 1'h0;
    1525: T462 = 1'h0;
    1526: T462 = 1'h0;
    1527: T462 = 1'h0;
    1528: T462 = 1'h0;
    1529: T462 = 1'h0;
    1530: T462 = 1'h0;
    1531: T462 = 1'h0;
    1532: T462 = 1'h0;
    1533: T462 = 1'h0;
    1534: T462 = 1'h0;
    1535: T462 = 1'h0;
    1536: T462 = 1'h0;
    1537: T462 = 1'h0;
    1538: T462 = 1'h0;
    1539: T462 = 1'h0;
    1540: T462 = 1'h0;
    1541: T462 = 1'h0;
    1542: T462 = 1'h0;
    1543: T462 = 1'h0;
    1544: T462 = 1'h0;
    1545: T462 = 1'h0;
    1546: T462 = 1'h0;
    1547: T462 = 1'h0;
    1548: T462 = 1'h0;
    1549: T462 = 1'h0;
    1550: T462 = 1'h0;
    1551: T462 = 1'h0;
    1552: T462 = 1'h0;
    1553: T462 = 1'h0;
    1554: T462 = 1'h0;
    1555: T462 = 1'h0;
    1556: T462 = 1'h0;
    1557: T462 = 1'h0;
    1558: T462 = 1'h0;
    1559: T462 = 1'h0;
    1560: T462 = 1'h0;
    1561: T462 = 1'h0;
    1562: T462 = 1'h0;
    1563: T462 = 1'h0;
    1564: T462 = 1'h0;
    1565: T462 = 1'h0;
    1566: T462 = 1'h0;
    1567: T462 = 1'h0;
    1568: T462 = 1'h0;
    1569: T462 = 1'h0;
    1570: T462 = 1'h0;
    1571: T462 = 1'h0;
    1572: T462 = 1'h0;
    1573: T462 = 1'h0;
    1574: T462 = 1'h0;
    1575: T462 = 1'h0;
    1576: T462 = 1'h0;
    1577: T462 = 1'h0;
    1578: T462 = 1'h0;
    1579: T462 = 1'h0;
    1580: T462 = 1'h0;
    1581: T462 = 1'h0;
    1582: T462 = 1'h0;
    1583: T462 = 1'h0;
    1584: T462 = 1'h0;
    1585: T462 = 1'h0;
    1586: T462 = 1'h0;
    1587: T462 = 1'h0;
    1588: T462 = 1'h0;
    1589: T462 = 1'h0;
    1590: T462 = 1'h0;
    1591: T462 = 1'h0;
    1592: T462 = 1'h0;
    1593: T462 = 1'h0;
    1594: T462 = 1'h0;
    1595: T462 = 1'h0;
    1596: T462 = 1'h0;
    1597: T462 = 1'h0;
    1598: T462 = 1'h0;
    1599: T462 = 1'h0;
    1600: T462 = 1'h0;
    1601: T462 = 1'h0;
    1602: T462 = 1'h0;
    1603: T462 = 1'h0;
    1604: T462 = 1'h0;
    1605: T462 = 1'h0;
    1606: T462 = 1'h0;
    1607: T462 = 1'h0;
    1608: T462 = 1'h0;
    1609: T462 = 1'h0;
    1610: T462 = 1'h0;
    1611: T462 = 1'h0;
    1612: T462 = 1'h0;
    1613: T462 = 1'h0;
    1614: T462 = 1'h0;
    1615: T462 = 1'h0;
    1616: T462 = 1'h0;
    1617: T462 = 1'h0;
    1618: T462 = 1'h0;
    1619: T462 = 1'h0;
    1620: T462 = 1'h0;
    1621: T462 = 1'h0;
    1622: T462 = 1'h0;
    1623: T462 = 1'h0;
    1624: T462 = 1'h0;
    1625: T462 = 1'h0;
    1626: T462 = 1'h0;
    1627: T462 = 1'h0;
    1628: T462 = 1'h0;
    1629: T462 = 1'h0;
    1630: T462 = 1'h0;
    1631: T462 = 1'h0;
    1632: T462 = 1'h0;
    1633: T462 = 1'h0;
    1634: T462 = 1'h0;
    1635: T462 = 1'h0;
    1636: T462 = 1'h0;
    1637: T462 = 1'h0;
    1638: T462 = 1'h0;
    1639: T462 = 1'h0;
    1640: T462 = 1'h0;
    1641: T462 = 1'h0;
    1642: T462 = 1'h0;
    1643: T462 = 1'h0;
    1644: T462 = 1'h0;
    1645: T462 = 1'h0;
    1646: T462 = 1'h0;
    1647: T462 = 1'h0;
    1648: T462 = 1'h0;
    1649: T462 = 1'h0;
    1650: T462 = 1'h0;
    1651: T462 = 1'h0;
    1652: T462 = 1'h0;
    1653: T462 = 1'h0;
    1654: T462 = 1'h0;
    1655: T462 = 1'h0;
    1656: T462 = 1'h0;
    1657: T462 = 1'h0;
    1658: T462 = 1'h0;
    1659: T462 = 1'h0;
    1660: T462 = 1'h0;
    1661: T462 = 1'h0;
    1662: T462 = 1'h0;
    1663: T462 = 1'h0;
    1664: T462 = 1'h0;
    1665: T462 = 1'h0;
    1666: T462 = 1'h0;
    1667: T462 = 1'h0;
    1668: T462 = 1'h0;
    1669: T462 = 1'h0;
    1670: T462 = 1'h0;
    1671: T462 = 1'h0;
    1672: T462 = 1'h0;
    1673: T462 = 1'h0;
    1674: T462 = 1'h0;
    1675: T462 = 1'h0;
    1676: T462 = 1'h0;
    1677: T462 = 1'h0;
    1678: T462 = 1'h0;
    1679: T462 = 1'h0;
    1680: T462 = 1'h0;
    1681: T462 = 1'h0;
    1682: T462 = 1'h0;
    1683: T462 = 1'h0;
    1684: T462 = 1'h0;
    1685: T462 = 1'h0;
    1686: T462 = 1'h0;
    1687: T462 = 1'h0;
    1688: T462 = 1'h0;
    1689: T462 = 1'h0;
    1690: T462 = 1'h0;
    1691: T462 = 1'h0;
    1692: T462 = 1'h0;
    1693: T462 = 1'h0;
    1694: T462 = 1'h0;
    1695: T462 = 1'h0;
    1696: T462 = 1'h0;
    1697: T462 = 1'h0;
    1698: T462 = 1'h0;
    1699: T462 = 1'h0;
    1700: T462 = 1'h0;
    1701: T462 = 1'h0;
    1702: T462 = 1'h0;
    1703: T462 = 1'h0;
    1704: T462 = 1'h0;
    1705: T462 = 1'h0;
    1706: T462 = 1'h0;
    1707: T462 = 1'h0;
    1708: T462 = 1'h0;
    1709: T462 = 1'h0;
    1710: T462 = 1'h0;
    1711: T462 = 1'h0;
    1712: T462 = 1'h0;
    1713: T462 = 1'h0;
    1714: T462 = 1'h0;
    1715: T462 = 1'h0;
    1716: T462 = 1'h0;
    1717: T462 = 1'h0;
    1718: T462 = 1'h0;
    1719: T462 = 1'h0;
    1720: T462 = 1'h0;
    1721: T462 = 1'h0;
    1722: T462 = 1'h0;
    1723: T462 = 1'h0;
    1724: T462 = 1'h0;
    1725: T462 = 1'h0;
    1726: T462 = 1'h0;
    1727: T462 = 1'h0;
    1728: T462 = 1'h0;
    1729: T462 = 1'h0;
    1730: T462 = 1'h0;
    1731: T462 = 1'h0;
    1732: T462 = 1'h0;
    1733: T462 = 1'h0;
    1734: T462 = 1'h0;
    1735: T462 = 1'h0;
    1736: T462 = 1'h0;
    1737: T462 = 1'h0;
    1738: T462 = 1'h0;
    1739: T462 = 1'h0;
    1740: T462 = 1'h0;
    1741: T462 = 1'h0;
    1742: T462 = 1'h0;
    1743: T462 = 1'h0;
    1744: T462 = 1'h0;
    1745: T462 = 1'h0;
    1746: T462 = 1'h0;
    1747: T462 = 1'h0;
    1748: T462 = 1'h0;
    1749: T462 = 1'h0;
    1750: T462 = 1'h0;
    1751: T462 = 1'h0;
    1752: T462 = 1'h0;
    1753: T462 = 1'h0;
    1754: T462 = 1'h0;
    1755: T462 = 1'h0;
    1756: T462 = 1'h0;
    1757: T462 = 1'h0;
    1758: T462 = 1'h0;
    1759: T462 = 1'h0;
    1760: T462 = 1'h0;
    1761: T462 = 1'h0;
    1762: T462 = 1'h0;
    1763: T462 = 1'h0;
    1764: T462 = 1'h0;
    1765: T462 = 1'h0;
    1766: T462 = 1'h0;
    1767: T462 = 1'h0;
    1768: T462 = 1'h0;
    1769: T462 = 1'h0;
    1770: T462 = 1'h0;
    1771: T462 = 1'h0;
    1772: T462 = 1'h0;
    1773: T462 = 1'h0;
    1774: T462 = 1'h0;
    1775: T462 = 1'h0;
    1776: T462 = 1'h0;
    1777: T462 = 1'h0;
    1778: T462 = 1'h0;
    1779: T462 = 1'h0;
    1780: T462 = 1'h0;
    1781: T462 = 1'h0;
    1782: T462 = 1'h0;
    1783: T462 = 1'h0;
    1784: T462 = 1'h0;
    1785: T462 = 1'h0;
    1786: T462 = 1'h0;
    1787: T462 = 1'h0;
    1788: T462 = 1'h0;
    1789: T462 = 1'h0;
    1790: T462 = 1'h0;
    1791: T462 = 1'h0;
    1792: T462 = 1'h0;
    1793: T462 = 1'h0;
    1794: T462 = 1'h0;
    1795: T462 = 1'h0;
    1796: T462 = 1'h0;
    1797: T462 = 1'h0;
    1798: T462 = 1'h0;
    1799: T462 = 1'h0;
    1800: T462 = 1'h0;
    1801: T462 = 1'h0;
    1802: T462 = 1'h0;
    1803: T462 = 1'h0;
    1804: T462 = 1'h0;
    1805: T462 = 1'h0;
    1806: T462 = 1'h0;
    1807: T462 = 1'h0;
    1808: T462 = 1'h0;
    1809: T462 = 1'h0;
    1810: T462 = 1'h0;
    1811: T462 = 1'h0;
    1812: T462 = 1'h0;
    1813: T462 = 1'h0;
    1814: T462 = 1'h0;
    1815: T462 = 1'h0;
    1816: T462 = 1'h0;
    1817: T462 = 1'h0;
    1818: T462 = 1'h0;
    1819: T462 = 1'h0;
    1820: T462 = 1'h0;
    1821: T462 = 1'h0;
    1822: T462 = 1'h0;
    1823: T462 = 1'h0;
    1824: T462 = 1'h0;
    1825: T462 = 1'h0;
    1826: T462 = 1'h0;
    1827: T462 = 1'h0;
    1828: T462 = 1'h0;
    1829: T462 = 1'h0;
    1830: T462 = 1'h0;
    1831: T462 = 1'h0;
    1832: T462 = 1'h0;
    1833: T462 = 1'h0;
    1834: T462 = 1'h0;
    1835: T462 = 1'h0;
    1836: T462 = 1'h0;
    1837: T462 = 1'h0;
    1838: T462 = 1'h0;
    1839: T462 = 1'h0;
    1840: T462 = 1'h0;
    1841: T462 = 1'h0;
    1842: T462 = 1'h0;
    1843: T462 = 1'h0;
    1844: T462 = 1'h0;
    1845: T462 = 1'h0;
    1846: T462 = 1'h0;
    1847: T462 = 1'h0;
    1848: T462 = 1'h0;
    1849: T462 = 1'h0;
    1850: T462 = 1'h0;
    1851: T462 = 1'h0;
    1852: T462 = 1'h0;
    1853: T462 = 1'h0;
    1854: T462 = 1'h0;
    1855: T462 = 1'h0;
    1856: T462 = 1'h0;
    1857: T462 = 1'h0;
    1858: T462 = 1'h0;
    1859: T462 = 1'h0;
    1860: T462 = 1'h0;
    1861: T462 = 1'h0;
    1862: T462 = 1'h0;
    1863: T462 = 1'h0;
    1864: T462 = 1'h0;
    1865: T462 = 1'h0;
    1866: T462 = 1'h0;
    1867: T462 = 1'h0;
    1868: T462 = 1'h0;
    1869: T462 = 1'h0;
    1870: T462 = 1'h0;
    1871: T462 = 1'h0;
    1872: T462 = 1'h0;
    1873: T462 = 1'h0;
    1874: T462 = 1'h0;
    1875: T462 = 1'h0;
    1876: T462 = 1'h0;
    1877: T462 = 1'h0;
    1878: T462 = 1'h0;
    1879: T462 = 1'h0;
    1880: T462 = 1'h0;
    1881: T462 = 1'h0;
    1882: T462 = 1'h0;
    1883: T462 = 1'h0;
    1884: T462 = 1'h0;
    1885: T462 = 1'h0;
    1886: T462 = 1'h0;
    1887: T462 = 1'h0;
    1888: T462 = 1'h0;
    1889: T462 = 1'h0;
    1890: T462 = 1'h0;
    1891: T462 = 1'h0;
    1892: T462 = 1'h0;
    1893: T462 = 1'h0;
    1894: T462 = 1'h0;
    1895: T462 = 1'h0;
    1896: T462 = 1'h0;
    1897: T462 = 1'h0;
    1898: T462 = 1'h0;
    1899: T462 = 1'h0;
    1900: T462 = 1'h0;
    1901: T462 = 1'h0;
    1902: T462 = 1'h0;
    1903: T462 = 1'h0;
    1904: T462 = 1'h0;
    1905: T462 = 1'h0;
    1906: T462 = 1'h0;
    1907: T462 = 1'h0;
    1908: T462 = 1'h0;
    1909: T462 = 1'h0;
    1910: T462 = 1'h0;
    1911: T462 = 1'h0;
    1912: T462 = 1'h0;
    1913: T462 = 1'h0;
    1914: T462 = 1'h0;
    1915: T462 = 1'h0;
    1916: T462 = 1'h0;
    1917: T462 = 1'h0;
    1918: T462 = 1'h0;
    1919: T462 = 1'h0;
    1920: T462 = 1'h0;
    1921: T462 = 1'h0;
    1922: T462 = 1'h0;
    1923: T462 = 1'h0;
    1924: T462 = 1'h0;
    1925: T462 = 1'h0;
    1926: T462 = 1'h0;
    1927: T462 = 1'h0;
    1928: T462 = 1'h0;
    1929: T462 = 1'h0;
    1930: T462 = 1'h0;
    1931: T462 = 1'h0;
    1932: T462 = 1'h0;
    1933: T462 = 1'h0;
    1934: T462 = 1'h0;
    1935: T462 = 1'h0;
    1936: T462 = 1'h0;
    1937: T462 = 1'h0;
    1938: T462 = 1'h0;
    1939: T462 = 1'h0;
    1940: T462 = 1'h0;
    1941: T462 = 1'h0;
    1942: T462 = 1'h0;
    1943: T462 = 1'h0;
    1944: T462 = 1'h0;
    1945: T462 = 1'h0;
    1946: T462 = 1'h0;
    1947: T462 = 1'h0;
    1948: T462 = 1'h0;
    1949: T462 = 1'h0;
    1950: T462 = 1'h0;
    1951: T462 = 1'h0;
    1952: T462 = 1'h0;
    1953: T462 = 1'h0;
    1954: T462 = 1'h0;
    1955: T462 = 1'h0;
    1956: T462 = 1'h0;
    1957: T462 = 1'h0;
    1958: T462 = 1'h0;
    1959: T462 = 1'h0;
    1960: T462 = 1'h0;
    1961: T462 = 1'h0;
    1962: T462 = 1'h0;
    1963: T462 = 1'h0;
    1964: T462 = 1'h0;
    1965: T462 = 1'h0;
    1966: T462 = 1'h0;
    1967: T462 = 1'h0;
    1968: T462 = 1'h0;
    1969: T462 = 1'h0;
    1970: T462 = 1'h0;
    1971: T462 = 1'h0;
    1972: T462 = 1'h0;
    1973: T462 = 1'h0;
    1974: T462 = 1'h0;
    1975: T462 = 1'h0;
    1976: T462 = 1'h0;
    1977: T462 = 1'h0;
    1978: T462 = 1'h0;
    1979: T462 = 1'h0;
    1980: T462 = 1'h0;
    1981: T462 = 1'h0;
    1982: T462 = 1'h0;
    1983: T462 = 1'h0;
    1984: T462 = 1'h0;
    1985: T462 = 1'h0;
    1986: T462 = 1'h0;
    1987: T462 = 1'h0;
    1988: T462 = 1'h0;
    1989: T462 = 1'h0;
    1990: T462 = 1'h0;
    1991: T462 = 1'h0;
    1992: T462 = 1'h0;
    1993: T462 = 1'h0;
    1994: T462 = 1'h0;
    1995: T462 = 1'h0;
    1996: T462 = 1'h0;
    1997: T462 = 1'h0;
    1998: T462 = 1'h0;
    1999: T462 = 1'h0;
    2000: T462 = 1'h0;
    2001: T462 = 1'h0;
    2002: T462 = 1'h0;
    2003: T462 = 1'h0;
    2004: T462 = 1'h0;
    2005: T462 = 1'h0;
    2006: T462 = 1'h0;
    2007: T462 = 1'h0;
    2008: T462 = 1'h0;
    2009: T462 = 1'h0;
    2010: T462 = 1'h0;
    2011: T462 = 1'h0;
    2012: T462 = 1'h0;
    2013: T462 = 1'h0;
    2014: T462 = 1'h0;
    2015: T462 = 1'h0;
    2016: T462 = 1'h0;
    2017: T462 = 1'h0;
    2018: T462 = 1'h0;
    2019: T462 = 1'h0;
    2020: T462 = 1'h0;
    2021: T462 = 1'h0;
    2022: T462 = 1'h0;
    2023: T462 = 1'h0;
    2024: T462 = 1'h0;
    2025: T462 = 1'h0;
    2026: T462 = 1'h0;
    2027: T462 = 1'h0;
    2028: T462 = 1'h0;
    2029: T462 = 1'h0;
    2030: T462 = 1'h0;
    2031: T462 = 1'h0;
    2032: T462 = 1'h0;
    2033: T462 = 1'h0;
    2034: T462 = 1'h0;
    2035: T462 = 1'h0;
    2036: T462 = 1'h0;
    2037: T462 = 1'h0;
    2038: T462 = 1'h0;
    2039: T462 = 1'h0;
    2040: T462 = 1'h0;
    2041: T462 = 1'h0;
    2042: T462 = 1'h0;
    2043: T462 = 1'h0;
    2044: T462 = 1'h0;
    2045: T462 = 1'h0;
    2046: T462 = 1'h0;
    2047: T462 = 1'h0;
    2048: T462 = 1'h0;
    2049: T462 = 1'h0;
    2050: T462 = 1'h0;
    2051: T462 = 1'h0;
    2052: T462 = 1'h0;
    2053: T462 = 1'h0;
    2054: T462 = 1'h0;
    2055: T462 = 1'h0;
    2056: T462 = 1'h0;
    2057: T462 = 1'h0;
    2058: T462 = 1'h0;
    2059: T462 = 1'h0;
    2060: T462 = 1'h0;
    2061: T462 = 1'h0;
    2062: T462 = 1'h0;
    2063: T462 = 1'h0;
    2064: T462 = 1'h0;
    2065: T462 = 1'h0;
    2066: T462 = 1'h0;
    2067: T462 = 1'h0;
    2068: T462 = 1'h0;
    2069: T462 = 1'h0;
    2070: T462 = 1'h0;
    2071: T462 = 1'h0;
    2072: T462 = 1'h0;
    2073: T462 = 1'h0;
    2074: T462 = 1'h0;
    2075: T462 = 1'h0;
    2076: T462 = 1'h0;
    2077: T462 = 1'h0;
    2078: T462 = 1'h0;
    2079: T462 = 1'h0;
    2080: T462 = 1'h0;
    2081: T462 = 1'h0;
    2082: T462 = 1'h0;
    2083: T462 = 1'h0;
    2084: T462 = 1'h0;
    2085: T462 = 1'h0;
    2086: T462 = 1'h0;
    2087: T462 = 1'h0;
    2088: T462 = 1'h0;
    2089: T462 = 1'h0;
    2090: T462 = 1'h0;
    2091: T462 = 1'h0;
    2092: T462 = 1'h0;
    2093: T462 = 1'h0;
    2094: T462 = 1'h0;
    2095: T462 = 1'h0;
    2096: T462 = 1'h0;
    2097: T462 = 1'h0;
    2098: T462 = 1'h0;
    2099: T462 = 1'h0;
    2100: T462 = 1'h0;
    2101: T462 = 1'h0;
    2102: T462 = 1'h0;
    2103: T462 = 1'h0;
    2104: T462 = 1'h0;
    2105: T462 = 1'h0;
    2106: T462 = 1'h0;
    2107: T462 = 1'h0;
    2108: T462 = 1'h0;
    2109: T462 = 1'h0;
    2110: T462 = 1'h0;
    2111: T462 = 1'h0;
    2112: T462 = 1'h0;
    2113: T462 = 1'h0;
    2114: T462 = 1'h0;
    2115: T462 = 1'h0;
    2116: T462 = 1'h0;
    2117: T462 = 1'h0;
    2118: T462 = 1'h0;
    2119: T462 = 1'h0;
    2120: T462 = 1'h0;
    2121: T462 = 1'h0;
    2122: T462 = 1'h0;
    2123: T462 = 1'h0;
    2124: T462 = 1'h0;
    2125: T462 = 1'h0;
    2126: T462 = 1'h0;
    2127: T462 = 1'h0;
    2128: T462 = 1'h0;
    2129: T462 = 1'h0;
    2130: T462 = 1'h0;
    2131: T462 = 1'h0;
    2132: T462 = 1'h0;
    2133: T462 = 1'h0;
    2134: T462 = 1'h0;
    2135: T462 = 1'h0;
    2136: T462 = 1'h0;
    2137: T462 = 1'h0;
    2138: T462 = 1'h0;
    2139: T462 = 1'h0;
    2140: T462 = 1'h0;
    2141: T462 = 1'h0;
    2142: T462 = 1'h0;
    2143: T462 = 1'h0;
    2144: T462 = 1'h0;
    2145: T462 = 1'h0;
    2146: T462 = 1'h0;
    2147: T462 = 1'h0;
    2148: T462 = 1'h0;
    2149: T462 = 1'h0;
    2150: T462 = 1'h0;
    2151: T462 = 1'h0;
    2152: T462 = 1'h0;
    2153: T462 = 1'h0;
    2154: T462 = 1'h0;
    2155: T462 = 1'h0;
    2156: T462 = 1'h0;
    2157: T462 = 1'h0;
    2158: T462 = 1'h0;
    2159: T462 = 1'h0;
    2160: T462 = 1'h0;
    2161: T462 = 1'h0;
    2162: T462 = 1'h0;
    2163: T462 = 1'h0;
    2164: T462 = 1'h0;
    2165: T462 = 1'h0;
    2166: T462 = 1'h0;
    2167: T462 = 1'h0;
    2168: T462 = 1'h0;
    2169: T462 = 1'h0;
    2170: T462 = 1'h0;
    2171: T462 = 1'h0;
    2172: T462 = 1'h0;
    2173: T462 = 1'h0;
    2174: T462 = 1'h0;
    2175: T462 = 1'h0;
    2176: T462 = 1'h0;
    2177: T462 = 1'h0;
    2178: T462 = 1'h0;
    2179: T462 = 1'h0;
    2180: T462 = 1'h0;
    2181: T462 = 1'h0;
    2182: T462 = 1'h0;
    2183: T462 = 1'h0;
    2184: T462 = 1'h0;
    2185: T462 = 1'h0;
    2186: T462 = 1'h0;
    2187: T462 = 1'h0;
    2188: T462 = 1'h0;
    2189: T462 = 1'h0;
    2190: T462 = 1'h0;
    2191: T462 = 1'h0;
    2192: T462 = 1'h0;
    2193: T462 = 1'h0;
    2194: T462 = 1'h0;
    2195: T462 = 1'h0;
    2196: T462 = 1'h0;
    2197: T462 = 1'h0;
    2198: T462 = 1'h0;
    2199: T462 = 1'h0;
    2200: T462 = 1'h0;
    2201: T462 = 1'h0;
    2202: T462 = 1'h0;
    2203: T462 = 1'h0;
    2204: T462 = 1'h0;
    2205: T462 = 1'h0;
    2206: T462 = 1'h0;
    2207: T462 = 1'h0;
    2208: T462 = 1'h0;
    2209: T462 = 1'h0;
    2210: T462 = 1'h0;
    2211: T462 = 1'h0;
    2212: T462 = 1'h0;
    2213: T462 = 1'h0;
    2214: T462 = 1'h0;
    2215: T462 = 1'h0;
    2216: T462 = 1'h0;
    2217: T462 = 1'h0;
    2218: T462 = 1'h0;
    2219: T462 = 1'h0;
    2220: T462 = 1'h0;
    2221: T462 = 1'h0;
    2222: T462 = 1'h0;
    2223: T462 = 1'h0;
    2224: T462 = 1'h0;
    2225: T462 = 1'h0;
    2226: T462 = 1'h0;
    2227: T462 = 1'h0;
    2228: T462 = 1'h0;
    2229: T462 = 1'h0;
    2230: T462 = 1'h0;
    2231: T462 = 1'h0;
    2232: T462 = 1'h0;
    2233: T462 = 1'h0;
    2234: T462 = 1'h0;
    2235: T462 = 1'h0;
    2236: T462 = 1'h0;
    2237: T462 = 1'h0;
    2238: T462 = 1'h0;
    2239: T462 = 1'h0;
    2240: T462 = 1'h0;
    2241: T462 = 1'h0;
    2242: T462 = 1'h0;
    2243: T462 = 1'h0;
    2244: T462 = 1'h0;
    2245: T462 = 1'h0;
    2246: T462 = 1'h0;
    2247: T462 = 1'h0;
    2248: T462 = 1'h0;
    2249: T462 = 1'h0;
    2250: T462 = 1'h0;
    2251: T462 = 1'h0;
    2252: T462 = 1'h0;
    2253: T462 = 1'h0;
    2254: T462 = 1'h0;
    2255: T462 = 1'h0;
    2256: T462 = 1'h0;
    2257: T462 = 1'h0;
    2258: T462 = 1'h0;
    2259: T462 = 1'h0;
    2260: T462 = 1'h0;
    2261: T462 = 1'h0;
    2262: T462 = 1'h0;
    2263: T462 = 1'h0;
    2264: T462 = 1'h0;
    2265: T462 = 1'h0;
    2266: T462 = 1'h0;
    2267: T462 = 1'h0;
    2268: T462 = 1'h0;
    2269: T462 = 1'h0;
    2270: T462 = 1'h0;
    2271: T462 = 1'h0;
    2272: T462 = 1'h0;
    2273: T462 = 1'h0;
    2274: T462 = 1'h0;
    2275: T462 = 1'h0;
    2276: T462 = 1'h0;
    2277: T462 = 1'h0;
    2278: T462 = 1'h0;
    2279: T462 = 1'h0;
    2280: T462 = 1'h0;
    2281: T462 = 1'h0;
    2282: T462 = 1'h0;
    2283: T462 = 1'h0;
    2284: T462 = 1'h0;
    2285: T462 = 1'h0;
    2286: T462 = 1'h0;
    2287: T462 = 1'h0;
    2288: T462 = 1'h0;
    2289: T462 = 1'h0;
    2290: T462 = 1'h0;
    2291: T462 = 1'h0;
    2292: T462 = 1'h0;
    2293: T462 = 1'h0;
    2294: T462 = 1'h0;
    2295: T462 = 1'h0;
    2296: T462 = 1'h0;
    2297: T462 = 1'h0;
    2298: T462 = 1'h0;
    2299: T462 = 1'h0;
    2300: T462 = 1'h0;
    2301: T462 = 1'h0;
    2302: T462 = 1'h0;
    2303: T462 = 1'h0;
    2304: T462 = 1'h0;
    2305: T462 = 1'h0;
    2306: T462 = 1'h0;
    2307: T462 = 1'h0;
    2308: T462 = 1'h0;
    2309: T462 = 1'h0;
    2310: T462 = 1'h0;
    2311: T462 = 1'h0;
    2312: T462 = 1'h0;
    2313: T462 = 1'h0;
    2314: T462 = 1'h0;
    2315: T462 = 1'h0;
    2316: T462 = 1'h0;
    2317: T462 = 1'h0;
    2318: T462 = 1'h0;
    2319: T462 = 1'h0;
    2320: T462 = 1'h0;
    2321: T462 = 1'h0;
    2322: T462 = 1'h0;
    2323: T462 = 1'h0;
    2324: T462 = 1'h0;
    2325: T462 = 1'h0;
    2326: T462 = 1'h0;
    2327: T462 = 1'h0;
    2328: T462 = 1'h0;
    2329: T462 = 1'h0;
    2330: T462 = 1'h0;
    2331: T462 = 1'h0;
    2332: T462 = 1'h0;
    2333: T462 = 1'h0;
    2334: T462 = 1'h0;
    2335: T462 = 1'h0;
    2336: T462 = 1'h0;
    2337: T462 = 1'h0;
    2338: T462 = 1'h0;
    2339: T462 = 1'h0;
    2340: T462 = 1'h0;
    2341: T462 = 1'h0;
    2342: T462 = 1'h0;
    2343: T462 = 1'h0;
    2344: T462 = 1'h0;
    2345: T462 = 1'h0;
    2346: T462 = 1'h0;
    2347: T462 = 1'h0;
    2348: T462 = 1'h0;
    2349: T462 = 1'h0;
    2350: T462 = 1'h0;
    2351: T462 = 1'h0;
    2352: T462 = 1'h0;
    2353: T462 = 1'h0;
    2354: T462 = 1'h0;
    2355: T462 = 1'h0;
    2356: T462 = 1'h0;
    2357: T462 = 1'h0;
    2358: T462 = 1'h0;
    2359: T462 = 1'h0;
    2360: T462 = 1'h0;
    2361: T462 = 1'h0;
    2362: T462 = 1'h0;
    2363: T462 = 1'h0;
    2364: T462 = 1'h0;
    2365: T462 = 1'h0;
    2366: T462 = 1'h0;
    2367: T462 = 1'h0;
    2368: T462 = 1'h0;
    2369: T462 = 1'h0;
    2370: T462 = 1'h0;
    2371: T462 = 1'h0;
    2372: T462 = 1'h0;
    2373: T462 = 1'h0;
    2374: T462 = 1'h0;
    2375: T462 = 1'h0;
    2376: T462 = 1'h0;
    2377: T462 = 1'h0;
    2378: T462 = 1'h0;
    2379: T462 = 1'h0;
    2380: T462 = 1'h0;
    2381: T462 = 1'h0;
    2382: T462 = 1'h0;
    2383: T462 = 1'h0;
    2384: T462 = 1'h0;
    2385: T462 = 1'h0;
    2386: T462 = 1'h0;
    2387: T462 = 1'h0;
    2388: T462 = 1'h0;
    2389: T462 = 1'h0;
    2390: T462 = 1'h0;
    2391: T462 = 1'h0;
    2392: T462 = 1'h0;
    2393: T462 = 1'h0;
    2394: T462 = 1'h0;
    2395: T462 = 1'h0;
    2396: T462 = 1'h0;
    2397: T462 = 1'h0;
    2398: T462 = 1'h0;
    2399: T462 = 1'h0;
    2400: T462 = 1'h0;
    2401: T462 = 1'h0;
    2402: T462 = 1'h0;
    2403: T462 = 1'h0;
    2404: T462 = 1'h0;
    2405: T462 = 1'h0;
    2406: T462 = 1'h0;
    2407: T462 = 1'h0;
    2408: T462 = 1'h0;
    2409: T462 = 1'h0;
    2410: T462 = 1'h0;
    2411: T462 = 1'h0;
    2412: T462 = 1'h0;
    2413: T462 = 1'h0;
    2414: T462 = 1'h0;
    2415: T462 = 1'h0;
    2416: T462 = 1'h0;
    2417: T462 = 1'h0;
    2418: T462 = 1'h0;
    2419: T462 = 1'h0;
    2420: T462 = 1'h0;
    2421: T462 = 1'h0;
    2422: T462 = 1'h0;
    2423: T462 = 1'h0;
    2424: T462 = 1'h0;
    2425: T462 = 1'h0;
    2426: T462 = 1'h0;
    2427: T462 = 1'h0;
    2428: T462 = 1'h0;
    2429: T462 = 1'h0;
    2430: T462 = 1'h0;
    2431: T462 = 1'h0;
    2432: T462 = 1'h0;
    2433: T462 = 1'h0;
    2434: T462 = 1'h0;
    2435: T462 = 1'h0;
    2436: T462 = 1'h0;
    2437: T462 = 1'h0;
    2438: T462 = 1'h0;
    2439: T462 = 1'h0;
    2440: T462 = 1'h0;
    2441: T462 = 1'h0;
    2442: T462 = 1'h0;
    2443: T462 = 1'h0;
    2444: T462 = 1'h0;
    2445: T462 = 1'h0;
    2446: T462 = 1'h0;
    2447: T462 = 1'h0;
    2448: T462 = 1'h0;
    2449: T462 = 1'h0;
    2450: T462 = 1'h0;
    2451: T462 = 1'h0;
    2452: T462 = 1'h0;
    2453: T462 = 1'h0;
    2454: T462 = 1'h0;
    2455: T462 = 1'h0;
    2456: T462 = 1'h0;
    2457: T462 = 1'h0;
    2458: T462 = 1'h0;
    2459: T462 = 1'h0;
    2460: T462 = 1'h0;
    2461: T462 = 1'h0;
    2462: T462 = 1'h0;
    2463: T462 = 1'h0;
    2464: T462 = 1'h0;
    2465: T462 = 1'h0;
    2466: T462 = 1'h0;
    2467: T462 = 1'h0;
    2468: T462 = 1'h0;
    2469: T462 = 1'h0;
    2470: T462 = 1'h0;
    2471: T462 = 1'h0;
    2472: T462 = 1'h0;
    2473: T462 = 1'h0;
    2474: T462 = 1'h0;
    2475: T462 = 1'h0;
    2476: T462 = 1'h0;
    2477: T462 = 1'h0;
    2478: T462 = 1'h0;
    2479: T462 = 1'h0;
    2480: T462 = 1'h0;
    2481: T462 = 1'h0;
    2482: T462 = 1'h0;
    2483: T462 = 1'h0;
    2484: T462 = 1'h0;
    2485: T462 = 1'h0;
    2486: T462 = 1'h0;
    2487: T462 = 1'h0;
    2488: T462 = 1'h0;
    2489: T462 = 1'h0;
    2490: T462 = 1'h0;
    2491: T462 = 1'h0;
    2492: T462 = 1'h0;
    2493: T462 = 1'h0;
    2494: T462 = 1'h0;
    2495: T462 = 1'h0;
    2496: T462 = 1'h0;
    2497: T462 = 1'h0;
    2498: T462 = 1'h0;
    2499: T462 = 1'h0;
    2500: T462 = 1'h0;
    2501: T462 = 1'h0;
    2502: T462 = 1'h0;
    2503: T462 = 1'h0;
    2504: T462 = 1'h0;
    2505: T462 = 1'h0;
    2506: T462 = 1'h0;
    2507: T462 = 1'h0;
    2508: T462 = 1'h0;
    2509: T462 = 1'h0;
    2510: T462 = 1'h0;
    2511: T462 = 1'h0;
    2512: T462 = 1'h0;
    2513: T462 = 1'h0;
    2514: T462 = 1'h0;
    2515: T462 = 1'h0;
    2516: T462 = 1'h0;
    2517: T462 = 1'h0;
    2518: T462 = 1'h0;
    2519: T462 = 1'h0;
    2520: T462 = 1'h0;
    2521: T462 = 1'h0;
    2522: T462 = 1'h0;
    2523: T462 = 1'h0;
    2524: T462 = 1'h0;
    2525: T462 = 1'h0;
    2526: T462 = 1'h0;
    2527: T462 = 1'h0;
    2528: T462 = 1'h0;
    2529: T462 = 1'h0;
    2530: T462 = 1'h0;
    2531: T462 = 1'h0;
    2532: T462 = 1'h0;
    2533: T462 = 1'h0;
    2534: T462 = 1'h0;
    2535: T462 = 1'h0;
    2536: T462 = 1'h0;
    2537: T462 = 1'h0;
    2538: T462 = 1'h0;
    2539: T462 = 1'h0;
    2540: T462 = 1'h0;
    2541: T462 = 1'h0;
    2542: T462 = 1'h0;
    2543: T462 = 1'h0;
    2544: T462 = 1'h0;
    2545: T462 = 1'h0;
    2546: T462 = 1'h0;
    2547: T462 = 1'h0;
    2548: T462 = 1'h0;
    2549: T462 = 1'h0;
    2550: T462 = 1'h0;
    2551: T462 = 1'h0;
    2552: T462 = 1'h0;
    2553: T462 = 1'h0;
    2554: T462 = 1'h0;
    2555: T462 = 1'h0;
    2556: T462 = 1'h0;
    2557: T462 = 1'h0;
    2558: T462 = 1'h0;
    2559: T462 = 1'h0;
    2560: T462 = 1'h0;
    2561: T462 = 1'h0;
    2562: T462 = 1'h0;
    2563: T462 = 1'h0;
    2564: T462 = 1'h0;
    2565: T462 = 1'h0;
    2566: T462 = 1'h0;
    2567: T462 = 1'h0;
    2568: T462 = 1'h0;
    2569: T462 = 1'h0;
    2570: T462 = 1'h0;
    2571: T462 = 1'h0;
    2572: T462 = 1'h0;
    2573: T462 = 1'h0;
    2574: T462 = 1'h0;
    2575: T462 = 1'h0;
    2576: T462 = 1'h0;
    2577: T462 = 1'h0;
    2578: T462 = 1'h0;
    2579: T462 = 1'h0;
    2580: T462 = 1'h0;
    2581: T462 = 1'h0;
    2582: T462 = 1'h0;
    2583: T462 = 1'h0;
    2584: T462 = 1'h0;
    2585: T462 = 1'h0;
    2586: T462 = 1'h0;
    2587: T462 = 1'h0;
    2588: T462 = 1'h0;
    2589: T462 = 1'h0;
    2590: T462 = 1'h0;
    2591: T462 = 1'h0;
    2592: T462 = 1'h0;
    2593: T462 = 1'h0;
    2594: T462 = 1'h0;
    2595: T462 = 1'h0;
    2596: T462 = 1'h0;
    2597: T462 = 1'h0;
    2598: T462 = 1'h0;
    2599: T462 = 1'h0;
    2600: T462 = 1'h0;
    2601: T462 = 1'h0;
    2602: T462 = 1'h0;
    2603: T462 = 1'h0;
    2604: T462 = 1'h0;
    2605: T462 = 1'h0;
    2606: T462 = 1'h0;
    2607: T462 = 1'h0;
    2608: T462 = 1'h0;
    2609: T462 = 1'h0;
    2610: T462 = 1'h0;
    2611: T462 = 1'h0;
    2612: T462 = 1'h0;
    2613: T462 = 1'h0;
    2614: T462 = 1'h0;
    2615: T462 = 1'h0;
    2616: T462 = 1'h0;
    2617: T462 = 1'h0;
    2618: T462 = 1'h0;
    2619: T462 = 1'h0;
    2620: T462 = 1'h0;
    2621: T462 = 1'h0;
    2622: T462 = 1'h0;
    2623: T462 = 1'h0;
    2624: T462 = 1'h0;
    2625: T462 = 1'h0;
    2626: T462 = 1'h0;
    2627: T462 = 1'h0;
    2628: T462 = 1'h0;
    2629: T462 = 1'h0;
    2630: T462 = 1'h0;
    2631: T462 = 1'h0;
    2632: T462 = 1'h0;
    2633: T462 = 1'h0;
    2634: T462 = 1'h0;
    2635: T462 = 1'h0;
    2636: T462 = 1'h0;
    2637: T462 = 1'h0;
    2638: T462 = 1'h0;
    2639: T462 = 1'h0;
    2640: T462 = 1'h0;
    2641: T462 = 1'h0;
    2642: T462 = 1'h0;
    2643: T462 = 1'h0;
    2644: T462 = 1'h0;
    2645: T462 = 1'h0;
    2646: T462 = 1'h0;
    2647: T462 = 1'h0;
    2648: T462 = 1'h0;
    2649: T462 = 1'h0;
    2650: T462 = 1'h0;
    2651: T462 = 1'h0;
    2652: T462 = 1'h0;
    2653: T462 = 1'h0;
    2654: T462 = 1'h0;
    2655: T462 = 1'h0;
    2656: T462 = 1'h0;
    2657: T462 = 1'h0;
    2658: T462 = 1'h0;
    2659: T462 = 1'h0;
    2660: T462 = 1'h0;
    2661: T462 = 1'h0;
    2662: T462 = 1'h0;
    2663: T462 = 1'h0;
    2664: T462 = 1'h0;
    2665: T462 = 1'h0;
    2666: T462 = 1'h0;
    2667: T462 = 1'h0;
    2668: T462 = 1'h0;
    2669: T462 = 1'h0;
    2670: T462 = 1'h0;
    2671: T462 = 1'h0;
    2672: T462 = 1'h0;
    2673: T462 = 1'h0;
    2674: T462 = 1'h0;
    2675: T462 = 1'h0;
    2676: T462 = 1'h0;
    2677: T462 = 1'h0;
    2678: T462 = 1'h0;
    2679: T462 = 1'h0;
    2680: T462 = 1'h0;
    2681: T462 = 1'h0;
    2682: T462 = 1'h0;
    2683: T462 = 1'h0;
    2684: T462 = 1'h0;
    2685: T462 = 1'h0;
    2686: T462 = 1'h0;
    2687: T462 = 1'h0;
    2688: T462 = 1'h0;
    2689: T462 = 1'h0;
    2690: T462 = 1'h0;
    2691: T462 = 1'h0;
    2692: T462 = 1'h0;
    2693: T462 = 1'h0;
    2694: T462 = 1'h0;
    2695: T462 = 1'h0;
    2696: T462 = 1'h0;
    2697: T462 = 1'h0;
    2698: T462 = 1'h0;
    2699: T462 = 1'h0;
    2700: T462 = 1'h0;
    2701: T462 = 1'h0;
    2702: T462 = 1'h0;
    2703: T462 = 1'h0;
    2704: T462 = 1'h0;
    2705: T462 = 1'h0;
    2706: T462 = 1'h0;
    2707: T462 = 1'h0;
    2708: T462 = 1'h0;
    2709: T462 = 1'h0;
    2710: T462 = 1'h0;
    2711: T462 = 1'h0;
    2712: T462 = 1'h0;
    2713: T462 = 1'h0;
    2714: T462 = 1'h0;
    2715: T462 = 1'h0;
    2716: T462 = 1'h0;
    2717: T462 = 1'h0;
    2718: T462 = 1'h0;
    2719: T462 = 1'h0;
    2720: T462 = 1'h0;
    2721: T462 = 1'h0;
    2722: T462 = 1'h0;
    2723: T462 = 1'h0;
    2724: T462 = 1'h0;
    2725: T462 = 1'h0;
    2726: T462 = 1'h0;
    2727: T462 = 1'h0;
    2728: T462 = 1'h0;
    2729: T462 = 1'h0;
    2730: T462 = 1'h0;
    2731: T462 = 1'h0;
    2732: T462 = 1'h0;
    2733: T462 = 1'h0;
    2734: T462 = 1'h0;
    2735: T462 = 1'h0;
    2736: T462 = 1'h0;
    2737: T462 = 1'h0;
    2738: T462 = 1'h0;
    2739: T462 = 1'h0;
    2740: T462 = 1'h0;
    2741: T462 = 1'h0;
    2742: T462 = 1'h0;
    2743: T462 = 1'h0;
    2744: T462 = 1'h0;
    2745: T462 = 1'h0;
    2746: T462 = 1'h0;
    2747: T462 = 1'h0;
    2748: T462 = 1'h0;
    2749: T462 = 1'h0;
    2750: T462 = 1'h0;
    2751: T462 = 1'h0;
    2752: T462 = 1'h0;
    2753: T462 = 1'h0;
    2754: T462 = 1'h0;
    2755: T462 = 1'h0;
    2756: T462 = 1'h0;
    2757: T462 = 1'h0;
    2758: T462 = 1'h0;
    2759: T462 = 1'h0;
    2760: T462 = 1'h0;
    2761: T462 = 1'h0;
    2762: T462 = 1'h0;
    2763: T462 = 1'h0;
    2764: T462 = 1'h0;
    2765: T462 = 1'h0;
    2766: T462 = 1'h0;
    2767: T462 = 1'h0;
    2768: T462 = 1'h0;
    2769: T462 = 1'h0;
    2770: T462 = 1'h0;
    2771: T462 = 1'h0;
    2772: T462 = 1'h0;
    2773: T462 = 1'h0;
    2774: T462 = 1'h0;
    2775: T462 = 1'h0;
    2776: T462 = 1'h0;
    2777: T462 = 1'h0;
    2778: T462 = 1'h0;
    2779: T462 = 1'h0;
    2780: T462 = 1'h0;
    2781: T462 = 1'h0;
    2782: T462 = 1'h0;
    2783: T462 = 1'h0;
    2784: T462 = 1'h0;
    2785: T462 = 1'h0;
    2786: T462 = 1'h0;
    2787: T462 = 1'h0;
    2788: T462 = 1'h0;
    2789: T462 = 1'h0;
    2790: T462 = 1'h0;
    2791: T462 = 1'h0;
    2792: T462 = 1'h0;
    2793: T462 = 1'h0;
    2794: T462 = 1'h0;
    2795: T462 = 1'h0;
    2796: T462 = 1'h0;
    2797: T462 = 1'h0;
    2798: T462 = 1'h0;
    2799: T462 = 1'h0;
    2800: T462 = 1'h0;
    2801: T462 = 1'h0;
    2802: T462 = 1'h0;
    2803: T462 = 1'h0;
    2804: T462 = 1'h0;
    2805: T462 = 1'h0;
    2806: T462 = 1'h0;
    2807: T462 = 1'h0;
    2808: T462 = 1'h0;
    2809: T462 = 1'h0;
    2810: T462 = 1'h0;
    2811: T462 = 1'h0;
    2812: T462 = 1'h0;
    2813: T462 = 1'h0;
    2814: T462 = 1'h0;
    2815: T462 = 1'h0;
    2816: T462 = 1'h0;
    2817: T462 = 1'h0;
    2818: T462 = 1'h0;
    2819: T462 = 1'h0;
    2820: T462 = 1'h0;
    2821: T462 = 1'h0;
    2822: T462 = 1'h0;
    2823: T462 = 1'h0;
    2824: T462 = 1'h0;
    2825: T462 = 1'h0;
    2826: T462 = 1'h0;
    2827: T462 = 1'h0;
    2828: T462 = 1'h0;
    2829: T462 = 1'h0;
    2830: T462 = 1'h0;
    2831: T462 = 1'h0;
    2832: T462 = 1'h0;
    2833: T462 = 1'h0;
    2834: T462 = 1'h0;
    2835: T462 = 1'h0;
    2836: T462 = 1'h0;
    2837: T462 = 1'h0;
    2838: T462 = 1'h0;
    2839: T462 = 1'h0;
    2840: T462 = 1'h0;
    2841: T462 = 1'h0;
    2842: T462 = 1'h0;
    2843: T462 = 1'h0;
    2844: T462 = 1'h0;
    2845: T462 = 1'h0;
    2846: T462 = 1'h0;
    2847: T462 = 1'h0;
    2848: T462 = 1'h0;
    2849: T462 = 1'h0;
    2850: T462 = 1'h0;
    2851: T462 = 1'h0;
    2852: T462 = 1'h0;
    2853: T462 = 1'h0;
    2854: T462 = 1'h0;
    2855: T462 = 1'h0;
    2856: T462 = 1'h0;
    2857: T462 = 1'h0;
    2858: T462 = 1'h0;
    2859: T462 = 1'h0;
    2860: T462 = 1'h0;
    2861: T462 = 1'h0;
    2862: T462 = 1'h0;
    2863: T462 = 1'h0;
    2864: T462 = 1'h0;
    2865: T462 = 1'h0;
    2866: T462 = 1'h0;
    2867: T462 = 1'h0;
    2868: T462 = 1'h0;
    2869: T462 = 1'h0;
    2870: T462 = 1'h0;
    2871: T462 = 1'h0;
    2872: T462 = 1'h0;
    2873: T462 = 1'h0;
    2874: T462 = 1'h0;
    2875: T462 = 1'h0;
    2876: T462 = 1'h0;
    2877: T462 = 1'h0;
    2878: T462 = 1'h0;
    2879: T462 = 1'h0;
    2880: T462 = 1'h0;
    2881: T462 = 1'h0;
    2882: T462 = 1'h0;
    2883: T462 = 1'h0;
    2884: T462 = 1'h0;
    2885: T462 = 1'h0;
    2886: T462 = 1'h0;
    2887: T462 = 1'h0;
    2888: T462 = 1'h0;
    2889: T462 = 1'h0;
    2890: T462 = 1'h0;
    2891: T462 = 1'h0;
    2892: T462 = 1'h0;
    2893: T462 = 1'h0;
    2894: T462 = 1'h0;
    2895: T462 = 1'h0;
    2896: T462 = 1'h0;
    2897: T462 = 1'h0;
    2898: T462 = 1'h0;
    2899: T462 = 1'h0;
    2900: T462 = 1'h0;
    2901: T462 = 1'h0;
    2902: T462 = 1'h0;
    2903: T462 = 1'h0;
    2904: T462 = 1'h0;
    2905: T462 = 1'h0;
    2906: T462 = 1'h0;
    2907: T462 = 1'h0;
    2908: T462 = 1'h0;
    2909: T462 = 1'h0;
    2910: T462 = 1'h0;
    2911: T462 = 1'h0;
    2912: T462 = 1'h0;
    2913: T462 = 1'h0;
    2914: T462 = 1'h0;
    2915: T462 = 1'h0;
    2916: T462 = 1'h0;
    2917: T462 = 1'h0;
    2918: T462 = 1'h0;
    2919: T462 = 1'h0;
    2920: T462 = 1'h0;
    2921: T462 = 1'h0;
    2922: T462 = 1'h0;
    2923: T462 = 1'h0;
    2924: T462 = 1'h0;
    2925: T462 = 1'h0;
    2926: T462 = 1'h0;
    2927: T462 = 1'h0;
    2928: T462 = 1'h0;
    2929: T462 = 1'h0;
    2930: T462 = 1'h0;
    2931: T462 = 1'h0;
    2932: T462 = 1'h0;
    2933: T462 = 1'h0;
    2934: T462 = 1'h0;
    2935: T462 = 1'h0;
    2936: T462 = 1'h0;
    2937: T462 = 1'h0;
    2938: T462 = 1'h0;
    2939: T462 = 1'h0;
    2940: T462 = 1'h0;
    2941: T462 = 1'h0;
    2942: T462 = 1'h0;
    2943: T462 = 1'h0;
    2944: T462 = 1'h0;
    2945: T462 = 1'h0;
    2946: T462 = 1'h0;
    2947: T462 = 1'h0;
    2948: T462 = 1'h0;
    2949: T462 = 1'h0;
    2950: T462 = 1'h0;
    2951: T462 = 1'h0;
    2952: T462 = 1'h0;
    2953: T462 = 1'h0;
    2954: T462 = 1'h0;
    2955: T462 = 1'h0;
    2956: T462 = 1'h0;
    2957: T462 = 1'h0;
    2958: T462 = 1'h0;
    2959: T462 = 1'h0;
    2960: T462 = 1'h0;
    2961: T462 = 1'h0;
    2962: T462 = 1'h0;
    2963: T462 = 1'h0;
    2964: T462 = 1'h0;
    2965: T462 = 1'h0;
    2966: T462 = 1'h0;
    2967: T462 = 1'h0;
    2968: T462 = 1'h0;
    2969: T462 = 1'h0;
    2970: T462 = 1'h0;
    2971: T462 = 1'h0;
    2972: T462 = 1'h0;
    2973: T462 = 1'h0;
    2974: T462 = 1'h0;
    2975: T462 = 1'h0;
    2976: T462 = 1'h0;
    2977: T462 = 1'h0;
    2978: T462 = 1'h0;
    2979: T462 = 1'h0;
    2980: T462 = 1'h0;
    2981: T462 = 1'h0;
    2982: T462 = 1'h0;
    2983: T462 = 1'h0;
    2984: T462 = 1'h0;
    2985: T462 = 1'h0;
    2986: T462 = 1'h0;
    2987: T462 = 1'h0;
    2988: T462 = 1'h0;
    2989: T462 = 1'h0;
    2990: T462 = 1'h0;
    2991: T462 = 1'h0;
    2992: T462 = 1'h0;
    2993: T462 = 1'h0;
    2994: T462 = 1'h0;
    2995: T462 = 1'h0;
    2996: T462 = 1'h0;
    2997: T462 = 1'h0;
    2998: T462 = 1'h0;
    2999: T462 = 1'h0;
    3000: T462 = 1'h0;
    3001: T462 = 1'h0;
    3002: T462 = 1'h0;
    3003: T462 = 1'h0;
    3004: T462 = 1'h0;
    3005: T462 = 1'h0;
    3006: T462 = 1'h0;
    3007: T462 = 1'h0;
    3008: T462 = 1'h0;
    3009: T462 = 1'h0;
    3010: T462 = 1'h0;
    3011: T462 = 1'h0;
    3012: T462 = 1'h0;
    3013: T462 = 1'h0;
    3014: T462 = 1'h0;
    3015: T462 = 1'h0;
    3016: T462 = 1'h0;
    3017: T462 = 1'h0;
    3018: T462 = 1'h0;
    3019: T462 = 1'h0;
    3020: T462 = 1'h0;
    3021: T462 = 1'h0;
    3022: T462 = 1'h0;
    3023: T462 = 1'h0;
    3024: T462 = 1'h0;
    3025: T462 = 1'h0;
    3026: T462 = 1'h0;
    3027: T462 = 1'h0;
    3028: T462 = 1'h0;
    3029: T462 = 1'h0;
    3030: T462 = 1'h0;
    3031: T462 = 1'h0;
    3032: T462 = 1'h0;
    3033: T462 = 1'h0;
    3034: T462 = 1'h0;
    3035: T462 = 1'h0;
    3036: T462 = 1'h0;
    3037: T462 = 1'h0;
    3038: T462 = 1'h0;
    3039: T462 = 1'h0;
    3040: T462 = 1'h0;
    3041: T462 = 1'h0;
    3042: T462 = 1'h0;
    3043: T462 = 1'h0;
    3044: T462 = 1'h0;
    3045: T462 = 1'h0;
    3046: T462 = 1'h0;
    3047: T462 = 1'h0;
    3048: T462 = 1'h0;
    3049: T462 = 1'h0;
    3050: T462 = 1'h0;
    3051: T462 = 1'h0;
    3052: T462 = 1'h0;
    3053: T462 = 1'h0;
    3054: T462 = 1'h0;
    3055: T462 = 1'h0;
    3056: T462 = 1'h0;
    3057: T462 = 1'h0;
    3058: T462 = 1'h0;
    3059: T462 = 1'h0;
    3060: T462 = 1'h0;
    3061: T462 = 1'h0;
    3062: T462 = 1'h0;
    3063: T462 = 1'h0;
    3064: T462 = 1'h0;
    3065: T462 = 1'h0;
    3066: T462 = 1'h0;
    3067: T462 = 1'h0;
    3068: T462 = 1'h0;
    3069: T462 = 1'h0;
    3070: T462 = 1'h0;
    3071: T462 = 1'h0;
    3072: T462 = 1'h1;
    3073: T462 = 1'h1;
    3074: T462 = 1'h1;
    3075: T462 = 1'h0;
    3076: T462 = 1'h0;
    3077: T462 = 1'h0;
    3078: T462 = 1'h0;
    3079: T462 = 1'h0;
    3080: T462 = 1'h0;
    3081: T462 = 1'h0;
    3082: T462 = 1'h0;
    3083: T462 = 1'h0;
    3084: T462 = 1'h0;
    3085: T462 = 1'h0;
    3086: T462 = 1'h0;
    3087: T462 = 1'h0;
    3088: T462 = 1'h0;
    3089: T462 = 1'h0;
    3090: T462 = 1'h0;
    3091: T462 = 1'h0;
    3092: T462 = 1'h0;
    3093: T462 = 1'h0;
    3094: T462 = 1'h0;
    3095: T462 = 1'h0;
    3096: T462 = 1'h0;
    3097: T462 = 1'h0;
    3098: T462 = 1'h0;
    3099: T462 = 1'h0;
    3100: T462 = 1'h0;
    3101: T462 = 1'h0;
    3102: T462 = 1'h0;
    3103: T462 = 1'h0;
    3104: T462 = 1'h0;
    3105: T462 = 1'h0;
    3106: T462 = 1'h0;
    3107: T462 = 1'h0;
    3108: T462 = 1'h0;
    3109: T462 = 1'h0;
    3110: T462 = 1'h0;
    3111: T462 = 1'h0;
    3112: T462 = 1'h0;
    3113: T462 = 1'h0;
    3114: T462 = 1'h0;
    3115: T462 = 1'h0;
    3116: T462 = 1'h0;
    3117: T462 = 1'h0;
    3118: T462 = 1'h0;
    3119: T462 = 1'h0;
    3120: T462 = 1'h0;
    3121: T462 = 1'h0;
    3122: T462 = 1'h0;
    3123: T462 = 1'h0;
    3124: T462 = 1'h0;
    3125: T462 = 1'h0;
    3126: T462 = 1'h0;
    3127: T462 = 1'h0;
    3128: T462 = 1'h0;
    3129: T462 = 1'h0;
    3130: T462 = 1'h0;
    3131: T462 = 1'h0;
    3132: T462 = 1'h0;
    3133: T462 = 1'h0;
    3134: T462 = 1'h0;
    3135: T462 = 1'h0;
    3136: T462 = 1'h0;
    3137: T462 = 1'h0;
    3138: T462 = 1'h0;
    3139: T462 = 1'h0;
    3140: T462 = 1'h0;
    3141: T462 = 1'h0;
    3142: T462 = 1'h0;
    3143: T462 = 1'h0;
    3144: T462 = 1'h0;
    3145: T462 = 1'h0;
    3146: T462 = 1'h0;
    3147: T462 = 1'h0;
    3148: T462 = 1'h0;
    3149: T462 = 1'h0;
    3150: T462 = 1'h0;
    3151: T462 = 1'h0;
    3152: T462 = 1'h0;
    3153: T462 = 1'h0;
    3154: T462 = 1'h0;
    3155: T462 = 1'h0;
    3156: T462 = 1'h0;
    3157: T462 = 1'h0;
    3158: T462 = 1'h0;
    3159: T462 = 1'h0;
    3160: T462 = 1'h0;
    3161: T462 = 1'h0;
    3162: T462 = 1'h0;
    3163: T462 = 1'h0;
    3164: T462 = 1'h0;
    3165: T462 = 1'h0;
    3166: T462 = 1'h0;
    3167: T462 = 1'h0;
    3168: T462 = 1'h0;
    3169: T462 = 1'h0;
    3170: T462 = 1'h0;
    3171: T462 = 1'h0;
    3172: T462 = 1'h0;
    3173: T462 = 1'h0;
    3174: T462 = 1'h0;
    3175: T462 = 1'h0;
    3176: T462 = 1'h0;
    3177: T462 = 1'h0;
    3178: T462 = 1'h0;
    3179: T462 = 1'h0;
    3180: T462 = 1'h0;
    3181: T462 = 1'h0;
    3182: T462 = 1'h0;
    3183: T462 = 1'h0;
    3184: T462 = 1'h0;
    3185: T462 = 1'h0;
    3186: T462 = 1'h0;
    3187: T462 = 1'h0;
    3188: T462 = 1'h0;
    3189: T462 = 1'h0;
    3190: T462 = 1'h0;
    3191: T462 = 1'h0;
    3192: T462 = 1'h0;
    3193: T462 = 1'h0;
    3194: T462 = 1'h0;
    3195: T462 = 1'h0;
    3196: T462 = 1'h0;
    3197: T462 = 1'h0;
    3198: T462 = 1'h0;
    3199: T462 = 1'h0;
    3200: T462 = 1'h0;
    3201: T462 = 1'h0;
    3202: T462 = 1'h0;
    3203: T462 = 1'h0;
    3204: T462 = 1'h0;
    3205: T462 = 1'h0;
    3206: T462 = 1'h0;
    3207: T462 = 1'h0;
    3208: T462 = 1'h0;
    3209: T462 = 1'h0;
    3210: T462 = 1'h0;
    3211: T462 = 1'h0;
    3212: T462 = 1'h0;
    3213: T462 = 1'h0;
    3214: T462 = 1'h0;
    3215: T462 = 1'h0;
    3216: T462 = 1'h0;
    3217: T462 = 1'h0;
    3218: T462 = 1'h0;
    3219: T462 = 1'h0;
    3220: T462 = 1'h0;
    3221: T462 = 1'h0;
    3222: T462 = 1'h0;
    3223: T462 = 1'h0;
    3224: T462 = 1'h0;
    3225: T462 = 1'h0;
    3226: T462 = 1'h0;
    3227: T462 = 1'h0;
    3228: T462 = 1'h0;
    3229: T462 = 1'h0;
    3230: T462 = 1'h0;
    3231: T462 = 1'h0;
    3232: T462 = 1'h0;
    3233: T462 = 1'h0;
    3234: T462 = 1'h0;
    3235: T462 = 1'h0;
    3236: T462 = 1'h0;
    3237: T462 = 1'h0;
    3238: T462 = 1'h0;
    3239: T462 = 1'h0;
    3240: T462 = 1'h0;
    3241: T462 = 1'h0;
    3242: T462 = 1'h0;
    3243: T462 = 1'h0;
    3244: T462 = 1'h0;
    3245: T462 = 1'h0;
    3246: T462 = 1'h0;
    3247: T462 = 1'h0;
    3248: T462 = 1'h0;
    3249: T462 = 1'h0;
    3250: T462 = 1'h0;
    3251: T462 = 1'h0;
    3252: T462 = 1'h0;
    3253: T462 = 1'h0;
    3254: T462 = 1'h0;
    3255: T462 = 1'h0;
    3256: T462 = 1'h0;
    3257: T462 = 1'h0;
    3258: T462 = 1'h0;
    3259: T462 = 1'h0;
    3260: T462 = 1'h0;
    3261: T462 = 1'h0;
    3262: T462 = 1'h0;
    3263: T462 = 1'h0;
    3264: T462 = 1'h1;
    3265: T462 = 1'h1;
    3266: T462 = 1'h1;
    3267: T462 = 1'h1;
    3268: T462 = 1'h1;
    3269: T462 = 1'h1;
    3270: T462 = 1'h1;
    3271: T462 = 1'h1;
    3272: T462 = 1'h1;
    3273: T462 = 1'h1;
    3274: T462 = 1'h1;
    3275: T462 = 1'h1;
    3276: T462 = 1'h1;
    3277: T462 = 1'h1;
    3278: T462 = 1'h1;
    3279: T462 = 1'h1;
    3280: T462 = 1'h0;
    3281: T462 = 1'h0;
    3282: T462 = 1'h0;
    3283: T462 = 1'h0;
    3284: T462 = 1'h0;
    3285: T462 = 1'h0;
    3286: T462 = 1'h0;
    3287: T462 = 1'h0;
    3288: T462 = 1'h0;
    3289: T462 = 1'h0;
    3290: T462 = 1'h0;
    3291: T462 = 1'h0;
    3292: T462 = 1'h0;
    3293: T462 = 1'h0;
    3294: T462 = 1'h0;
    3295: T462 = 1'h0;
    3296: T462 = 1'h0;
    3297: T462 = 1'h0;
    3298: T462 = 1'h0;
    3299: T462 = 1'h0;
    3300: T462 = 1'h0;
    3301: T462 = 1'h0;
    3302: T462 = 1'h0;
    3303: T462 = 1'h0;
    3304: T462 = 1'h0;
    3305: T462 = 1'h0;
    3306: T462 = 1'h0;
    3307: T462 = 1'h0;
    3308: T462 = 1'h0;
    3309: T462 = 1'h0;
    3310: T462 = 1'h0;
    3311: T462 = 1'h0;
    3312: T462 = 1'h0;
    3313: T462 = 1'h0;
    3314: T462 = 1'h0;
    3315: T462 = 1'h0;
    3316: T462 = 1'h0;
    3317: T462 = 1'h0;
    3318: T462 = 1'h0;
    3319: T462 = 1'h0;
    3320: T462 = 1'h0;
    3321: T462 = 1'h0;
    3322: T462 = 1'h0;
    3323: T462 = 1'h0;
    3324: T462 = 1'h0;
    3325: T462 = 1'h0;
    3326: T462 = 1'h0;
    3327: T462 = 1'h0;
    3328: T462 = 1'h0;
    3329: T462 = 1'h0;
    3330: T462 = 1'h0;
    3331: T462 = 1'h0;
    3332: T462 = 1'h0;
    3333: T462 = 1'h0;
    3334: T462 = 1'h0;
    3335: T462 = 1'h0;
    3336: T462 = 1'h0;
    3337: T462 = 1'h0;
    3338: T462 = 1'h0;
    3339: T462 = 1'h0;
    3340: T462 = 1'h0;
    3341: T462 = 1'h0;
    3342: T462 = 1'h0;
    3343: T462 = 1'h0;
    3344: T462 = 1'h0;
    3345: T462 = 1'h0;
    3346: T462 = 1'h0;
    3347: T462 = 1'h0;
    3348: T462 = 1'h0;
    3349: T462 = 1'h0;
    3350: T462 = 1'h0;
    3351: T462 = 1'h0;
    3352: T462 = 1'h0;
    3353: T462 = 1'h0;
    3354: T462 = 1'h0;
    3355: T462 = 1'h0;
    3356: T462 = 1'h0;
    3357: T462 = 1'h0;
    3358: T462 = 1'h0;
    3359: T462 = 1'h0;
    3360: T462 = 1'h0;
    3361: T462 = 1'h0;
    3362: T462 = 1'h0;
    3363: T462 = 1'h0;
    3364: T462 = 1'h0;
    3365: T462 = 1'h0;
    3366: T462 = 1'h0;
    3367: T462 = 1'h0;
    3368: T462 = 1'h0;
    3369: T462 = 1'h0;
    3370: T462 = 1'h0;
    3371: T462 = 1'h0;
    3372: T462 = 1'h0;
    3373: T462 = 1'h0;
    3374: T462 = 1'h0;
    3375: T462 = 1'h0;
    3376: T462 = 1'h0;
    3377: T462 = 1'h0;
    3378: T462 = 1'h0;
    3379: T462 = 1'h0;
    3380: T462 = 1'h0;
    3381: T462 = 1'h0;
    3382: T462 = 1'h0;
    3383: T462 = 1'h0;
    3384: T462 = 1'h0;
    3385: T462 = 1'h0;
    3386: T462 = 1'h0;
    3387: T462 = 1'h0;
    3388: T462 = 1'h0;
    3389: T462 = 1'h0;
    3390: T462 = 1'h0;
    3391: T462 = 1'h0;
    3392: T462 = 1'h0;
    3393: T462 = 1'h0;
    3394: T462 = 1'h0;
    3395: T462 = 1'h0;
    3396: T462 = 1'h0;
    3397: T462 = 1'h0;
    3398: T462 = 1'h0;
    3399: T462 = 1'h0;
    3400: T462 = 1'h0;
    3401: T462 = 1'h0;
    3402: T462 = 1'h0;
    3403: T462 = 1'h0;
    3404: T462 = 1'h0;
    3405: T462 = 1'h0;
    3406: T462 = 1'h0;
    3407: T462 = 1'h0;
    3408: T462 = 1'h0;
    3409: T462 = 1'h0;
    3410: T462 = 1'h0;
    3411: T462 = 1'h0;
    3412: T462 = 1'h0;
    3413: T462 = 1'h0;
    3414: T462 = 1'h0;
    3415: T462 = 1'h0;
    3416: T462 = 1'h0;
    3417: T462 = 1'h0;
    3418: T462 = 1'h0;
    3419: T462 = 1'h0;
    3420: T462 = 1'h0;
    3421: T462 = 1'h0;
    3422: T462 = 1'h0;
    3423: T462 = 1'h0;
    3424: T462 = 1'h0;
    3425: T462 = 1'h0;
    3426: T462 = 1'h0;
    3427: T462 = 1'h0;
    3428: T462 = 1'h0;
    3429: T462 = 1'h0;
    3430: T462 = 1'h0;
    3431: T462 = 1'h0;
    3432: T462 = 1'h0;
    3433: T462 = 1'h0;
    3434: T462 = 1'h0;
    3435: T462 = 1'h0;
    3436: T462 = 1'h0;
    3437: T462 = 1'h0;
    3438: T462 = 1'h0;
    3439: T462 = 1'h0;
    3440: T462 = 1'h0;
    3441: T462 = 1'h0;
    3442: T462 = 1'h0;
    3443: T462 = 1'h0;
    3444: T462 = 1'h0;
    3445: T462 = 1'h0;
    3446: T462 = 1'h0;
    3447: T462 = 1'h0;
    3448: T462 = 1'h0;
    3449: T462 = 1'h0;
    3450: T462 = 1'h0;
    3451: T462 = 1'h0;
    3452: T462 = 1'h0;
    3453: T462 = 1'h0;
    3454: T462 = 1'h0;
    3455: T462 = 1'h0;
    3456: T462 = 1'h0;
    3457: T462 = 1'h0;
    3458: T462 = 1'h0;
    3459: T462 = 1'h0;
    3460: T462 = 1'h0;
    3461: T462 = 1'h0;
    3462: T462 = 1'h0;
    3463: T462 = 1'h0;
    3464: T462 = 1'h0;
    3465: T462 = 1'h0;
    3466: T462 = 1'h0;
    3467: T462 = 1'h0;
    3468: T462 = 1'h0;
    3469: T462 = 1'h0;
    3470: T462 = 1'h0;
    3471: T462 = 1'h0;
    3472: T462 = 1'h0;
    3473: T462 = 1'h0;
    3474: T462 = 1'h0;
    3475: T462 = 1'h0;
    3476: T462 = 1'h0;
    3477: T462 = 1'h0;
    3478: T462 = 1'h0;
    3479: T462 = 1'h0;
    3480: T462 = 1'h0;
    3481: T462 = 1'h0;
    3482: T462 = 1'h0;
    3483: T462 = 1'h0;
    3484: T462 = 1'h0;
    3485: T462 = 1'h0;
    3486: T462 = 1'h0;
    3487: T462 = 1'h0;
    3488: T462 = 1'h0;
    3489: T462 = 1'h0;
    3490: T462 = 1'h0;
    3491: T462 = 1'h0;
    3492: T462 = 1'h0;
    3493: T462 = 1'h0;
    3494: T462 = 1'h0;
    3495: T462 = 1'h0;
    3496: T462 = 1'h0;
    3497: T462 = 1'h0;
    3498: T462 = 1'h0;
    3499: T462 = 1'h0;
    3500: T462 = 1'h0;
    3501: T462 = 1'h0;
    3502: T462 = 1'h0;
    3503: T462 = 1'h0;
    3504: T462 = 1'h0;
    3505: T462 = 1'h0;
    3506: T462 = 1'h0;
    3507: T462 = 1'h0;
    3508: T462 = 1'h0;
    3509: T462 = 1'h0;
    3510: T462 = 1'h0;
    3511: T462 = 1'h0;
    3512: T462 = 1'h0;
    3513: T462 = 1'h0;
    3514: T462 = 1'h0;
    3515: T462 = 1'h0;
    3516: T462 = 1'h0;
    3517: T462 = 1'h0;
    3518: T462 = 1'h0;
    3519: T462 = 1'h0;
    3520: T462 = 1'h0;
    3521: T462 = 1'h0;
    3522: T462 = 1'h0;
    3523: T462 = 1'h0;
    3524: T462 = 1'h0;
    3525: T462 = 1'h0;
    3526: T462 = 1'h0;
    3527: T462 = 1'h0;
    3528: T462 = 1'h0;
    3529: T462 = 1'h0;
    3530: T462 = 1'h0;
    3531: T462 = 1'h0;
    3532: T462 = 1'h0;
    3533: T462 = 1'h0;
    3534: T462 = 1'h0;
    3535: T462 = 1'h0;
    3536: T462 = 1'h0;
    3537: T462 = 1'h0;
    3538: T462 = 1'h0;
    3539: T462 = 1'h0;
    3540: T462 = 1'h0;
    3541: T462 = 1'h0;
    3542: T462 = 1'h0;
    3543: T462 = 1'h0;
    3544: T462 = 1'h0;
    3545: T462 = 1'h0;
    3546: T462 = 1'h0;
    3547: T462 = 1'h0;
    3548: T462 = 1'h0;
    3549: T462 = 1'h0;
    3550: T462 = 1'h0;
    3551: T462 = 1'h0;
    3552: T462 = 1'h0;
    3553: T462 = 1'h0;
    3554: T462 = 1'h0;
    3555: T462 = 1'h0;
    3556: T462 = 1'h0;
    3557: T462 = 1'h0;
    3558: T462 = 1'h0;
    3559: T462 = 1'h0;
    3560: T462 = 1'h0;
    3561: T462 = 1'h0;
    3562: T462 = 1'h0;
    3563: T462 = 1'h0;
    3564: T462 = 1'h0;
    3565: T462 = 1'h0;
    3566: T462 = 1'h0;
    3567: T462 = 1'h0;
    3568: T462 = 1'h0;
    3569: T462 = 1'h0;
    3570: T462 = 1'h0;
    3571: T462 = 1'h0;
    3572: T462 = 1'h0;
    3573: T462 = 1'h0;
    3574: T462 = 1'h0;
    3575: T462 = 1'h0;
    3576: T462 = 1'h0;
    3577: T462 = 1'h0;
    3578: T462 = 1'h0;
    3579: T462 = 1'h0;
    3580: T462 = 1'h0;
    3581: T462 = 1'h0;
    3582: T462 = 1'h0;
    3583: T462 = 1'h0;
    3584: T462 = 1'h0;
    3585: T462 = 1'h0;
    3586: T462 = 1'h0;
    3587: T462 = 1'h0;
    3588: T462 = 1'h0;
    3589: T462 = 1'h0;
    3590: T462 = 1'h0;
    3591: T462 = 1'h0;
    3592: T462 = 1'h0;
    3593: T462 = 1'h0;
    3594: T462 = 1'h0;
    3595: T462 = 1'h0;
    3596: T462 = 1'h0;
    3597: T462 = 1'h0;
    3598: T462 = 1'h0;
    3599: T462 = 1'h0;
    3600: T462 = 1'h0;
    3601: T462 = 1'h0;
    3602: T462 = 1'h0;
    3603: T462 = 1'h0;
    3604: T462 = 1'h0;
    3605: T462 = 1'h0;
    3606: T462 = 1'h0;
    3607: T462 = 1'h0;
    3608: T462 = 1'h0;
    3609: T462 = 1'h0;
    3610: T462 = 1'h0;
    3611: T462 = 1'h0;
    3612: T462 = 1'h0;
    3613: T462 = 1'h0;
    3614: T462 = 1'h0;
    3615: T462 = 1'h0;
    3616: T462 = 1'h0;
    3617: T462 = 1'h0;
    3618: T462 = 1'h0;
    3619: T462 = 1'h0;
    3620: T462 = 1'h0;
    3621: T462 = 1'h0;
    3622: T462 = 1'h0;
    3623: T462 = 1'h0;
    3624: T462 = 1'h0;
    3625: T462 = 1'h0;
    3626: T462 = 1'h0;
    3627: T462 = 1'h0;
    3628: T462 = 1'h0;
    3629: T462 = 1'h0;
    3630: T462 = 1'h0;
    3631: T462 = 1'h0;
    3632: T462 = 1'h0;
    3633: T462 = 1'h0;
    3634: T462 = 1'h0;
    3635: T462 = 1'h0;
    3636: T462 = 1'h0;
    3637: T462 = 1'h0;
    3638: T462 = 1'h0;
    3639: T462 = 1'h0;
    3640: T462 = 1'h0;
    3641: T462 = 1'h0;
    3642: T462 = 1'h0;
    3643: T462 = 1'h0;
    3644: T462 = 1'h0;
    3645: T462 = 1'h0;
    3646: T462 = 1'h0;
    3647: T462 = 1'h0;
    3648: T462 = 1'h0;
    3649: T462 = 1'h0;
    3650: T462 = 1'h0;
    3651: T462 = 1'h0;
    3652: T462 = 1'h0;
    3653: T462 = 1'h0;
    3654: T462 = 1'h0;
    3655: T462 = 1'h0;
    3656: T462 = 1'h0;
    3657: T462 = 1'h0;
    3658: T462 = 1'h0;
    3659: T462 = 1'h0;
    3660: T462 = 1'h0;
    3661: T462 = 1'h0;
    3662: T462 = 1'h0;
    3663: T462 = 1'h0;
    3664: T462 = 1'h0;
    3665: T462 = 1'h0;
    3666: T462 = 1'h0;
    3667: T462 = 1'h0;
    3668: T462 = 1'h0;
    3669: T462 = 1'h0;
    3670: T462 = 1'h0;
    3671: T462 = 1'h0;
    3672: T462 = 1'h0;
    3673: T462 = 1'h0;
    3674: T462 = 1'h0;
    3675: T462 = 1'h0;
    3676: T462 = 1'h0;
    3677: T462 = 1'h0;
    3678: T462 = 1'h0;
    3679: T462 = 1'h0;
    3680: T462 = 1'h0;
    3681: T462 = 1'h0;
    3682: T462 = 1'h0;
    3683: T462 = 1'h0;
    3684: T462 = 1'h0;
    3685: T462 = 1'h0;
    3686: T462 = 1'h0;
    3687: T462 = 1'h0;
    3688: T462 = 1'h0;
    3689: T462 = 1'h0;
    3690: T462 = 1'h0;
    3691: T462 = 1'h0;
    3692: T462 = 1'h0;
    3693: T462 = 1'h0;
    3694: T462 = 1'h0;
    3695: T462 = 1'h0;
    3696: T462 = 1'h0;
    3697: T462 = 1'h0;
    3698: T462 = 1'h0;
    3699: T462 = 1'h0;
    3700: T462 = 1'h0;
    3701: T462 = 1'h0;
    3702: T462 = 1'h0;
    3703: T462 = 1'h0;
    3704: T462 = 1'h0;
    3705: T462 = 1'h0;
    3706: T462 = 1'h0;
    3707: T462 = 1'h0;
    3708: T462 = 1'h0;
    3709: T462 = 1'h0;
    3710: T462 = 1'h0;
    3711: T462 = 1'h0;
    3712: T462 = 1'h0;
    3713: T462 = 1'h0;
    3714: T462 = 1'h0;
    3715: T462 = 1'h0;
    3716: T462 = 1'h0;
    3717: T462 = 1'h0;
    3718: T462 = 1'h0;
    3719: T462 = 1'h0;
    3720: T462 = 1'h0;
    3721: T462 = 1'h0;
    3722: T462 = 1'h0;
    3723: T462 = 1'h0;
    3724: T462 = 1'h0;
    3725: T462 = 1'h0;
    3726: T462 = 1'h0;
    3727: T462 = 1'h0;
    3728: T462 = 1'h0;
    3729: T462 = 1'h0;
    3730: T462 = 1'h0;
    3731: T462 = 1'h0;
    3732: T462 = 1'h0;
    3733: T462 = 1'h0;
    3734: T462 = 1'h0;
    3735: T462 = 1'h0;
    3736: T462 = 1'h0;
    3737: T462 = 1'h0;
    3738: T462 = 1'h0;
    3739: T462 = 1'h0;
    3740: T462 = 1'h0;
    3741: T462 = 1'h0;
    3742: T462 = 1'h0;
    3743: T462 = 1'h0;
    3744: T462 = 1'h0;
    3745: T462 = 1'h0;
    3746: T462 = 1'h0;
    3747: T462 = 1'h0;
    3748: T462 = 1'h0;
    3749: T462 = 1'h0;
    3750: T462 = 1'h0;
    3751: T462 = 1'h0;
    3752: T462 = 1'h0;
    3753: T462 = 1'h0;
    3754: T462 = 1'h0;
    3755: T462 = 1'h0;
    3756: T462 = 1'h0;
    3757: T462 = 1'h0;
    3758: T462 = 1'h0;
    3759: T462 = 1'h0;
    3760: T462 = 1'h0;
    3761: T462 = 1'h0;
    3762: T462 = 1'h0;
    3763: T462 = 1'h0;
    3764: T462 = 1'h0;
    3765: T462 = 1'h0;
    3766: T462 = 1'h0;
    3767: T462 = 1'h0;
    3768: T462 = 1'h0;
    3769: T462 = 1'h0;
    3770: T462 = 1'h0;
    3771: T462 = 1'h0;
    3772: T462 = 1'h0;
    3773: T462 = 1'h0;
    3774: T462 = 1'h0;
    3775: T462 = 1'h0;
    3776: T462 = 1'h0;
    3777: T462 = 1'h0;
    3778: T462 = 1'h0;
    3779: T462 = 1'h0;
    3780: T462 = 1'h0;
    3781: T462 = 1'h0;
    3782: T462 = 1'h0;
    3783: T462 = 1'h0;
    3784: T462 = 1'h0;
    3785: T462 = 1'h0;
    3786: T462 = 1'h0;
    3787: T462 = 1'h0;
    3788: T462 = 1'h0;
    3789: T462 = 1'h0;
    3790: T462 = 1'h0;
    3791: T462 = 1'h0;
    3792: T462 = 1'h0;
    3793: T462 = 1'h0;
    3794: T462 = 1'h0;
    3795: T462 = 1'h0;
    3796: T462 = 1'h0;
    3797: T462 = 1'h0;
    3798: T462 = 1'h0;
    3799: T462 = 1'h0;
    3800: T462 = 1'h0;
    3801: T462 = 1'h0;
    3802: T462 = 1'h0;
    3803: T462 = 1'h0;
    3804: T462 = 1'h0;
    3805: T462 = 1'h0;
    3806: T462 = 1'h0;
    3807: T462 = 1'h0;
    3808: T462 = 1'h0;
    3809: T462 = 1'h0;
    3810: T462 = 1'h0;
    3811: T462 = 1'h0;
    3812: T462 = 1'h0;
    3813: T462 = 1'h0;
    3814: T462 = 1'h0;
    3815: T462 = 1'h0;
    3816: T462 = 1'h0;
    3817: T462 = 1'h0;
    3818: T462 = 1'h0;
    3819: T462 = 1'h0;
    3820: T462 = 1'h0;
    3821: T462 = 1'h0;
    3822: T462 = 1'h0;
    3823: T462 = 1'h0;
    3824: T462 = 1'h0;
    3825: T462 = 1'h0;
    3826: T462 = 1'h0;
    3827: T462 = 1'h0;
    3828: T462 = 1'h0;
    3829: T462 = 1'h0;
    3830: T462 = 1'h0;
    3831: T462 = 1'h0;
    3832: T462 = 1'h0;
    3833: T462 = 1'h0;
    3834: T462 = 1'h0;
    3835: T462 = 1'h0;
    3836: T462 = 1'h0;
    3837: T462 = 1'h0;
    3838: T462 = 1'h0;
    3839: T462 = 1'h0;
    3840: T462 = 1'h0;
    3841: T462 = 1'h0;
    3842: T462 = 1'h0;
    3843: T462 = 1'h0;
    3844: T462 = 1'h0;
    3845: T462 = 1'h0;
    3846: T462 = 1'h0;
    3847: T462 = 1'h0;
    3848: T462 = 1'h0;
    3849: T462 = 1'h0;
    3850: T462 = 1'h0;
    3851: T462 = 1'h0;
    3852: T462 = 1'h0;
    3853: T462 = 1'h0;
    3854: T462 = 1'h0;
    3855: T462 = 1'h0;
    3856: T462 = 1'h0;
    3857: T462 = 1'h0;
    3858: T462 = 1'h0;
    3859: T462 = 1'h0;
    3860: T462 = 1'h0;
    3861: T462 = 1'h0;
    3862: T462 = 1'h0;
    3863: T462 = 1'h0;
    3864: T462 = 1'h0;
    3865: T462 = 1'h0;
    3866: T462 = 1'h0;
    3867: T462 = 1'h0;
    3868: T462 = 1'h0;
    3869: T462 = 1'h0;
    3870: T462 = 1'h0;
    3871: T462 = 1'h0;
    3872: T462 = 1'h0;
    3873: T462 = 1'h0;
    3874: T462 = 1'h0;
    3875: T462 = 1'h0;
    3876: T462 = 1'h0;
    3877: T462 = 1'h0;
    3878: T462 = 1'h0;
    3879: T462 = 1'h0;
    3880: T462 = 1'h0;
    3881: T462 = 1'h0;
    3882: T462 = 1'h0;
    3883: T462 = 1'h0;
    3884: T462 = 1'h0;
    3885: T462 = 1'h0;
    3886: T462 = 1'h0;
    3887: T462 = 1'h0;
    3888: T462 = 1'h0;
    3889: T462 = 1'h0;
    3890: T462 = 1'h0;
    3891: T462 = 1'h0;
    3892: T462 = 1'h0;
    3893: T462 = 1'h0;
    3894: T462 = 1'h0;
    3895: T462 = 1'h0;
    3896: T462 = 1'h0;
    3897: T462 = 1'h0;
    3898: T462 = 1'h0;
    3899: T462 = 1'h0;
    3900: T462 = 1'h0;
    3901: T462 = 1'h0;
    3902: T462 = 1'h0;
    3903: T462 = 1'h0;
    3904: T462 = 1'h0;
    3905: T462 = 1'h0;
    3906: T462 = 1'h0;
    3907: T462 = 1'h0;
    3908: T462 = 1'h0;
    3909: T462 = 1'h0;
    3910: T462 = 1'h0;
    3911: T462 = 1'h0;
    3912: T462 = 1'h0;
    3913: T462 = 1'h0;
    3914: T462 = 1'h0;
    3915: T462 = 1'h0;
    3916: T462 = 1'h0;
    3917: T462 = 1'h0;
    3918: T462 = 1'h0;
    3919: T462 = 1'h0;
    3920: T462 = 1'h0;
    3921: T462 = 1'h0;
    3922: T462 = 1'h0;
    3923: T462 = 1'h0;
    3924: T462 = 1'h0;
    3925: T462 = 1'h0;
    3926: T462 = 1'h0;
    3927: T462 = 1'h0;
    3928: T462 = 1'h0;
    3929: T462 = 1'h0;
    3930: T462 = 1'h0;
    3931: T462 = 1'h0;
    3932: T462 = 1'h0;
    3933: T462 = 1'h0;
    3934: T462 = 1'h0;
    3935: T462 = 1'h0;
    3936: T462 = 1'h0;
    3937: T462 = 1'h0;
    3938: T462 = 1'h0;
    3939: T462 = 1'h0;
    3940: T462 = 1'h0;
    3941: T462 = 1'h0;
    3942: T462 = 1'h0;
    3943: T462 = 1'h0;
    3944: T462 = 1'h0;
    3945: T462 = 1'h0;
    3946: T462 = 1'h0;
    3947: T462 = 1'h0;
    3948: T462 = 1'h0;
    3949: T462 = 1'h0;
    3950: T462 = 1'h0;
    3951: T462 = 1'h0;
    3952: T462 = 1'h0;
    3953: T462 = 1'h0;
    3954: T462 = 1'h0;
    3955: T462 = 1'h0;
    3956: T462 = 1'h0;
    3957: T462 = 1'h0;
    3958: T462 = 1'h0;
    3959: T462 = 1'h0;
    3960: T462 = 1'h0;
    3961: T462 = 1'h0;
    3962: T462 = 1'h0;
    3963: T462 = 1'h0;
    3964: T462 = 1'h0;
    3965: T462 = 1'h0;
    3966: T462 = 1'h0;
    3967: T462 = 1'h0;
    3968: T462 = 1'h0;
    3969: T462 = 1'h0;
    3970: T462 = 1'h0;
    3971: T462 = 1'h0;
    3972: T462 = 1'h0;
    3973: T462 = 1'h0;
    3974: T462 = 1'h0;
    3975: T462 = 1'h0;
    3976: T462 = 1'h0;
    3977: T462 = 1'h0;
    3978: T462 = 1'h0;
    3979: T462 = 1'h0;
    3980: T462 = 1'h0;
    3981: T462 = 1'h0;
    3982: T462 = 1'h0;
    3983: T462 = 1'h0;
    3984: T462 = 1'h0;
    3985: T462 = 1'h0;
    3986: T462 = 1'h0;
    3987: T462 = 1'h0;
    3988: T462 = 1'h0;
    3989: T462 = 1'h0;
    3990: T462 = 1'h0;
    3991: T462 = 1'h0;
    3992: T462 = 1'h0;
    3993: T462 = 1'h0;
    3994: T462 = 1'h0;
    3995: T462 = 1'h0;
    3996: T462 = 1'h0;
    3997: T462 = 1'h0;
    3998: T462 = 1'h0;
    3999: T462 = 1'h0;
    4000: T462 = 1'h0;
    4001: T462 = 1'h0;
    4002: T462 = 1'h0;
    4003: T462 = 1'h0;
    4004: T462 = 1'h0;
    4005: T462 = 1'h0;
    4006: T462 = 1'h0;
    4007: T462 = 1'h0;
    4008: T462 = 1'h0;
    4009: T462 = 1'h0;
    4010: T462 = 1'h0;
    4011: T462 = 1'h0;
    4012: T462 = 1'h0;
    4013: T462 = 1'h0;
    4014: T462 = 1'h0;
    4015: T462 = 1'h0;
    4016: T462 = 1'h0;
    4017: T462 = 1'h0;
    4018: T462 = 1'h0;
    4019: T462 = 1'h0;
    4020: T462 = 1'h0;
    4021: T462 = 1'h0;
    4022: T462 = 1'h0;
    4023: T462 = 1'h0;
    4024: T462 = 1'h0;
    4025: T462 = 1'h0;
    4026: T462 = 1'h0;
    4027: T462 = 1'h0;
    4028: T462 = 1'h0;
    4029: T462 = 1'h0;
    4030: T462 = 1'h0;
    4031: T462 = 1'h0;
    4032: T462 = 1'h0;
    4033: T462 = 1'h0;
    4034: T462 = 1'h0;
    4035: T462 = 1'h0;
    4036: T462 = 1'h0;
    4037: T462 = 1'h0;
    4038: T462 = 1'h0;
    4039: T462 = 1'h0;
    4040: T462 = 1'h0;
    4041: T462 = 1'h0;
    4042: T462 = 1'h0;
    4043: T462 = 1'h0;
    4044: T462 = 1'h0;
    4045: T462 = 1'h0;
    4046: T462 = 1'h0;
    4047: T462 = 1'h0;
    4048: T462 = 1'h0;
    4049: T462 = 1'h0;
    4050: T462 = 1'h0;
    4051: T462 = 1'h0;
    4052: T462 = 1'h0;
    4053: T462 = 1'h0;
    4054: T462 = 1'h0;
    4055: T462 = 1'h0;
    4056: T462 = 1'h0;
    4057: T462 = 1'h0;
    4058: T462 = 1'h0;
    4059: T462 = 1'h0;
    4060: T462 = 1'h0;
    4061: T462 = 1'h0;
    4062: T462 = 1'h0;
    4063: T462 = 1'h0;
    4064: T462 = 1'h0;
    4065: T462 = 1'h0;
    4066: T462 = 1'h0;
    4067: T462 = 1'h0;
    4068: T462 = 1'h0;
    4069: T462 = 1'h0;
    4070: T462 = 1'h0;
    4071: T462 = 1'h0;
    4072: T462 = 1'h0;
    4073: T462 = 1'h0;
    4074: T462 = 1'h0;
    4075: T462 = 1'h0;
    4076: T462 = 1'h0;
    4077: T462 = 1'h0;
    4078: T462 = 1'h0;
    4079: T462 = 1'h0;
    4080: T462 = 1'h0;
    4081: T462 = 1'h0;
    4082: T462 = 1'h0;
    4083: T462 = 1'h0;
    4084: T462 = 1'h0;
    4085: T462 = 1'h0;
    4086: T462 = 1'h0;
    4087: T462 = 1'h0;
    4088: T462 = 1'h0;
    4089: T462 = 1'h0;
    4090: T462 = 1'h0;
    4091: T462 = 1'h0;
    4092: T462 = 1'h0;
    4093: T462 = 1'h0;
    4094: T462 = 1'h0;
    4095: T462 = 1'h0;
`ifndef SYNTHESIS
    default: T462 = {1{$random}};
`else
    default: T462 = 1'bx;
`endif
  endcase
  assign T464 = id_int_val ^ 1'h1;
  assign id_int_val = T467 | T465;
  assign T465 = T466 == 32'h33;
  assign T466 = io_dpath_inst & 32'hfc007077;
  assign T467 = T470 | T468;
  assign T468 = T469 == 32'h4063;
  assign T469 = io_dpath_inst & 32'h407f;
  assign T470 = T473 | T471;
  assign T471 = T472 == 32'h1063;
  assign T472 = io_dpath_inst & 32'h306f;
  assign T473 = T476 | T474;
  assign T474 = T475 == 32'h23;
  assign T475 = io_dpath_inst & 32'h603f;
  assign T476 = T479 | T477;
  assign T477 = T478 == 32'he0000053;
  assign T478 = io_dpath_inst & 32'hedf0707f;
  assign T479 = T482 | T480;
  assign T480 = T481 == 32'he0000053;
  assign T481 = io_dpath_inst & 32'hfdf0607f;
  assign T482 = T485 | T483;
  assign T483 = T484 == 32'hc0000053;
  assign T484 = io_dpath_inst & 32'hedc0007f;
  assign T485 = T488 | T486;
  assign T486 = T487 == 32'h42000053;
  assign T487 = io_dpath_inst & 32'h7ff0007f;
  assign T488 = T491 | T489;
  assign T489 = T490 == 32'h40100053;
  assign T490 = io_dpath_inst & 32'h7ff0007f;
  assign T491 = T494 | T492;
  assign T492 = T493 == 32'h20000053;
  assign T493 = io_dpath_inst & 32'h7c00507f;
  assign T494 = T497 | T495;
  assign T495 = T496 == 32'h20000053;
  assign T496 = io_dpath_inst & 32'h7c00607f;
  assign T497 = T500 | T498;
  assign T498 = T499 == 32'h20000053;
  assign T499 = io_dpath_inst & 32'hf400607f;
  assign T500 = T501 | T63;
  assign T501 = T502 | T66;
  assign T502 = T505 | T503;
  assign T503 = T504 == 32'h2004033;
  assign T504 = io_dpath_inst & 32'hfe004077;
  assign T505 = T508 | T506;
  assign T506 = T507 == 32'h5033;
  assign T507 = io_dpath_inst & 32'hbe007077;
  assign T508 = T511 | T509;
  assign T509 = T510 == 32'h501b;
  assign T510 = io_dpath_inst & 32'hbe00705f;
  assign T511 = T514 | T512;
  assign T512 = T513 == 32'h5013;
  assign T513 = io_dpath_inst & 32'hbc00707f;
  assign T514 = T517 | T515;
  assign T515 = T516 == 32'h2073;
  assign T516 = io_dpath_inst & 32'h207f;
  assign T517 = T518 | T69;
  assign T518 = T521 | T519;
  assign T519 = T520 == 32'h2013;
  assign T520 = io_dpath_inst & 32'h207f;
  assign T521 = T522 | T72;
  assign T522 = T525 | T523;
  assign T523 = T524 == 32'h101b;
  assign T524 = io_dpath_inst & 32'hfe00305f;
  assign T525 = T528 | T526;
  assign T526 = T527 == 32'h1013;
  assign T527 = io_dpath_inst & 32'hfc00305f;
  assign T528 = T531 | T529;
  assign T529 = T530 == 32'h73;
  assign T530 = io_dpath_inst & 32'h7fffffff;
  assign T531 = T534 | T532;
  assign T532 = T533 == 32'h6f;
  assign T533 = io_dpath_inst & 32'h7f;
  assign T534 = T537 | T535;
  assign T535 = T536 == 32'h63;
  assign T536 = io_dpath_inst & 32'h707b;
  assign T537 = T540 | T538;
  assign T538 = T539 == 32'h53;
  assign T539 = io_dpath_inst & 32'hec00007f;
  assign T540 = T543 | T541;
  assign T541 = T542 == 32'h53;
  assign T542 = io_dpath_inst & 32'hf400007f;
  assign T543 = T546 | T544;
  assign T544 = T545 == 32'h43;
  assign T545 = io_dpath_inst & 32'h4000073;
  assign T546 = T549 | T547;
  assign T547 = T548 == 32'h33;
  assign T548 = io_dpath_inst & 32'hbe007077;
  assign T549 = T552 | T550;
  assign T550 = T551 == 32'h33;
  assign T551 = io_dpath_inst & 32'hfc00007f;
  assign T552 = T555 | T553;
  assign T553 = T554 == 32'h17;
  assign T554 = io_dpath_inst & 32'h5f;
  assign T555 = T558 | T556;
  assign T556 = T557 == 32'h13;
  assign T557 = io_dpath_inst & 32'h7077;
  assign T558 = T561 | T559;
  assign T559 = T560 == 32'hf;
  assign T560 = io_dpath_inst & 32'h607f;
  assign T561 = T78 | T562;
  assign T562 = T563 == 32'h3;
  assign T563 = io_dpath_inst & 32'h106f;
  assign T564 = T565 | io_imem_resp_bits_xcpt_if;
  assign T565 = id_interrupt | io_imem_resp_bits_xcpt_ma;
  assign T566 = T567 & io_imem_resp_valid;
  assign T567 = id_interrupt & T568;
  assign T568 = take_pc ^ 1'h1;
  assign T569 = dcache_kill_mem | take_pc_wb;
  assign T570 = replay_wb | wb_reg_xcpt;
  assign mem_xcpt = T572 | T571;
  assign T571 = mem_reg_mem_val & io_dmem_xcpt_pf_st;
  assign T572 = T574 | T573;
  assign T573 = mem_reg_mem_val & io_dmem_xcpt_pf_ld;
  assign T574 = T576 | T575;
  assign T575 = mem_reg_mem_val & io_dmem_xcpt_ma_st;
  assign T576 = T578 | T577;
  assign T577 = mem_reg_mem_val & io_dmem_xcpt_ma_ld;
  assign T578 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T579 = T581 & T580;
  assign T580 = mem_reg_replay_next ^ 1'h1;
  assign T581 = T582 & ex_reg_xcpt_interrupt;
  assign T582 = take_pc ^ 1'h1;
  assign io_rocc_s = io_dpath_status_s;
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = wb_reg_rocc_val & T583;
  assign T583 = replay_wb_common ^ 1'h1;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T584;
  assign T584 = T585 & id_fp_val;
  assign T585 = ctrl_killd ^ 1'h1;
  assign io_dmem_req_bits_cmd = ex_reg_mem_cmd;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_typ = ex_reg_mem_type;
  assign io_dmem_req_bits_kill = T586;
  assign T586 = killm_common | mem_xcpt;
  assign io_dmem_req_valid = ex_reg_mem_val;
  assign io_imem_invalidate = wb_reg_flush_inst;
  assign T587 = ctrl_killm ? 1'h0 : mem_reg_flush_inst;
  assign T588 = ctrl_killx ? 1'h0 : ex_reg_flush_inst;
  assign T589 = ctrl_killd ? 1'h0 : id_fence_i;
  assign io_imem_btb_update_bits_mispredict = take_pc_mem;
  assign io_imem_btb_update_bits_isReturn = T590;
  assign T590 = mem_reg_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_btb_update_bits_isCall = T591;
  assign T591 = mem_reg_wen & T592;
  assign T592 = io_dpath_mem_waddr[1'h0:1'h0];
  assign io_imem_btb_update_bits_isJump = T593;
  assign T593 = mem_reg_jal | mem_reg_jalr;
  assign io_imem_btb_update_bits_taken = T594;
  assign T594 = T595 | io_imem_btb_update_bits_isJump;
  assign T595 = mem_reg_branch & io_dpath_mem_br_taken;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T596 = T599 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T597 = T598 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T598 = T320 & io_imem_btb_resp_valid;
  assign T599 = T352 & ex_reg_btb_hit;
  assign T600 = ctrl_killd ? 1'h0 : io_imem_btb_resp_valid;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T601 = T599 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T602 = T598 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T603 = T599 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T604 = T598 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T605 = T599 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T606 = T598 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T607 = T599 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T608 = T598 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T609 = T352 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T610;
  assign T610 = T612 & T611;
  assign T611 = take_pc_wb ^ 1'h1;
  assign T612 = mem_reg_branch | io_imem_btb_update_bits_isJump;
  assign io_imem_resp_ready = T613;
  assign T613 = T614 | ctrl_draind;
  assign T614 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_valid = take_pc;
  assign io_dpath_badvaddr_wen = wb_reg_xcpt;
  assign io_dpath_cause = wb_reg_cause;
  assign T615 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T578 ? mem_reg_cause : T796;
  assign T796 = {60'h0, T616};
  assign T616 = T577 ? 4'h8 : T617;
  assign T617 = T575 ? 4'h9 : T618;
  assign T618 = T573 ? 4'ha : 4'hb;
  assign T619 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T426 ? ex_reg_cause : 64'h2;
  assign T620 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = id_interrupt ? id_interrupt_cause : T797;
  assign T797 = {60'h0, T621};
  assign T621 = io_imem_resp_bits_xcpt_ma ? 4'h0 : T622;
  assign T622 = io_imem_resp_bits_xcpt_if ? 4'h1 : T623;
  assign T623 = T460 ? 4'h2 : T624;
  assign T624 = id_csr_privileged ? 4'h3 : T625;
  assign T625 = T436 ? 4'h3 : T626;
  assign T626 = T430 ? 4'h4 : T627;
  assign T627 = id_syscall ? 4'h6 : 4'hc;
  assign id_interrupt_cause = T56 ? 64'h8000000000000000 : T628;
  assign T628 = T53 ? 64'h8000000000000001 : T629;
  assign T629 = T49 ? 64'h8000000000000002 : T630;
  assign T630 = T45 ? 64'h8000000000000003 : T631;
  assign T631 = T41 ? 64'h8000000000000004 : T632;
  assign T632 = T37 ? 64'h8000000000000005 : T633;
  assign T633 = T33 ? 64'h8000000000000006 : 64'h8000000000000007;
  assign io_dpath_exception = wb_reg_xcpt;
  assign io_dpath_retire = T634;
  assign T634 = wb_reg_valid & T635;
  assign T635 = replay_wb ^ 1'h1;
  assign T636 = ctrl_killm ? 1'h0 : mem_reg_valid;
  assign io_dpath_ll_ready = T637;
  assign T637 = wb_reg_wen ^ 1'h1;
  assign io_dpath_bypass_src_0 = T638;
  assign T638 = T647 ? 2'h0 : T639;
  assign T639 = T645 ? 2'h1 : T640;
  assign T640 = T641 ? 2'h2 : 2'h3;
  assign T641 = T643 & T642;
  assign T642 = io_dpath_mem_waddr == id_raddr1;
  assign T643 = mem_reg_wen & T644;
  assign T644 = mem_reg_mem_val ^ 1'h1;
  assign T645 = ex_reg_wen & T646;
  assign T646 = io_dpath_ex_waddr == id_raddr1;
  assign T647 = 5'h0 == id_raddr1;
  assign io_dpath_bypass_src_1 = T648;
  assign T648 = T655 ? 2'h0 : T649;
  assign T649 = T653 ? 2'h1 : T650;
  assign T650 = T651 ? 2'h2 : 2'h3;
  assign T651 = T643 & T652;
  assign T652 = io_dpath_mem_waddr == id_raddr2;
  assign T653 = ex_reg_wen & T654;
  assign T654 = io_dpath_ex_waddr == id_raddr2;
  assign T655 = 5'h0 == id_raddr2;
  assign io_dpath_bypass_0 = T656;
  assign T656 = T659 | T657;
  assign T657 = mem_reg_wen & T658;
  assign T658 = io_dpath_mem_waddr == id_raddr1;
  assign T659 = T660 | T641;
  assign T660 = T647 | T645;
  assign io_dpath_bypass_1 = T661;
  assign T661 = T664 | T662;
  assign T662 = mem_reg_wen & T663;
  assign T663 = io_dpath_mem_waddr == id_raddr2;
  assign T664 = T665 | T651;
  assign T665 = T655 | T653;
  assign io_dpath_mem_rocc_val = mem_reg_rocc_val;
  assign io_dpath_ex_rocc_val = ex_reg_rocc_val;
  assign io_dpath_ex_rs2_val = T666;
  assign T666 = T667 | ex_reg_rocc_val;
  assign T667 = ex_reg_mem_val & T668;
  assign T668 = T672 | T669;
  assign T669 = T671 | T670;
  assign T670 = ex_reg_mem_cmd == 5'h4;
  assign T671 = ex_reg_mem_cmd[2'h3:2'h3];
  assign T672 = T674 | T673;
  assign T673 = ex_reg_mem_cmd == 5'h7;
  assign T674 = ex_reg_mem_cmd == 5'h1;
  assign io_dpath_ex_mem_type = ex_reg_mem_type;
  assign io_dpath_wb_wen = T675;
  assign T675 = wb_reg_wen & T676;
  assign T676 = replay_wb ^ 1'h1;
  assign io_dpath_mem_wen = mem_reg_wen;
  assign io_dpath_mem_branch = mem_reg_branch;
  assign io_dpath_mem_jalr = mem_reg_jalr;
  assign io_dpath_ex_valid = ex_reg_valid;
  assign io_dpath_ex_wen = ex_reg_wen;
  assign io_dpath_mem_fp_val = mem_reg_fp_val;
  assign io_dpath_ex_fp_val = ex_reg_fp_val;
  assign io_dpath_wb_load = T677;
  assign T677 = wb_reg_mem_val & wb_reg_wen;
  assign io_dpath_mem_load = T678;
  assign T678 = mem_reg_mem_val & mem_reg_wen;
  assign io_dpath_sret = wb_reg_sret;
  assign io_dpath_csr = T798;
  assign T798 = {1'h0, wb_reg_csr};
  assign T679 = ctrl_killm ? 2'h0 : mem_reg_csr;
  assign io_dpath_div_mul_kill = T680;
  assign T680 = mem_reg_div_mul_val & killm_common;
  assign io_dpath_div_mul_val = ex_reg_div_mul_val;
  assign io_dpath_fn_alu = T681;
  assign T681 = id_fn_alu;
  assign id_fn_alu = {T717, T682};
  assign T682 = {T706, T683};
  assign T683 = {T692, T684};
  assign T684 = T687 | T685;
  assign T685 = T686 == 32'h7000;
  assign T686 = io_dpath_inst & 32'h7044;
  assign T687 = T690 | T688;
  assign T688 = T689 == 32'h1040;
  assign T689 = io_dpath_inst & 32'h1058;
  assign T690 = T691 == 32'h1010;
  assign T691 = io_dpath_inst & 32'h3054;
  assign T692 = T695 | T693;
  assign T693 = T694 == 32'h40001010;
  assign T694 = io_dpath_inst & 32'h40001054;
  assign T695 = T698 | T696;
  assign T696 = T697 == 32'h40000030;
  assign T697 = io_dpath_inst & 32'h40003034;
  assign T698 = T701 | T699;
  assign T699 = T700 == 32'h6010;
  assign T700 = io_dpath_inst & 32'h6054;
  assign T701 = T704 | T702;
  assign T702 = T703 == 32'h3010;
  assign T703 = io_dpath_inst & 32'h3054;
  assign T704 = T705 == 32'h2040;
  assign T705 = io_dpath_inst & 32'h2058;
  assign T706 = T709 | T707;
  assign T707 = T708 == 32'h4040;
  assign T708 = io_dpath_inst & 32'h4058;
  assign T709 = T712 | T710;
  assign T710 = T711 == 32'h4010;
  assign T711 = io_dpath_inst & 32'h5054;
  assign T712 = T715 | T713;
  assign T713 = T714 == 32'h4010;
  assign T714 = io_dpath_inst & 32'h40004054;
  assign T715 = T716 == 32'h2010;
  assign T716 = io_dpath_inst & 32'h2054;
  assign T717 = T720 | T718;
  assign T718 = T719 == 32'h40001010;
  assign T719 = io_dpath_inst & 32'h40003054;
  assign T720 = T721 | T696;
  assign T721 = T724 | T722;
  assign T722 = T723 == 32'h2010;
  assign T723 = io_dpath_inst & 32'h6054;
  assign T724 = T725 == 32'h40;
  assign T725 = io_dpath_inst & 32'h54;
  assign io_dpath_fn_dw = T726;
  assign T726 = id_fn_dw;
  assign id_fn_dw = T729 | T727;
  assign T727 = T728 == 32'h0;
  assign T728 = io_dpath_inst & 32'h8;
  assign T729 = T730 == 32'h0;
  assign T730 = io_dpath_inst & 32'h10;
  assign io_dpath_sel_imm = T731;
  assign T731 = id_sel_imm;
  assign id_sel_imm = {T741, T732};
  assign T732 = {T738, T733};
  assign T733 = T736 | T734;
  assign T734 = T735 == 32'h40;
  assign T735 = io_dpath_inst & 32'h44;
  assign T736 = T737 == 32'h8;
  assign T737 = io_dpath_inst & 32'h18;
  assign T738 = T736 | T739;
  assign T739 = T740 == 32'h14;
  assign T740 = io_dpath_inst & 32'h14;
  assign T741 = T744 | T742;
  assign T742 = T743 == 32'h10;
  assign T743 = io_dpath_inst & 32'h14;
  assign T744 = T747 | T745;
  assign T745 = T746 == 32'h4;
  assign T746 = io_dpath_inst & 32'h201c;
  assign T747 = T748 == 32'h0;
  assign T748 = io_dpath_inst & 32'h30;
  assign io_dpath_sel_alu1 = T749;
  assign T749 = id_sel_alu1;
  assign id_sel_alu1 = {T762, T750};
  assign T750 = T753 | T751;
  assign T751 = T752 == 32'h0;
  assign T752 = io_dpath_inst & 32'h18;
  assign T753 = T756 | T754;
  assign T754 = T755 == 32'h0;
  assign T755 = io_dpath_inst & 32'h24;
  assign T756 = T757 | T262;
  assign T757 = T760 | T758;
  assign T758 = T759 == 32'h0;
  assign T759 = io_dpath_inst & 32'h50;
  assign T760 = T761 == 32'h0;
  assign T761 = io_dpath_inst & 32'h4004;
  assign T762 = T765 | T763;
  assign T763 = T764 == 32'h48;
  assign T764 = io_dpath_inst & 32'h48;
  assign T765 = T766 == 32'h14;
  assign T766 = io_dpath_inst & 32'h34;
  assign io_dpath_sel_alu2 = T799;
  assign T799 = {1'h0, T767};
  assign T767 = id_sel_alu2;
  assign id_sel_alu2 = {T780, T768};
  assign T768 = T771 | T769;
  assign T769 = T770 == 32'h4050;
  assign T770 = io_dpath_inst & 32'h4050;
  assign T771 = T772 | T763;
  assign T772 = T775 | T773;
  assign T773 = T774 == 32'h4;
  assign T774 = io_dpath_inst & 32'hc;
  assign T775 = T778 | T776;
  assign T776 = T777 == 32'h0;
  assign T777 = io_dpath_inst & 32'h20;
  assign T778 = T779 == 32'h0;
  assign T779 = io_dpath_inst & 32'h58;
  assign T780 = T783 | T781;
  assign T781 = T782 == 32'h4000;
  assign T782 = io_dpath_inst & 32'h4008;
  assign T783 = T784 | T751;
  assign T784 = T785 | T262;
  assign T785 = T786 == 32'h0;
  assign T786 = io_dpath_inst & 32'h48;
  assign io_dpath_ren_0 = id_renx1;
  assign io_dpath_ren_1 = id_renx2;
  assign io_dpath_killd = T787;
  assign T787 = take_pc | T788;
  assign T788 = ctrl_stalld & T789;
  assign T789 = ctrl_draind ^ 1'h1;
  assign io_dpath_sel_pc = T800;
  assign T800 = {1'h0, T790};
  assign T790 = wb_reg_xcpt ? 2'h3 : T791;
  assign T791 = wb_reg_sret ? 2'h3 : T792;
  assign T792 = replay_wb ? 2'h2 : 2'h1;

  always @(posedge clk) begin
    wb_reg_xcpt <= T1;
    if(ctrl_killm) begin
      wb_reg_sret <= 1'h0;
    end else begin
      wb_reg_sret <= T5;
    end
    mem_reg_replay <= T7;
    if(ctrl_killx) begin
      mem_reg_replay_next <= 1'h0;
    end else begin
      mem_reg_replay_next <= ex_reg_replay_next;
    end
    if(ctrl_killd) begin
      ex_reg_replay_next <= 1'h0;
    end else begin
      ex_reg_replay_next <= T10;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T82;
    end
    if(ctrl_killd) begin
      ex_reg_mem_val <= 1'h0;
    end else begin
      ex_reg_mem_val <= T91;
    end
    if(reset) begin
      R105 <= 32'h0;
    end else if(T165) begin
      R105 <= T161;
    end else if(T160) begin
      R105 <= T156;
    end else if(T112) begin
      R105 <= T109;
    end
    if(ctrl_killm) begin
      wb_reg_rocc_val <= 1'h0;
    end else begin
      wb_reg_rocc_val <= mem_reg_rocc_val;
    end
    if(ctrl_killx) begin
      mem_reg_rocc_val <= 1'h0;
    end else begin
      mem_reg_rocc_val <= ex_reg_rocc_val;
    end
    if(ctrl_killd) begin
      ex_reg_rocc_val <= 1'h0;
    end else begin
      ex_reg_rocc_val <= T119;
    end
    wb_reg_replay <= T121;
    if(ctrl_killx) begin
      mem_reg_fp_val <= 1'h0;
    end else begin
      mem_reg_fp_val <= ex_reg_fp_val;
    end
    if(ctrl_killd) begin
      ex_reg_fp_val <= 1'h0;
    end else begin
      ex_reg_fp_val <= id_fp_val;
    end
    if(ctrl_killx) begin
      mem_reg_wen <= 1'h0;
    end else begin
      mem_reg_wen <= ex_reg_wen;
    end
    if(ctrl_killd) begin
      ex_reg_wen <= 1'h0;
    end else begin
      ex_reg_wen <= id_wen;
    end
    if(ctrl_killm) begin
      wb_reg_fp_wen <= 1'h0;
    end else begin
      wb_reg_fp_wen <= mem_reg_fp_wen;
    end
    if(ctrl_killx) begin
      mem_reg_fp_wen <= 1'h0;
    end else begin
      mem_reg_fp_wen <= ex_reg_fp_wen;
    end
    if(ctrl_killd) begin
      ex_reg_fp_wen <= 1'h0;
    end else begin
      ex_reg_fp_wen <= T152;
    end
    if(ctrl_killm) begin
      wb_reg_mem_val <= 1'h0;
    end else begin
      wb_reg_mem_val <= mem_reg_mem_val;
    end
    if(ctrl_killx) begin
      mem_reg_mem_val <= 1'h0;
    end else begin
      mem_reg_mem_val <= ex_reg_mem_val;
    end
    if(reset) begin
      R208 <= 32'h0;
    end else if(T222) begin
      R208 <= T211;
    end else if(io_dpath_ll_wen) begin
      R208 <= T204;
    end
    if(ctrl_killm) begin
      wb_reg_div_mul_val <= 1'h0;
    end else begin
      wb_reg_div_mul_val <= mem_reg_div_mul_val;
    end
    mem_reg_div_mul_val <= T217;
    if(ctrl_killd) begin
      ex_reg_div_mul_val <= 1'h0;
    end else begin
      ex_reg_div_mul_val <= T219;
    end
    if(ctrl_killm) begin
      wb_reg_fp_val <= 1'h0;
    end else begin
      wb_reg_fp_val <= mem_reg_fp_val;
    end
    if(ctrl_killm) begin
      wb_reg_wen <= 1'h0;
    end else begin
      wb_reg_wen <= mem_reg_wen;
    end
    if(T352) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T320) begin
      ex_reg_mem_type <= T312;
    end
    if(T320) begin
      ex_reg_mem_cmd <= id_mem_cmd;
    end
    if(ctrl_killx) begin
      mem_reg_csr <= 2'h0;
    end else begin
      mem_reg_csr <= ex_reg_csr;
    end
    if(ctrl_killd) begin
      ex_reg_csr <= 2'h0;
    end else begin
      ex_reg_csr <= id_csr;
    end
    if(ctrl_killd) begin
      ex_reg_jalr <= 1'h0;
    end else begin
      ex_reg_jalr <= id_jalr;
    end
    if(ctrl_killx) begin
      mem_reg_jal <= 1'h0;
    end else begin
      mem_reg_jal <= ex_reg_jal;
    end
    if(ctrl_killd) begin
      ex_reg_jal <= 1'h0;
    end else begin
      ex_reg_jal <= id_jal;
    end
    if(ctrl_killx) begin
      mem_reg_jalr <= 1'h0;
    end else begin
      mem_reg_jalr <= ex_reg_jalr;
    end
    if(ctrl_killx) begin
      mem_reg_branch <= 1'h0;
    end else begin
      mem_reg_branch <= ex_reg_branch;
    end
    if(ctrl_killd) begin
      ex_reg_branch <= 1'h0;
    end else begin
      ex_reg_branch <= id_branch;
    end
    if(ctrl_killd) begin
      ex_reg_load_use <= 1'h0;
    end else begin
      ex_reg_load_use <= id_load_use;
    end
    if(ctrl_killx) begin
      mem_reg_sret <= 1'h0;
    end else begin
      mem_reg_sret <= ex_reg_sret;
    end
    if(ctrl_killd) begin
      ex_reg_sret <= 1'h0;
    end else begin
      ex_reg_sret <= id_sret;
    end
    if(ctrl_killx) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ex_reg_valid;
    end
    if(ctrl_killd) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= 1'h1;
    end
    if(ctrl_killx) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ex_xcpt;
    end
    if(ctrl_killd) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= id_xcpt;
    end
    ex_reg_xcpt_interrupt <= T566;
    mem_reg_xcpt_interrupt <= T579;
    if(ctrl_killm) begin
      wb_reg_flush_inst <= 1'h0;
    end else begin
      wb_reg_flush_inst <= mem_reg_flush_inst;
    end
    if(ctrl_killx) begin
      mem_reg_flush_inst <= 1'h0;
    end else begin
      mem_reg_flush_inst <= ex_reg_flush_inst;
    end
    if(ctrl_killd) begin
      ex_reg_flush_inst <= 1'h0;
    end else begin
      ex_reg_flush_inst <= id_fence_i;
    end
    if(T599) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T598) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(ctrl_killd) begin
      ex_reg_btb_hit <= 1'h0;
    end else begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T599) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T598) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T599) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T598) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T599) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T598) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T599) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T598) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T352) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(ctrl_killm) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= mem_reg_valid;
    end
    if(ctrl_killm) begin
      wb_reg_csr <= 2'h0;
    end else begin
      wb_reg_csr <= mem_reg_csr;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T133;
  wire cmp;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] T29;
  wire T30;
  wire[63:0] shout_l;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[62:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[61:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[59:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[55:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[47:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T134;
  wire[31:0] T55;
  wire[63:0] T56;
  wire[63:0] T135;
  wire[47:0] T57;
  wire[63:0] T58;
  wire[63:0] T136;
  wire[55:0] T59;
  wire[63:0] T60;
  wire[63:0] T137;
  wire[59:0] T61;
  wire[63:0] T62;
  wire[63:0] T138;
  wire[61:0] T63;
  wire[63:0] T64;
  wire[63:0] T139;
  wire[62:0] T65;
  wire T66;
  wire[63:0] shout_r;
  wire[64:0] T67;
  wire[5:0] shamt;
  wire[5:0] T68;
  wire[4:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[64:0] T73;
  wire[64:0] T74;
  wire[63:0] shin;
  wire[63:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[62:0] T78;
  wire[63:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[61:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[59:0] T86;
  wire[63:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[55:0] T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[47:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[31:0] T98;
  wire[63:0] T99;
  wire[63:0] T140;
  wire[31:0] T100;
  wire[63:0] T101;
  wire[63:0] T141;
  wire[47:0] T102;
  wire[63:0] T103;
  wire[63:0] T142;
  wire[55:0] T104;
  wire[63:0] T105;
  wire[63:0] T143;
  wire[59:0] T106;
  wire[63:0] T107;
  wire[63:0] T144;
  wire[61:0] T108;
  wire[63:0] T109;
  wire[63:0] T145;
  wire[62:0] T110;
  wire[63:0] shin_r;
  wire[31:0] T111;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T112;
  wire[31:0] T146;
  wire T113;
  wire T114;
  wire[31:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[31:0] out_hi;
  wire[31:0] T129;
  wire[31:0] T147;
  wire T130;
  wire[31:0] T131;
  wire T132;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T126 ? sum : T6;
  assign T6 = T123 ? shout_r : T7;
  assign T7 = T66 ? shout_l : T8;
  assign T8 = T30 ? T29 : T9;
  assign T9 = T28 ? T27 : T10;
  assign T10 = T26 ? T25 : T133;
  assign T133 = {63'h0, cmp};
  assign cmp = T24 ^ T11;
  assign T11 = T22 ? T21 : T12;
  assign T12 = T18 ? T17 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = io_in1[6'h3f:6'h3f];
  assign T15 = io_in2[6'h3f:6'h3f];
  assign T16 = io_fn[1'h1:1'h1];
  assign T17 = sum[6'h3f:6'h3f];
  assign T18 = T20 == T19;
  assign T19 = io_in2[6'h3f:6'h3f];
  assign T20 = io_in1[6'h3f:6'h3f];
  assign T21 = sum == 64'h0;
  assign T22 = T23 ^ 1'h1;
  assign T23 = io_fn[2'h2:2'h2];
  assign T24 = io_fn[1'h0:1'h0];
  assign T25 = io_in1 ^ io_in2;
  assign T26 = io_fn == 4'h4;
  assign T27 = io_in1 | io_in2;
  assign T28 = io_fn == 4'h6;
  assign T29 = io_in1 & io_in2;
  assign T30 = io_fn == 4'h7;
  assign shout_l = T64 | T31;
  assign T31 = T32 & 64'haaaaaaaaaaaaaaaa;
  assign T32 = T33 << 1'h1;
  assign T33 = T34[6'h3e:1'h0];
  assign T34 = T62 | T35;
  assign T35 = T36 & 64'hcccccccccccccccc;
  assign T36 = T37 << 2'h2;
  assign T37 = T38[6'h3d:1'h0];
  assign T38 = T60 | T39;
  assign T39 = T40 & 64'hf0f0f0f0f0f0f0f0;
  assign T40 = T41 << 3'h4;
  assign T41 = T42[6'h3b:1'h0];
  assign T42 = T58 | T43;
  assign T43 = T44 & 64'hff00ff00ff00ff00;
  assign T44 = T45 << 4'h8;
  assign T45 = T46[6'h37:1'h0];
  assign T46 = T56 | T47;
  assign T47 = T48 & 64'hffff0000ffff0000;
  assign T48 = T49 << 5'h10;
  assign T49 = T50[6'h2f:1'h0];
  assign T50 = T54 | T51;
  assign T51 = T52 & 64'hffffffff00000000;
  assign T52 = T53 << 6'h20;
  assign T53 = shout_r[5'h1f:1'h0];
  assign T54 = T134 & 64'hffffffff;
  assign T134 = {32'h0, T55};
  assign T55 = shout_r >> 6'h20;
  assign T56 = T135 & 64'hffff0000ffff;
  assign T135 = {16'h0, T57};
  assign T57 = T50 >> 5'h10;
  assign T58 = T136 & 64'hff00ff00ff00ff;
  assign T136 = {8'h0, T59};
  assign T59 = T46 >> 4'h8;
  assign T60 = T137 & 64'hf0f0f0f0f0f0f0f;
  assign T137 = {4'h0, T61};
  assign T61 = T42 >> 3'h4;
  assign T62 = T138 & 64'h3333333333333333;
  assign T138 = {2'h0, T63};
  assign T63 = T38 >> 2'h2;
  assign T64 = T139 & 64'h5555555555555555;
  assign T139 = {1'h0, T65};
  assign T65 = T34 >> 1'h1;
  assign T66 = io_fn == 4'h1;
  assign shout_r = T67[6'h3f:1'h0];
  assign T67 = $signed(T73) >>> shamt;
  assign shamt = T68;
  assign T68 = {T70, T69};
  assign T69 = io_in2[3'h4:1'h0];
  assign T70 = T72 & T71;
  assign T71 = io_dw == 1'h1;
  assign T72 = io_in2[3'h5:3'h5];
  assign T73 = T74;
  assign T74 = {T120, shin};
  assign shin = T117 ? shin_r : T75;
  assign T75 = T109 | T76;
  assign T76 = T77 & 64'haaaaaaaaaaaaaaaa;
  assign T77 = T78 << 1'h1;
  assign T78 = T79[6'h3e:1'h0];
  assign T79 = T107 | T80;
  assign T80 = T81 & 64'hcccccccccccccccc;
  assign T81 = T82 << 2'h2;
  assign T82 = T83[6'h3d:1'h0];
  assign T83 = T105 | T84;
  assign T84 = T85 & 64'hf0f0f0f0f0f0f0f0;
  assign T85 = T86 << 3'h4;
  assign T86 = T87[6'h3b:1'h0];
  assign T87 = T103 | T88;
  assign T88 = T89 & 64'hff00ff00ff00ff00;
  assign T89 = T90 << 4'h8;
  assign T90 = T91[6'h37:1'h0];
  assign T91 = T101 | T92;
  assign T92 = T93 & 64'hffff0000ffff0000;
  assign T93 = T94 << 5'h10;
  assign T94 = T95[6'h2f:1'h0];
  assign T95 = T99 | T96;
  assign T96 = T97 & 64'hffffffff00000000;
  assign T97 = T98 << 6'h20;
  assign T98 = shin_r[5'h1f:1'h0];
  assign T99 = T140 & 64'hffffffff;
  assign T140 = {32'h0, T100};
  assign T100 = shin_r >> 6'h20;
  assign T101 = T141 & 64'hffff0000ffff;
  assign T141 = {16'h0, T102};
  assign T102 = T95 >> 5'h10;
  assign T103 = T142 & 64'hff00ff00ff00ff;
  assign T142 = {8'h0, T104};
  assign T104 = T91 >> 4'h8;
  assign T105 = T143 & 64'hf0f0f0f0f0f0f0f;
  assign T143 = {4'h0, T106};
  assign T106 = T87 >> 3'h4;
  assign T107 = T144 & 64'h3333333333333333;
  assign T144 = {2'h0, T108};
  assign T108 = T83 >> 2'h2;
  assign T109 = T145 & 64'h5555555555555555;
  assign T145 = {1'h0, T110};
  assign T110 = T79 >> 1'h1;
  assign shin_r = {shin_hi, T111};
  assign T111 = io_in1[5'h1f:1'h0];
  assign shin_hi = T116 ? T115 : shin_hi_32;
  assign shin_hi_32 = T114 ? T112 : 32'h0;
  assign T112 = 32'h0 - T146;
  assign T146 = {31'h0, T113};
  assign T113 = io_in1[5'h1f:5'h1f];
  assign T114 = io_fn[2'h3:2'h3];
  assign T115 = io_in1[6'h3f:6'h20];
  assign T116 = io_dw == 1'h1;
  assign T117 = T119 | T118;
  assign T118 = io_fn == 4'hb;
  assign T119 = io_fn == 4'h5;
  assign T120 = T122 & T121;
  assign T121 = shin[6'h3f:6'h3f];
  assign T122 = io_fn[2'h3:2'h3];
  assign T123 = T125 | T124;
  assign T124 = io_fn == 4'hb;
  assign T125 = io_fn == 4'h5;
  assign T126 = T128 | T127;
  assign T127 = io_fn == 4'ha;
  assign T128 = io_fn == 4'h0;
  assign out_hi = T132 ? T131 : T129;
  assign T129 = 32'h0 - T147;
  assign T147 = {31'h0, T130};
  assign T130 = out64[5'h1f:5'h1f];
  assign T131 = out64[6'h3f:6'h20];
  assign T132 = io_dw == 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[129:0] T180;
  wire[63:0] negated_remainder;
  wire[63:0] T119;
  wire T11;
  wire T12;
  reg  isMul;
  wire T13;
  wire cmdMul;
  wire T14;
  wire[3:0] T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  reg [2:0] state;
  wire[2:0] T181;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  reg  neg_out;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  isHi;
  wire T33;
  wire cmdHi;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire T37;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T41;
  wire[64:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[64:0] T46;
  wire[63:0] rhs_in;
  wire[31:0] T47;
  wire[31:0] T48;
  wire[31:0] T49;
  wire[31:0] T182;
  wire[31:0] T50;
  wire T51;
  wire rhs_sign;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire rhsSigned;
  wire T56;
  wire[3:0] T57;
  wire[64:0] T58;
  wire T59;
  reg [6:0] count;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire[6:0] T65;
  wire[6:0] T183;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[5:0] T184;
  wire[5:0] T185;
  wire[5:0] T186;
  wire[5:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[5:0] T190;
  wire[5:0] T191;
  wire[5:0] T192;
  wire[5:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire[5:0] T196;
  wire[5:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[4:0] T216;
  wire[4:0] T217;
  wire[4:0] T218;
  wire[4:0] T219;
  wire[4:0] T220;
  wire[4:0] T221;
  wire[4:0] T222;
  wire[4:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[4:0] T226;
  wire[4:0] T227;
  wire[4:0] T228;
  wire[4:0] T229;
  wire[4:0] T230;
  wire[4:0] T231;
  wire[3:0] T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[3:0] T238;
  wire[3:0] T239;
  wire[2:0] T240;
  wire[2:0] T241;
  wire[2:0] T242;
  wire[2:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire T246;
  wire[63:0] T70;
  wire[63:0] T71;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire[5:0] T72;
  wire[5:0] T309;
  wire[5:0] T310;
  wire[5:0] T311;
  wire[5:0] T312;
  wire[5:0] T313;
  wire[5:0] T314;
  wire[5:0] T315;
  wire[5:0] T316;
  wire[5:0] T317;
  wire[5:0] T318;
  wire[5:0] T319;
  wire[5:0] T320;
  wire[5:0] T321;
  wire[5:0] T322;
  wire[5:0] T323;
  wire[5:0] T324;
  wire[5:0] T325;
  wire[5:0] T326;
  wire[5:0] T327;
  wire[5:0] T328;
  wire[5:0] T329;
  wire[5:0] T330;
  wire[5:0] T331;
  wire[5:0] T332;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[4:0] T341;
  wire[4:0] T342;
  wire[4:0] T343;
  wire[4:0] T344;
  wire[4:0] T345;
  wire[4:0] T346;
  wire[4:0] T347;
  wire[4:0] T348;
  wire[4:0] T349;
  wire[4:0] T350;
  wire[4:0] T351;
  wire[4:0] T352;
  wire[4:0] T353;
  wire[4:0] T354;
  wire[4:0] T355;
  wire[4:0] T356;
  wire[3:0] T357;
  wire[3:0] T358;
  wire[3:0] T359;
  wire[3:0] T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[2:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire T371;
  wire[63:0] T74;
  wire[63:0] T75;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire lhs_sign;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire lhsSigned;
  wire T84;
  wire[3:0] T85;
  wire T86;
  wire T87;
  wire[2:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[64:0] T97;
  wire[5:0] T98;
  wire[10:0] T99;
  wire[63:0] T100;
  wire[128:0] T101;
  wire[63:0] T102;
  wire[64:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire[129:0] T434;
  wire T120;
  wire[129:0] T435;
  wire[63:0] T121;
  wire T122;
  wire[129:0] T123;
  wire[129:0] T124;
  wire[64:0] T125;
  wire[63:0] T126;
  wire[128:0] T127;
  wire[63:0] T128;
  wire[128:0] T129;
  wire[128:0] T130;
  wire[128:0] T131;
  wire[55:0] T132;
  wire[72:0] T133;
  wire[72:0] T436;
  wire[64:0] T134;
  wire[64:0] T135;
  wire[7:0] T437;
  wire T438;
  wire[72:0] T136;
  wire[8:0] T137;
  wire[8:0] T138;
  wire[7:0] T139;
  wire[64:0] T140;
  wire[128:0] T141;
  wire[5:0] T142;
  wire[10:0] T143;
  wire[10:0] T144;
  wire[64:0] T145;
  wire[64:0] T146;
  wire T147;
  wire T148;
  wire[129:0] T439;
  wire[128:0] T149;
  wire[64:0] T150;
  wire T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[63:0] T154;
  wire[63:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[129:0] T440;
  wire[126:0] T159;
  wire[63:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire[129:0] T441;
  wire[63:0] lhs_in;
  wire[31:0] T167;
  wire[31:0] T168;
  wire[31:0] T169;
  wire[31:0] T442;
  wire[31:0] T170;
  wire T171;
  wire[63:0] T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T443;
  wire T175;
  wire T176;
  reg  req_dw;
  wire T177;
  wire T178;
  wire T179;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T176 ? T172 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T441 : T5;
  assign T5 = T161 ? T440 : T6;
  assign T6 = T156 ? T439 : T7;
  assign T7 = T147 ? T123 : T8;
  assign T8 = T122 ? T435 : T9;
  assign T9 = T120 ? T434 : T10;
  assign T10 = T11 ? T180 : remainder;
  assign T180 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T119;
  assign T119 = remainder[6'h3f:1'h0];
  assign T11 = T19 & T12;
  assign T12 = T18 | isMul;
  assign T13 = T1 ? cmdMul : isMul;
  assign cmdMul = T16 | T14;
  assign T14 = T15 == 4'h8;
  assign T15 = io_req_bits_fn & 4'h8;
  assign T16 = T17 == 4'h0;
  assign T17 = io_req_bits_fn & 4'h4;
  assign T18 = remainder[6'h3f:6'h3f];
  assign T19 = state == 3'h1;
  assign T181 = reset ? 3'h0 : T20;
  assign T20 = T1 ? T115 : T21;
  assign T21 = T113 ? 3'h0 : T22;
  assign T22 = T111 ? T109 : T23;
  assign T23 = T89 ? T88 : T24;
  assign T24 = T122 ? T27 : T25;
  assign T25 = T120 ? 3'h5 : T26;
  assign T26 = T19 ? 3'h2 : state;
  assign T27 = neg_out ? 3'h4 : 3'h5;
  assign T28 = T1 ? T77 : T29;
  assign T29 = T30 ? 1'h0 : neg_out;
  assign T30 = T156 & T31;
  assign T31 = T39 & T32;
  assign T32 = isHi ^ 1'h1;
  assign T33 = T1 ? cmdHi : isHi;
  assign cmdHi = T34 | T14;
  assign T34 = T37 | T35;
  assign T35 = T36 == 4'h2;
  assign T36 = io_req_bits_fn & 4'h2;
  assign T37 = T38 == 4'h1;
  assign T38 = io_req_bits_fn & 4'h5;
  assign T39 = T59 & T40;
  assign T40 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T58 - divisor;
  assign T41 = T1 ? T46 : T42;
  assign T42 = T43 ? subtractor : divisor;
  assign T43 = T19 & T44;
  assign T44 = T45 | isMul;
  assign T45 = divisor[6'h3f:6'h3f];
  assign T46 = {rhs_sign, rhs_in};
  assign rhs_in = {T48, T47};
  assign T47 = io_req_bits_in2[5'h1f:1'h0];
  assign T48 = T51 ? T50 : T49;
  assign T49 = 32'h0 - T182;
  assign T182 = {31'h0, rhs_sign};
  assign T50 = io_req_bits_in2[6'h3f:6'h20];
  assign T51 = io_req_bits_dw == 1'h1;
  assign rhs_sign = rhsSigned & T52;
  assign T52 = T55 ? T54 : T53;
  assign T53 = io_req_bits_in2[5'h1f:5'h1f];
  assign T54 = io_req_bits_in2[6'h3f:6'h3f];
  assign T55 = io_req_bits_dw == 1'h1;
  assign rhsSigned = T56 | T16;
  assign T56 = T57 == 4'h0;
  assign T57 = io_req_bits_fn & 4'h9;
  assign T58 = remainder[8'h80:7'h40];
  assign T59 = count == 7'h0;
  assign T60 = T1 ? 7'h0 : T61;
  assign T61 = T161 ? T183 : T62;
  assign T62 = T156 ? T65 : T63;
  assign T63 = T147 ? T64 : count;
  assign T64 = count + 7'h1;
  assign T65 = count + 7'h1;
  assign T183 = {1'h0, T66};
  assign T66 = T76 ? 6'h3f : T67;
  assign T67 = T68[3'h5:1'h0];
  assign T68 = T72 - T184;
  assign T184 = T308 ? 6'h3f : T185;
  assign T185 = T307 ? 6'h3e : T186;
  assign T186 = T306 ? 6'h3d : T187;
  assign T187 = T305 ? 6'h3c : T188;
  assign T188 = T304 ? 6'h3b : T189;
  assign T189 = T303 ? 6'h3a : T190;
  assign T190 = T302 ? 6'h39 : T191;
  assign T191 = T301 ? 6'h38 : T192;
  assign T192 = T300 ? 6'h37 : T193;
  assign T193 = T299 ? 6'h36 : T194;
  assign T194 = T298 ? 6'h35 : T195;
  assign T195 = T297 ? 6'h34 : T196;
  assign T196 = T296 ? 6'h33 : T197;
  assign T197 = T295 ? 6'h32 : T198;
  assign T198 = T294 ? 6'h31 : T199;
  assign T199 = T293 ? 6'h30 : T200;
  assign T200 = T292 ? 6'h2f : T201;
  assign T201 = T291 ? 6'h2e : T202;
  assign T202 = T290 ? 6'h2d : T203;
  assign T203 = T289 ? 6'h2c : T204;
  assign T204 = T288 ? 6'h2b : T205;
  assign T205 = T287 ? 6'h2a : T206;
  assign T206 = T286 ? 6'h29 : T207;
  assign T207 = T285 ? 6'h28 : T208;
  assign T208 = T284 ? 6'h27 : T209;
  assign T209 = T283 ? 6'h26 : T210;
  assign T210 = T282 ? 6'h25 : T211;
  assign T211 = T281 ? 6'h24 : T212;
  assign T212 = T280 ? 6'h23 : T213;
  assign T213 = T279 ? 6'h22 : T214;
  assign T214 = T278 ? 6'h21 : T215;
  assign T215 = T277 ? 6'h20 : T216;
  assign T216 = T276 ? 5'h1f : T217;
  assign T217 = T275 ? 5'h1e : T218;
  assign T218 = T274 ? 5'h1d : T219;
  assign T219 = T273 ? 5'h1c : T220;
  assign T220 = T272 ? 5'h1b : T221;
  assign T221 = T271 ? 5'h1a : T222;
  assign T222 = T270 ? 5'h19 : T223;
  assign T223 = T269 ? 5'h18 : T224;
  assign T224 = T268 ? 5'h17 : T225;
  assign T225 = T267 ? 5'h16 : T226;
  assign T226 = T266 ? 5'h15 : T227;
  assign T227 = T265 ? 5'h14 : T228;
  assign T228 = T264 ? 5'h13 : T229;
  assign T229 = T263 ? 5'h12 : T230;
  assign T230 = T262 ? 5'h11 : T231;
  assign T231 = T261 ? 5'h10 : T232;
  assign T232 = T260 ? 4'hf : T233;
  assign T233 = T259 ? 4'he : T234;
  assign T234 = T258 ? 4'hd : T235;
  assign T235 = T257 ? 4'hc : T236;
  assign T236 = T256 ? 4'hb : T237;
  assign T237 = T255 ? 4'ha : T238;
  assign T238 = T254 ? 4'h9 : T239;
  assign T239 = T253 ? 4'h8 : T240;
  assign T240 = T252 ? 3'h7 : T241;
  assign T241 = T251 ? 3'h6 : T242;
  assign T242 = T250 ? 3'h5 : T243;
  assign T243 = T249 ? 3'h4 : T244;
  assign T244 = T248 ? 2'h3 : T245;
  assign T245 = T247 ? 2'h2 : T246;
  assign T246 = T70[1'h1:1'h1];
  assign T70 = T71[6'h3f:1'h0];
  assign T71 = remainder[6'h3f:1'h0];
  assign T247 = T70[2'h2:2'h2];
  assign T248 = T70[2'h3:2'h3];
  assign T249 = T70[3'h4:3'h4];
  assign T250 = T70[3'h5:3'h5];
  assign T251 = T70[3'h6:3'h6];
  assign T252 = T70[3'h7:3'h7];
  assign T253 = T70[4'h8:4'h8];
  assign T254 = T70[4'h9:4'h9];
  assign T255 = T70[4'ha:4'ha];
  assign T256 = T70[4'hb:4'hb];
  assign T257 = T70[4'hc:4'hc];
  assign T258 = T70[4'hd:4'hd];
  assign T259 = T70[4'he:4'he];
  assign T260 = T70[4'hf:4'hf];
  assign T261 = T70[5'h10:5'h10];
  assign T262 = T70[5'h11:5'h11];
  assign T263 = T70[5'h12:5'h12];
  assign T264 = T70[5'h13:5'h13];
  assign T265 = T70[5'h14:5'h14];
  assign T266 = T70[5'h15:5'h15];
  assign T267 = T70[5'h16:5'h16];
  assign T268 = T70[5'h17:5'h17];
  assign T269 = T70[5'h18:5'h18];
  assign T270 = T70[5'h19:5'h19];
  assign T271 = T70[5'h1a:5'h1a];
  assign T272 = T70[5'h1b:5'h1b];
  assign T273 = T70[5'h1c:5'h1c];
  assign T274 = T70[5'h1d:5'h1d];
  assign T275 = T70[5'h1e:5'h1e];
  assign T276 = T70[5'h1f:5'h1f];
  assign T277 = T70[6'h20:6'h20];
  assign T278 = T70[6'h21:6'h21];
  assign T279 = T70[6'h22:6'h22];
  assign T280 = T70[6'h23:6'h23];
  assign T281 = T70[6'h24:6'h24];
  assign T282 = T70[6'h25:6'h25];
  assign T283 = T70[6'h26:6'h26];
  assign T284 = T70[6'h27:6'h27];
  assign T285 = T70[6'h28:6'h28];
  assign T286 = T70[6'h29:6'h29];
  assign T287 = T70[6'h2a:6'h2a];
  assign T288 = T70[6'h2b:6'h2b];
  assign T289 = T70[6'h2c:6'h2c];
  assign T290 = T70[6'h2d:6'h2d];
  assign T291 = T70[6'h2e:6'h2e];
  assign T292 = T70[6'h2f:6'h2f];
  assign T293 = T70[6'h30:6'h30];
  assign T294 = T70[6'h31:6'h31];
  assign T295 = T70[6'h32:6'h32];
  assign T296 = T70[6'h33:6'h33];
  assign T297 = T70[6'h34:6'h34];
  assign T298 = T70[6'h35:6'h35];
  assign T299 = T70[6'h36:6'h36];
  assign T300 = T70[6'h37:6'h37];
  assign T301 = T70[6'h38:6'h38];
  assign T302 = T70[6'h39:6'h39];
  assign T303 = T70[6'h3a:6'h3a];
  assign T304 = T70[6'h3b:6'h3b];
  assign T305 = T70[6'h3c:6'h3c];
  assign T306 = T70[6'h3d:6'h3d];
  assign T307 = T70[6'h3e:6'h3e];
  assign T308 = T70[6'h3f:6'h3f];
  assign T72 = 6'h3f + T309;
  assign T309 = T433 ? 6'h3f : T310;
  assign T310 = T432 ? 6'h3e : T311;
  assign T311 = T431 ? 6'h3d : T312;
  assign T312 = T430 ? 6'h3c : T313;
  assign T313 = T429 ? 6'h3b : T314;
  assign T314 = T428 ? 6'h3a : T315;
  assign T315 = T427 ? 6'h39 : T316;
  assign T316 = T426 ? 6'h38 : T317;
  assign T317 = T425 ? 6'h37 : T318;
  assign T318 = T424 ? 6'h36 : T319;
  assign T319 = T423 ? 6'h35 : T320;
  assign T320 = T422 ? 6'h34 : T321;
  assign T321 = T421 ? 6'h33 : T322;
  assign T322 = T420 ? 6'h32 : T323;
  assign T323 = T419 ? 6'h31 : T324;
  assign T324 = T418 ? 6'h30 : T325;
  assign T325 = T417 ? 6'h2f : T326;
  assign T326 = T416 ? 6'h2e : T327;
  assign T327 = T415 ? 6'h2d : T328;
  assign T328 = T414 ? 6'h2c : T329;
  assign T329 = T413 ? 6'h2b : T330;
  assign T330 = T412 ? 6'h2a : T331;
  assign T331 = T411 ? 6'h29 : T332;
  assign T332 = T410 ? 6'h28 : T333;
  assign T333 = T409 ? 6'h27 : T334;
  assign T334 = T408 ? 6'h26 : T335;
  assign T335 = T407 ? 6'h25 : T336;
  assign T336 = T406 ? 6'h24 : T337;
  assign T337 = T405 ? 6'h23 : T338;
  assign T338 = T404 ? 6'h22 : T339;
  assign T339 = T403 ? 6'h21 : T340;
  assign T340 = T402 ? 6'h20 : T341;
  assign T341 = T401 ? 5'h1f : T342;
  assign T342 = T400 ? 5'h1e : T343;
  assign T343 = T399 ? 5'h1d : T344;
  assign T344 = T398 ? 5'h1c : T345;
  assign T345 = T397 ? 5'h1b : T346;
  assign T346 = T396 ? 5'h1a : T347;
  assign T347 = T395 ? 5'h19 : T348;
  assign T348 = T394 ? 5'h18 : T349;
  assign T349 = T393 ? 5'h17 : T350;
  assign T350 = T392 ? 5'h16 : T351;
  assign T351 = T391 ? 5'h15 : T352;
  assign T352 = T390 ? 5'h14 : T353;
  assign T353 = T389 ? 5'h13 : T354;
  assign T354 = T388 ? 5'h12 : T355;
  assign T355 = T387 ? 5'h11 : T356;
  assign T356 = T386 ? 5'h10 : T357;
  assign T357 = T385 ? 4'hf : T358;
  assign T358 = T384 ? 4'he : T359;
  assign T359 = T383 ? 4'hd : T360;
  assign T360 = T382 ? 4'hc : T361;
  assign T361 = T381 ? 4'hb : T362;
  assign T362 = T380 ? 4'ha : T363;
  assign T363 = T379 ? 4'h9 : T364;
  assign T364 = T378 ? 4'h8 : T365;
  assign T365 = T377 ? 3'h7 : T366;
  assign T366 = T376 ? 3'h6 : T367;
  assign T367 = T375 ? 3'h5 : T368;
  assign T368 = T374 ? 3'h4 : T369;
  assign T369 = T373 ? 2'h3 : T370;
  assign T370 = T372 ? 2'h2 : T371;
  assign T371 = T74[1'h1:1'h1];
  assign T74 = T75[6'h3f:1'h0];
  assign T75 = divisor[6'h3f:1'h0];
  assign T372 = T74[2'h2:2'h2];
  assign T373 = T74[2'h3:2'h3];
  assign T374 = T74[3'h4:3'h4];
  assign T375 = T74[3'h5:3'h5];
  assign T376 = T74[3'h6:3'h6];
  assign T377 = T74[3'h7:3'h7];
  assign T378 = T74[4'h8:4'h8];
  assign T379 = T74[4'h9:4'h9];
  assign T380 = T74[4'ha:4'ha];
  assign T381 = T74[4'hb:4'hb];
  assign T382 = T74[4'hc:4'hc];
  assign T383 = T74[4'hd:4'hd];
  assign T384 = T74[4'he:4'he];
  assign T385 = T74[4'hf:4'hf];
  assign T386 = T74[5'h10:5'h10];
  assign T387 = T74[5'h11:5'h11];
  assign T388 = T74[5'h12:5'h12];
  assign T389 = T74[5'h13:5'h13];
  assign T390 = T74[5'h14:5'h14];
  assign T391 = T74[5'h15:5'h15];
  assign T392 = T74[5'h16:5'h16];
  assign T393 = T74[5'h17:5'h17];
  assign T394 = T74[5'h18:5'h18];
  assign T395 = T74[5'h19:5'h19];
  assign T396 = T74[5'h1a:5'h1a];
  assign T397 = T74[5'h1b:5'h1b];
  assign T398 = T74[5'h1c:5'h1c];
  assign T399 = T74[5'h1d:5'h1d];
  assign T400 = T74[5'h1e:5'h1e];
  assign T401 = T74[5'h1f:5'h1f];
  assign T402 = T74[6'h20:6'h20];
  assign T403 = T74[6'h21:6'h21];
  assign T404 = T74[6'h22:6'h22];
  assign T405 = T74[6'h23:6'h23];
  assign T406 = T74[6'h24:6'h24];
  assign T407 = T74[6'h25:6'h25];
  assign T408 = T74[6'h26:6'h26];
  assign T409 = T74[6'h27:6'h27];
  assign T410 = T74[6'h28:6'h28];
  assign T411 = T74[6'h29:6'h29];
  assign T412 = T74[6'h2a:6'h2a];
  assign T413 = T74[6'h2b:6'h2b];
  assign T414 = T74[6'h2c:6'h2c];
  assign T415 = T74[6'h2d:6'h2d];
  assign T416 = T74[6'h2e:6'h2e];
  assign T417 = T74[6'h2f:6'h2f];
  assign T418 = T74[6'h30:6'h30];
  assign T419 = T74[6'h31:6'h31];
  assign T420 = T74[6'h32:6'h32];
  assign T421 = T74[6'h33:6'h33];
  assign T422 = T74[6'h34:6'h34];
  assign T423 = T74[6'h35:6'h35];
  assign T424 = T74[6'h36:6'h36];
  assign T425 = T74[6'h37:6'h37];
  assign T426 = T74[6'h38:6'h38];
  assign T427 = T74[6'h39:6'h39];
  assign T428 = T74[6'h3a:6'h3a];
  assign T429 = T74[6'h3b:6'h3b];
  assign T430 = T74[6'h3c:6'h3c];
  assign T431 = T74[6'h3d:6'h3d];
  assign T432 = T74[6'h3e:6'h3e];
  assign T433 = T74[6'h3f:6'h3f];
  assign T76 = T184 < T309;
  assign T77 = T87 & T78;
  assign T78 = cmdHi ? lhs_sign : T79;
  assign T79 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T80;
  assign T80 = T83 ? T82 : T81;
  assign T81 = io_req_bits_in1[5'h1f:5'h1f];
  assign T82 = io_req_bits_in1[6'h3f:6'h3f];
  assign T83 = io_req_bits_dw == 1'h1;
  assign lhsSigned = T86 | T84;
  assign T84 = T85 == 4'h0;
  assign T85 = io_req_bits_fn & 4'h3;
  assign T86 = T56 | T16;
  assign T87 = cmdMul ^ 1'h1;
  assign T88 = isHi ? 3'h3 : 3'h5;
  assign T89 = T147 & T90;
  assign T90 = T92 | T91;
  assign T91 = count == 7'h7;
  assign T92 = T104 & T93;
  assign T93 = T94 == 64'h0;
  assign T94 = T100 & T95;
  assign T95 = ~ T96;
  assign T96 = T97[6'h3f:1'h0];
  assign T97 = $signed(65'h10000000000000000) >>> T98;
  assign T98 = T99[3'h5:1'h0];
  assign T99 = count * 4'h8;
  assign T100 = T101[6'h3f:1'h0];
  assign T101 = {T103, T102};
  assign T102 = remainder[6'h3f:1'h0];
  assign T103 = remainder[8'h81:7'h41];
  assign T104 = T106 & T105;
  assign T105 = isHi ^ 1'h1;
  assign T106 = T108 & T107;
  assign T107 = count != 7'h0;
  assign T108 = count != 7'h7;
  assign T109 = isHi ? 3'h3 : T110;
  assign T110 = neg_out ? 3'h4 : 3'h5;
  assign T111 = T156 & T112;
  assign T112 = count == 7'h40;
  assign T113 = T114 | io_kill;
  assign T114 = io_resp_ready & io_resp_valid;
  assign T115 = T116 ? 3'h1 : 3'h2;
  assign T116 = lhs_sign | T117;
  assign T117 = rhs_sign & T118;
  assign T118 = cmdMul ^ 1'h1;
  assign T434 = {66'h0, negated_remainder};
  assign T120 = state == 3'h4;
  assign T435 = {66'h0, T121};
  assign T121 = remainder[8'h80:7'h41];
  assign T122 = state == 3'h3;
  assign T123 = T124;
  assign T124 = {T146, T125};
  assign T125 = {1'h0, T126};
  assign T126 = T127[6'h3f:1'h0];
  assign T127 = {T145, T128};
  assign T128 = T129[6'h3f:1'h0];
  assign T129 = T92 ? T141 : T130;
  assign T130 = T131;
  assign T131 = {T133, T132};
  assign T132 = T100[6'h3f:4'h8];
  assign T133 = T136 + T436;
  assign T436 = {T437, T134};
  assign T134 = T135;
  assign T135 = T101[8'h80:7'h40];
  assign T437 = T438 ? 8'hff : 8'h0;
  assign T438 = T134[7'h40:7'h40];
  assign T136 = $signed(T140) * $signed(T137);
  assign T137 = T138;
  assign T138 = {1'h0, T139};
  assign T139 = T100[3'h7:1'h0];
  assign T140 = divisor;
  assign T141 = T101 >> T142;
  assign T142 = T143[3'h5:1'h0];
  assign T143 = 11'h40 - T144;
  assign T144 = count * 4'h8;
  assign T145 = T130[8'h80:7'h40];
  assign T146 = T127 >> 7'h40;
  assign T147 = T148 & isMul;
  assign T148 = state == 3'h2;
  assign T439 = {1'h0, T149};
  assign T149 = {T153, T150};
  assign T150 = {T152, T151};
  assign T151 = less ^ 1'h1;
  assign T152 = remainder[6'h3f:1'h0];
  assign T153 = less ? T155 : T154;
  assign T154 = subtractor[6'h3f:1'h0];
  assign T155 = remainder[7'h7f:7'h40];
  assign T156 = T158 & T157;
  assign T157 = isMul ^ 1'h1;
  assign T158 = state == 3'h2;
  assign T440 = {3'h0, T159};
  assign T159 = T160 << T66;
  assign T160 = remainder[6'h3f:1'h0];
  assign T161 = T156 & T162;
  assign T162 = T165 & T163;
  assign T163 = T164 | T76;
  assign T164 = 6'h0 < T68;
  assign T165 = T166 & less;
  assign T166 = count == 7'h0;
  assign T441 = {66'h0, lhs_in};
  assign lhs_in = {T168, T167};
  assign T167 = io_req_bits_in1[5'h1f:1'h0];
  assign T168 = T171 ? T170 : T169;
  assign T169 = 32'h0 - T442;
  assign T442 = {31'h0, lhs_sign};
  assign T170 = io_req_bits_in1[6'h3f:6'h20];
  assign T171 = io_req_bits_dw == 1'h1;
  assign T172 = {T174, T173};
  assign T173 = remainder[5'h1f:1'h0];
  assign T174 = 32'h0 - T443;
  assign T443 = {31'h0, T175};
  assign T175 = remainder[5'h1f:5'h1f];
  assign T176 = req_dw == 1'h0;
  assign T177 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T178;
  assign T178 = state == 3'h5;
  assign io_req_ready = T179;
  assign T179 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T441;
    end else if(T161) begin
      remainder <= T440;
    end else if(T156) begin
      remainder <= T439;
    end else if(T147) begin
      remainder <= T123;
    end else if(T122) begin
      remainder <= T435;
    end else if(T120) begin
      remainder <= T434;
    end else if(T11) begin
      remainder <= T180;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T115;
    end else if(T113) begin
      state <= 3'h0;
    end else if(T111) begin
      state <= T109;
    end else if(T89) begin
      state <= T88;
    end else if(T122) begin
      state <= T27;
    end else if(T120) begin
      state <= 3'h5;
    end else if(T19) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T77;
    end else if(T30) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T46;
    end else if(T43) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T161) begin
      count <= T183;
    end else if(T156) begin
      count <= T65;
    end else if(T147) begin
      count <= T64;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module ManagementMachine(input clk, input reset,
    output io_stall_out,
    input  io_write_to_cfga,
    input [63:0] io_cfgd_in,
    output io_s_axi_awvalid,
    input  io_s_axi_awready,
    output io_s_axi_wvalid,
    input  io_s_axi_wready,
    input [1:0] io_s_axi_bresp,
    input  io_s_axi_bvalid,
    output io_s_axi_bready,
    output io_s_axi_arvalid,
    //input  io_s_axi_arready
    input [31:0] io_s_axi_rdata,
    input [1:0] io_s_axi_rresp,
    input  io_s_axi_rvalid,
    output io_s_axi_rready
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T33;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  handled;
  wire T34;
  wire T29;
  wire T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    handled = {1{$random}};
  end
`endif

  assign io_s_axi_rready = 1'h0;
  assign io_s_axi_arvalid = 1'h0;
  assign io_s_axi_bready = T0;
  assign T0 = state == 2'h3;
  assign T33 = reset ? 2'h0 : T1;
  assign T1 = T16 ? 2'h0 : T2;
  assign T2 = T11 ? 2'h3 : T3;
  assign T3 = T7 ? 2'h2 : T4;
  assign T4 = T5 ? 2'h1 : 2'h0;
  assign T5 = T6 & io_write_to_cfga;
  assign T6 = state == 2'h0;
  assign T7 = T8 & io_s_axi_awready;
  assign T8 = T10 & T9;
  assign T9 = state == 2'h1;
  assign T10 = T6 ^ 1'h1;
  assign T11 = T12 & io_s_axi_wready;
  assign T12 = T14 & T13;
  assign T13 = state == 2'h2;
  assign T14 = T15 ^ 1'h1;
  assign T15 = T6 | T9;
  assign T16 = T17 & io_s_axi_bvalid;
  assign T17 = T19 & T18;
  assign T18 = state == 2'h3;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T15 | T13;
  assign io_s_axi_wvalid = T21;
  assign T21 = T23 & T22;
  assign T22 = io_cfgd_in[6'h20:6'h20];
  assign T23 = state == 2'h2;
  assign io_s_axi_awvalid = T24;
  assign T24 = T26 & T25;
  assign T25 = io_cfgd_in[6'h20:6'h20];
  assign T26 = state == 2'h1;
  assign io_stall_out = T27;
  assign T27 = T31 & T28;
  assign T28 = handled == 1'h0;
  assign T34 = reset ? 1'h0 : T29;
  assign T29 = T16 ? 1'h1 : T30;
  assign T30 = T6 ? 1'h0 : handled;
  assign T31 = T32 | io_write_to_cfga;
  assign T32 = state != 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T16) begin
      state <= 2'h0;
    end else if(T11) begin
      state <= 2'h3;
    end else if(T7) begin
      state <= 2'h2;
    end else if(T5) begin
      state <= 2'h1;
    end else begin
      state <= 2'h0;
    end
    if(reset) begin
      handled <= 1'h0;
    end else if(T16) begin
      handled <= 1'h1;
    end else if(T6) begin
      handled <= 1'h0;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [1:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready,
    output[7:0] io_status_ip,
    output[7:0] io_status_im,
    output[6:0] io_status_zero,
    output io_status_er,
    output io_status_vm,
    output io_status_s64,
    output io_status_u64,
    output io_status_ef,
    output io_status_pei,
    output io_status_ei,
    output io_status_ps,
    output io_status_s,
    output[31:0] io_ptbr,
    output[43:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input  io_badvaddr_wen,
    input [43:0] io_pc,
    input  io_sret,
    output io_fatc,
    output io_replay,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  reg [63:0] reg_cfgd;
  wire[63:0] T506;
  wire[63:0] T135;
  wire[63:0] wdata;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T2;
  wire[63:0] T3;
  wire T4;
  wire host_pcr_req_fire;
  wire T5;
  reg  host_pcr_req_valid;
  wire T6;
  wire T7;
  wire cpu_req_valid;
  wire T136;
  wire T137;
  reg [45:0] T10;
  wire[11:0] addr;
  wire[11:0] T494;
  wire[10:0] T12;
  wire[10:0] T495;
  reg [4:0] host_pcr_bits_addr;
  wire[4:0] T13;
  wire wen;
  wire T14;
  reg  host_pcr_bits_rw;
  wire T15;
  wire T132;
  wire T133;
  reg [2:0] reg_frm;
  wire[2:0] T492;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T493;
  wire T8;
  wire T9;
  wire[63:0] T496;
  wire[58:0] T16;
  wire T17;
  wire T18;
  wire[63:0] T19;
  reg [5:0] R20;
  wire[5:0] T497;
  wire[5:0] T21;
  wire[5:0] T22;
  wire[6:0] T23;
  wire[6:0] T498;
  wire[5:0] T24;
  wire[63:0] T25;
  wire T26;
  wire T27;
  reg [57:0] R28;
  wire[57:0] T499;
  wire[57:0] T29;
  wire[57:0] T30;
  wire[57:0] T31;
  wire T32;
  wire[57:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[43:0] T38;
  wire[43:0] T39;
  reg [43:0] reg_epc;
  wire[43:0] T40;
  wire[43:0] T41;
  wire[43:0] T42;
  wire[43:0] T43;
  wire[43:0] T44;
  wire T45;
  wire T46;
  wire[43:0] T500;
  wire[42:0] T47;
  reg [42:0] reg_evec;
  wire[42:0] T48;
  wire[42:0] T49;
  wire[42:0] T50;
  wire T51;
  wire T52;
  wire T501;
  reg [31:0] reg_ptbr;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[18:0] T56;
  wire T57;
  wire T58;
  reg  reg_status_s;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  reg_status_ps;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg  reg_status_ei;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  reg_status_pei;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg  reg_status_ef;
  wire T79;
  wire T80;
  wire T81;
  reg  reg_status_u64;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  reg  reg_status_s64;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  reg_status_vm;
  wire T90;
  wire T91;
  wire T92;
  reg  reg_status_er;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  reg [6:0] reg_status_zero;
  wire[6:0] T97;
  wire[6:0] T98;
  wire[6:0] T99;
  wire[6:0] T100;
  reg [7:0] reg_status_im;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[3:0] T105;
  wire[1:0] T106;
  reg  r_irq_ipi;
  wire T502;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[1:0] T112;
  wire T113;
  reg [63:0] reg_fromhost;
  wire[63:0] T503;
  wire[63:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg  r_irq_timer;
  wire T504;
  wire T121;
  wire T122;
  wire T123;
  reg [31:0] reg_compare;
  wire[31:0] T124;
  wire[31:0] T125;
  wire[31:0] T126;
  wire[31:0] T127;
  wire T128;
  wire T129;
  wire[11:0] T130;
  reg [63:0] reg_cfga;
  wire[63:0] T505;
  wire[63:0] T131;
  wire[31:0] T134;
  wire[11:0] T138;
  wire[63:0] T139;
  wire[63:0] T140;
  wire[63:0] T141;
  reg [5:0] R142;
  wire[5:0] T507;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[6:0] T145;
  wire[6:0] T508;
  wire T146;
  reg [57:0] R147;
  wire[57:0] T509;
  wire[57:0] T148;
  wire[57:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire[63:0] T153;
  wire[63:0] T154;
  wire[63:0] T155;
  reg [5:0] R156;
  wire[5:0] T510;
  wire[5:0] T157;
  wire[5:0] T158;
  wire[6:0] T159;
  wire[6:0] T511;
  wire T160;
  reg [57:0] R161;
  wire[57:0] T512;
  wire[57:0] T162;
  wire[57:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire[63:0] T167;
  wire[63:0] T168;
  wire[63:0] T169;
  reg [5:0] R170;
  wire[5:0] T513;
  wire[5:0] T171;
  wire[5:0] T172;
  wire[6:0] T173;
  wire[6:0] T514;
  wire T174;
  reg [57:0] R175;
  wire[57:0] T515;
  wire[57:0] T176;
  wire[57:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire[63:0] T181;
  wire[63:0] T182;
  wire[63:0] T183;
  reg [5:0] R184;
  wire[5:0] T516;
  wire[5:0] T185;
  wire[5:0] T186;
  wire[6:0] T187;
  wire[6:0] T517;
  wire T188;
  reg [57:0] R189;
  wire[57:0] T518;
  wire[57:0] T190;
  wire[57:0] T191;
  wire T192;
  wire T193;
  wire T194;
  wire[63:0] T195;
  wire[63:0] T196;
  wire[63:0] T197;
  reg [5:0] R198;
  wire[5:0] T519;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[6:0] T201;
  wire[6:0] T520;
  wire T202;
  reg [57:0] R203;
  wire[57:0] T521;
  wire[57:0] T204;
  wire[57:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire[63:0] T209;
  wire[63:0] T210;
  wire[63:0] T211;
  reg [5:0] R212;
  wire[5:0] T522;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[6:0] T215;
  wire[6:0] T523;
  wire T216;
  reg [57:0] R217;
  wire[57:0] T524;
  wire[57:0] T218;
  wire[57:0] T219;
  wire T220;
  wire T221;
  wire T222;
  wire[63:0] T223;
  wire[63:0] T224;
  wire[63:0] T225;
  reg [5:0] R226;
  wire[5:0] T525;
  wire[5:0] T227;
  wire[5:0] T228;
  wire[6:0] T229;
  wire[6:0] T526;
  wire T230;
  reg [57:0] R231;
  wire[57:0] T527;
  wire[57:0] T232;
  wire[57:0] T233;
  wire T234;
  wire T235;
  wire T236;
  wire[63:0] T237;
  wire[63:0] T238;
  wire[63:0] T239;
  reg [5:0] R240;
  wire[5:0] T528;
  wire[5:0] T241;
  wire[5:0] T242;
  wire[6:0] T243;
  wire[6:0] T529;
  wire T244;
  reg [57:0] R245;
  wire[57:0] T530;
  wire[57:0] T246;
  wire[57:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[63:0] T251;
  wire[63:0] T252;
  wire[63:0] T253;
  reg [5:0] R254;
  wire[5:0] T531;
  wire[5:0] T255;
  wire[5:0] T256;
  wire[6:0] T257;
  wire[6:0] T532;
  wire T258;
  reg [57:0] R259;
  wire[57:0] T533;
  wire[57:0] T260;
  wire[57:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire[63:0] T265;
  wire[63:0] T266;
  wire[63:0] T267;
  reg [5:0] R268;
  wire[5:0] T534;
  wire[5:0] T269;
  wire[5:0] T270;
  wire[6:0] T271;
  wire[6:0] T535;
  wire T272;
  reg [57:0] R273;
  wire[57:0] T536;
  wire[57:0] T274;
  wire[57:0] T275;
  wire T276;
  wire T277;
  wire T278;
  wire[63:0] T279;
  wire[63:0] T280;
  wire[63:0] T281;
  reg [5:0] R282;
  wire[5:0] T537;
  wire[5:0] T283;
  wire[5:0] T284;
  wire[6:0] T285;
  wire[6:0] T538;
  wire T286;
  reg [57:0] R287;
  wire[57:0] T539;
  wire[57:0] T288;
  wire[57:0] T289;
  wire T290;
  wire T291;
  wire T292;
  wire[63:0] T293;
  wire[63:0] T294;
  wire[63:0] T295;
  reg [5:0] R296;
  wire[5:0] T540;
  wire[5:0] T297;
  wire[5:0] T298;
  wire[6:0] T299;
  wire[6:0] T541;
  wire T300;
  reg [57:0] R301;
  wire[57:0] T542;
  wire[57:0] T302;
  wire[57:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[63:0] T307;
  wire[63:0] T308;
  wire[63:0] T309;
  reg [5:0] R310;
  wire[5:0] T543;
  wire[5:0] T311;
  wire[5:0] T312;
  wire[6:0] T313;
  wire[6:0] T544;
  wire T314;
  reg [57:0] R315;
  wire[57:0] T545;
  wire[57:0] T316;
  wire[57:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[63:0] T321;
  wire[63:0] T322;
  wire[63:0] T323;
  reg [5:0] R324;
  wire[5:0] T546;
  wire[5:0] T325;
  wire[5:0] T326;
  wire[6:0] T327;
  wire[6:0] T547;
  wire T328;
  reg [57:0] R329;
  wire[57:0] T548;
  wire[57:0] T330;
  wire[57:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire[63:0] T335;
  wire[63:0] T336;
  wire[63:0] T337;
  reg [5:0] R338;
  wire[5:0] T549;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[6:0] T341;
  wire[6:0] T550;
  wire T342;
  reg [57:0] R343;
  wire[57:0] T551;
  wire[57:0] T344;
  wire[57:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire[63:0] T349;
  wire[63:0] T350;
  wire[63:0] T351;
  reg [5:0] R352;
  wire[5:0] T552;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[6:0] T355;
  wire[6:0] T553;
  wire T356;
  reg [57:0] R357;
  wire[57:0] T554;
  wire[57:0] T358;
  wire[57:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[63:0] T363;
  wire[63:0] T364;
  wire[63:0] T365;
  wire[63:0] T366;
  wire[63:0] T367;
  wire[63:0] T368;
  wire[63:0] T369;
  wire[63:0] T370;
  reg [63:0] reg_tohost;
  wire[63:0] T555;
  wire[63:0] T371;
  wire[63:0] T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire[63:0] T381;
  wire[63:0] T556;
  wire T382;
  reg  reg_stats;
  wire T557;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire[63:0] T387;
  wire[63:0] T558;
  wire[1:0] T388;
  wire[63:0] T389;
  wire[63:0] T559;
  wire[1:0] T390;
  wire T391;
  wire[63:0] T392;
  wire[63:0] T560;
  wire[1:0] T393;
  wire[63:0] T394;
  wire[63:0] T561;
  wire[1:0] T395;
  wire T396;
  wire[63:0] T397;
  wire[63:0] T562;
  wire T398;
  wire T399;
  wire[63:0] T400;
  wire[63:0] T563;
  wire[31:0] T401;
  wire[31:0] T402;
  wire[31:0] T403;
  wire[5:0] T404;
  wire[2:0] T405;
  wire[1:0] T406;
  wire[2:0] T407;
  wire[1:0] T408;
  wire[25:0] T409;
  wire[2:0] T410;
  wire[1:0] T411;
  wire[22:0] T412;
  wire[14:0] T413;
  wire[63:0] T414;
  wire[63:0] T415;
  reg [63:0] reg_cause;
  wire[63:0] T416;
  wire T417;
  wire[63:0] T418;
  wire[63:0] T564;
  wire[42:0] T419;
  wire[63:0] T420;
  wire[63:0] T565;
  wire[31:0] T421;
  wire[63:0] T422;
  wire[63:0] T423;
  wire[63:0] T424;
  wire[63:0] T425;
  wire[63:0] T566;
  wire[31:0] T426;
  wire[31:0] read_ptbr;
  wire[18:0] T427;
  wire[63:0] T428;
  wire[63:0] T567;
  wire[42:0] T429;
  reg [42:0] reg_badvaddr;
  wire[42:0] T568;
  wire[43:0] T430;
  wire[43:0] T569;
  wire[43:0] T431;
  wire[43:0] T432;
  wire[42:0] T433;
  wire T434;
  wire T435;
  wire[20:0] T436;
  wire T437;
  wire T438;
  wire[42:0] T439;
  wire T440;
  wire[63:0] T441;
  wire[63:0] T570;
  wire[43:0] T442;
  wire[63:0] T443;
  wire[63:0] T444;
  reg [63:0] reg_sup1;
  wire[63:0] T445;
  wire T446;
  wire T447;
  wire[63:0] T448;
  wire[63:0] T449;
  reg [63:0] reg_sup0;
  wire[63:0] T450;
  wire T451;
  wire T452;
  wire[63:0] T453;
  wire[63:0] T454;
  wire[63:0] T455;
  reg [5:0] R456;
  wire[5:0] T571;
  wire[5:0] T457;
  wire[5:0] T458;
  wire[6:0] T459;
  wire[6:0] T572;
  wire T460;
  reg [57:0] R461;
  wire[57:0] T573;
  wire[57:0] T462;
  wire[57:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[63:0] T467;
  wire[63:0] T468;
  wire T469;
  wire[63:0] T470;
  wire[63:0] T471;
  wire T472;
  wire[63:0] T574;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  reg [4:0] reg_fflags;
  wire[4:0] T575;
  wire[63:0] T476;
  wire[63:0] T477;
  wire[63:0] T576;
  wire[4:0] T478;
  wire[4:0] T479;
  wire T480;
  wire T481;
  wire[7:0] T577;
  wire[4:0] T482;
  wire[4:0] T578;
  wire[2:0] T483;
  wire[4:0] T484;
  wire T579;
  wire T485;
  reg  host_pcr_rep_valid;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire temac_manage_io_s_axi_awvalid;
  wire temac_manage_io_s_axi_wvalid;
  wire temac_manage_io_s_axi_bready;
  wire temac_manage_io_s_axi_arvalid;
  wire temac_manage_io_s_axi_rready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    reg_cfgd = {2{$random}};
    host_pcr_bits_data = {2{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    reg_frm = {1{$random}};
    R20 = {1{$random}};
    R28 = {2{$random}};
    reg_epc = {2{$random}};
    reg_evec = {2{$random}};
    reg_ptbr = {1{$random}};
    reg_status_s = {1{$random}};
    reg_status_ps = {1{$random}};
    reg_status_ei = {1{$random}};
    reg_status_pei = {1{$random}};
    reg_status_ef = {1{$random}};
    reg_status_u64 = {1{$random}};
    reg_status_s64 = {1{$random}};
    reg_status_vm = {1{$random}};
    reg_status_er = {1{$random}};
    reg_status_zero = {1{$random}};
    reg_status_im = {1{$random}};
    r_irq_ipi = {1{$random}};
    reg_fromhost = {2{$random}};
    r_irq_timer = {1{$random}};
    reg_compare = {1{$random}};
    reg_cfga = {2{$random}};
    R142 = {1{$random}};
    R147 = {2{$random}};
    R156 = {1{$random}};
    R161 = {2{$random}};
    R170 = {1{$random}};
    R175 = {2{$random}};
    R184 = {1{$random}};
    R189 = {2{$random}};
    R198 = {1{$random}};
    R203 = {2{$random}};
    R212 = {1{$random}};
    R217 = {2{$random}};
    R226 = {1{$random}};
    R231 = {2{$random}};
    R240 = {1{$random}};
    R245 = {2{$random}};
    R254 = {1{$random}};
    R259 = {2{$random}};
    R268 = {1{$random}};
    R273 = {2{$random}};
    R282 = {1{$random}};
    R287 = {2{$random}};
    R296 = {1{$random}};
    R301 = {2{$random}};
    R310 = {1{$random}};
    R315 = {2{$random}};
    R324 = {1{$random}};
    R329 = {2{$random}};
    R338 = {1{$random}};
    R343 = {2{$random}};
    R352 = {1{$random}};
    R357 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_cause = {2{$random}};
    reg_badvaddr = {2{$random}};
    reg_sup1 = {2{$random}};
    reg_sup0 = {2{$random}};
    R456 = {1{$random}};
    R461 = {2{$random}};
    reg_fflags = {1{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
`endif

  assign T506 = reset ? 64'h0 : T135;
  assign T135 = T136 ? wdata : reg_cfgd;
  assign wdata = cpu_req_valid ? io_rw_wdata : host_pcr_bits_data;
  assign T2 = host_pcr_req_fire ? io_rw_rdata : T3;
  assign T3 = T4 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T4 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign host_pcr_req_fire = host_pcr_req_valid & T5;
  assign T5 = cpu_req_valid ^ 1'h1;
  assign T6 = host_pcr_req_fire ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : host_pcr_req_valid;
  assign cpu_req_valid = io_rw_cmd != 2'h0;
  assign T136 = wen & T137;
  assign T137 = T10[5'h1a:5'h1a];
  always @(*) case (addr)
    1: T10 = 46'h1;
    2: T10 = 46'h2;
    3: T10 = 46'h4;
    192: T10 = 46'h8;
    1280: T10 = 46'h10;
    1281: T10 = 46'h20;
    1282: T10 = 46'h40;
    1283: T10 = 46'h80;
    1284: T10 = 46'h100;
    1285: T10 = 46'h200;
    1286: T10 = 46'h400;
    1287: T10 = 46'h800;
    1288: T10 = 46'h1000;
    1289: T10 = 46'h2000;
    1290: T10 = 46'h4000;
    1291: T10 = 46'h8000;
    1292: T10 = 46'h10000;
    1293: T10 = 46'h20000;
    1294: T10 = 46'h40000;
    1295: T10 = 46'h80000;
    1309: T10 = 46'h100000;
    1310: T10 = 46'h200000;
    1311: T10 = 46'h400000;
    1312: T10 = 46'h800000;
    1313: T10 = 46'h1000000;
    1314: T10 = 46'h2000000;
    1315: T10 = 46'h4000000;
    3072: T10 = 46'h8000000;
    3073: T10 = 46'h10000000;
    3074: T10 = 46'h20000000;
    3264: T10 = 46'h40000000;
    3265: T10 = 46'h80000000;
    3266: T10 = 46'h100000000;
    3267: T10 = 46'h200000000;
    3268: T10 = 46'h400000000;
    3269: T10 = 46'h800000000;
    3270: T10 = 46'h1000000000;
    3271: T10 = 46'h2000000000;
    3272: T10 = 46'h4000000000;
    3273: T10 = 46'h8000000000;
    3274: T10 = 46'h10000000000;
    3275: T10 = 46'h20000000000;
    3276: T10 = 46'h40000000000;
    3277: T10 = 46'h80000000000;
    3278: T10 = 46'h100000000000;
    3279: T10 = 46'h200000000000;
`ifndef SYNTHESIS
    default: T10 = {2{$random}};
`else
    default: T10 = 46'bx;
`endif
  endcase
  assign addr = cpu_req_valid ? io_rw_addr : T494;
  assign T494 = {1'h0, T12};
  assign T12 = T495 | 11'h500;
  assign T495 = {6'h0, host_pcr_bits_addr};
  assign T13 = T4 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign wen = cpu_req_valid | T14;
  assign T14 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T15 = T4 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign T132 = wen & T133;
  assign T133 = T10[5'h19:5'h19];
  assign io_fcsr_rm = reg_frm;
  assign T492 = T0[2'h2:1'h0];
  assign T0 = T17 ? T496 : T1;
  assign T1 = T8 ? wdata : T493;
  assign T493 = {61'h0, reg_frm};
  assign T8 = wen & T9;
  assign T9 = T10[1'h1:1'h1];
  assign T496 = {5'h0, T16};
  assign T16 = wdata >> 3'h5;
  assign T17 = wen & T18;
  assign T18 = T10[2'h2:2'h2];
  assign io_time = T19;
  assign T19 = {R28, R20};
  assign T497 = reset ? 6'h0 : T21;
  assign T21 = T26 ? T24 : T22;
  assign T22 = T23[3'h5:1'h0];
  assign T23 = T498 + 7'h1;
  assign T498 = {1'h0, R20};
  assign T24 = T25[3'h5:1'h0];
  assign T25 = wdata;
  assign T26 = wen & T27;
  assign T27 = T10[4'ha:4'ha];
  assign T499 = reset ? 58'h0 : T29;
  assign T29 = T26 ? T33 : T30;
  assign T30 = T32 ? T31 : R28;
  assign T31 = R28 + 58'h1;
  assign T32 = T23[3'h6:3'h6];
  assign T33 = T25[6'h3f:3'h6];
  assign io_replay = T34;
  assign T34 = io_host_ipi_req_valid & T35;
  assign T35 = io_host_ipi_req_ready ^ 1'h1;
  assign io_fatc = T36;
  assign T36 = wen & T37;
  assign T37 = T10[5'h11:5'h11];
  assign io_evec = T38;
  assign T38 = T39;
  assign T39 = io_exception ? T500 : reg_epc;
  assign T40 = T45 ? T43 : T41;
  assign T41 = io_exception ? T42 : reg_epc;
  assign T42 = io_pc;
  assign T43 = T44;
  assign T44 = wdata[6'h2b:1'h0];
  assign T45 = wen & T46;
  assign T46 = T10[3'h6:3'h6];
  assign T500 = {T501, T47};
  assign T47 = reg_evec;
  assign T48 = T51 ? T49 : reg_evec;
  assign T49 = T50;
  assign T50 = wdata[6'h2a:1'h0];
  assign T51 = wen & T52;
  assign T52 = T10[4'hc:4'hc];
  assign T501 = T47[6'h2a:6'h2a];
  assign io_ptbr = reg_ptbr;
  assign T53 = T57 ? T54 : reg_ptbr;
  assign T54 = T55;
  assign T55 = {T56, 13'h0};
  assign T56 = wdata[5'h1f:4'hd];
  assign T57 = wen & T58;
  assign T58 = T10[4'h8:4'h8];
  assign io_status_s = reg_status_s;
  assign T59 = reset ? 1'h1 : T60;
  assign T60 = T68 ? T67 : T61;
  assign T61 = io_sret ? reg_status_ps : T62;
  assign T62 = io_exception ? 1'h1 : reg_status_s;
  assign T63 = reset ? 1'h0 : T64;
  assign T64 = T68 ? T66 : T65;
  assign T65 = io_exception ? reg_status_s : reg_status_ps;
  assign T66 = wdata[1'h1:1'h1];
  assign T67 = wdata[1'h0:1'h0];
  assign T68 = wen & T69;
  assign T69 = T10[4'he:4'he];
  assign io_status_ps = reg_status_ps;
  assign io_status_ei = reg_status_ei;
  assign T70 = reset ? 1'h0 : T71;
  assign T71 = T68 ? T78 : T72;
  assign T72 = io_sret ? reg_status_pei : T73;
  assign T73 = io_exception ? 1'h0 : reg_status_ei;
  assign T74 = reset ? 1'h0 : T75;
  assign T75 = T68 ? T77 : T76;
  assign T76 = io_exception ? reg_status_ei : reg_status_pei;
  assign T77 = wdata[2'h3:2'h3];
  assign T78 = wdata[2'h2:2'h2];
  assign io_status_pei = reg_status_pei;
  assign io_status_ef = reg_status_ef;
  assign T79 = reset ? 1'h0 : T80;
  assign T80 = T68 ? T81 : reg_status_ef;
  assign T81 = wdata[3'h4:3'h4];
  assign io_status_u64 = reg_status_u64;
  assign T82 = reset ? 1'h1 : T83;
  assign T83 = T68 ? 1'h1 : T84;
  assign T84 = T68 ? T85 : reg_status_u64;
  assign T85 = wdata[3'h5:3'h5];
  assign io_status_s64 = reg_status_s64;
  assign T86 = reset ? 1'h1 : T87;
  assign T87 = T68 ? 1'h1 : T88;
  assign T88 = T68 ? T89 : reg_status_s64;
  assign T89 = wdata[3'h6:3'h6];
  assign io_status_vm = reg_status_vm;
  assign T90 = reset ? 1'h0 : T91;
  assign T91 = T68 ? T92 : reg_status_vm;
  assign T92 = wdata[3'h7:3'h7];
  assign io_status_er = reg_status_er;
  assign T93 = reset ? 1'h0 : T94;
  assign T94 = T68 ? 1'h0 : T95;
  assign T95 = T68 ? T96 : reg_status_er;
  assign T96 = wdata[4'h8:4'h8];
  assign io_status_zero = reg_status_zero;
  assign T97 = reset ? 7'h0 : T98;
  assign T98 = T68 ? 7'h0 : T99;
  assign T99 = T68 ? T100 : reg_status_zero;
  assign T100 = wdata[4'hf:4'h9];
  assign io_status_im = reg_status_im;
  assign T101 = reset ? 8'h0 : T102;
  assign T102 = T68 ? T103 : reg_status_im;
  assign T103 = wdata[5'h17:5'h10];
  assign io_status_ip = T104;
  assign T104 = {T105, 4'h0};
  assign T105 = {T112, T106};
  assign T106 = {r_irq_ipi, 1'h0};
  assign T502 = reset ? 1'h1 : T107;
  assign T107 = io_host_ipi_rep_valid ? 1'h1 : T108;
  assign T108 = T110 ? T109 : r_irq_ipi;
  assign T109 = wdata[1'h0:1'h0];
  assign T110 = wen & T111;
  assign T111 = T10[5'h13:5'h13];
  assign T112 = {r_irq_timer, T113};
  assign T113 = reg_fromhost != 64'h0;
  assign T503 = reset ? 64'h0 : T114;
  assign T114 = T115 ? wdata : reg_fromhost;
  assign T115 = T119 & T116;
  assign T116 = T118 | T117;
  assign T117 = host_pcr_req_fire ^ 1'h1;
  assign T118 = reg_fromhost == 64'h0;
  assign T119 = wen & T120;
  assign T120 = T10[5'h16:5'h16];
  assign T504 = reset ? 1'h0 : T121;
  assign T121 = T128 ? 1'h0 : T122;
  assign T122 = T123 ? 1'h1 : r_irq_timer;
  assign T123 = T127 == reg_compare;
  assign T124 = T128 ? T125 : reg_compare;
  assign T125 = T126;
  assign T126 = wdata[5'h1f:1'h0];
  assign T127 = T19[5'h1f:1'h0];
  assign T128 = wen & T129;
  assign T129 = T10[4'hb:4'hb];
  assign io_temac_s_axi_rready = temac_manage_io_s_axi_rready;
  assign io_temac_s_axi_arvalid = temac_manage_io_s_axi_arvalid;
  assign io_temac_s_axi_araddr = T130;
  assign T130 = reg_cfga[4'hb:1'h0];
  assign T505 = reset ? 64'h0 : T131;
  assign T131 = T132 ? wdata : reg_cfga;
  assign io_temac_s_axi_bready = temac_manage_io_s_axi_bready;
  assign io_temac_s_axi_wvalid = temac_manage_io_s_axi_wvalid;
  assign io_temac_s_axi_wdata = T134;
  assign T134 = reg_cfgd[5'h1f:1'h0];
  assign io_temac_s_axi_awvalid = temac_manage_io_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = T138;
  assign T138 = reg_cfga[4'hb:1'h0];
  assign io_temac_tx_axis_fifo_tlast = 1'h0;
  assign io_temac_tx_axis_fifo_tvalid = 1'h0;
  assign io_temac_tx_axis_fifo_tdata = 8'hff;
  assign io_temac_rx_axis_fifo_tready = 1'h0;
  assign io_rw_rdata = T139;
  assign T139 = T153 | T140;
  assign T140 = T152 ? T141 : 64'h0;
  assign T141 = {R147, R142};
  assign T507 = reset ? 6'h0 : T143;
  assign T143 = T146 ? T144 : R142;
  assign T144 = T145[3'h5:1'h0];
  assign T145 = T508 + 7'h1;
  assign T508 = {1'h0, R142};
  assign T146 = io_uarch_counters_15 != 1'h0;
  assign T509 = reset ? 58'h0 : T148;
  assign T148 = T150 ? T149 : R147;
  assign T149 = R147 + 58'h1;
  assign T150 = T146 & T151;
  assign T151 = T145[3'h6:3'h6];
  assign T152 = T10[6'h2d:6'h2d];
  assign T153 = T167 | T154;
  assign T154 = T166 ? T155 : 64'h0;
  assign T155 = {R161, R156};
  assign T510 = reset ? 6'h0 : T157;
  assign T157 = T160 ? T158 : R156;
  assign T158 = T159[3'h5:1'h0];
  assign T159 = T511 + 7'h1;
  assign T511 = {1'h0, R156};
  assign T160 = io_uarch_counters_14 != 1'h0;
  assign T512 = reset ? 58'h0 : T162;
  assign T162 = T164 ? T163 : R161;
  assign T163 = R161 + 58'h1;
  assign T164 = T160 & T165;
  assign T165 = T159[3'h6:3'h6];
  assign T166 = T10[6'h2c:6'h2c];
  assign T167 = T181 | T168;
  assign T168 = T180 ? T169 : 64'h0;
  assign T169 = {R175, R170};
  assign T513 = reset ? 6'h0 : T171;
  assign T171 = T174 ? T172 : R170;
  assign T172 = T173[3'h5:1'h0];
  assign T173 = T514 + 7'h1;
  assign T514 = {1'h0, R170};
  assign T174 = io_uarch_counters_13 != 1'h0;
  assign T515 = reset ? 58'h0 : T176;
  assign T176 = T178 ? T177 : R175;
  assign T177 = R175 + 58'h1;
  assign T178 = T174 & T179;
  assign T179 = T173[3'h6:3'h6];
  assign T180 = T10[6'h2b:6'h2b];
  assign T181 = T195 | T182;
  assign T182 = T194 ? T183 : 64'h0;
  assign T183 = {R189, R184};
  assign T516 = reset ? 6'h0 : T185;
  assign T185 = T188 ? T186 : R184;
  assign T186 = T187[3'h5:1'h0];
  assign T187 = T517 + 7'h1;
  assign T517 = {1'h0, R184};
  assign T188 = io_uarch_counters_12 != 1'h0;
  assign T518 = reset ? 58'h0 : T190;
  assign T190 = T192 ? T191 : R189;
  assign T191 = R189 + 58'h1;
  assign T192 = T188 & T193;
  assign T193 = T187[3'h6:3'h6];
  assign T194 = T10[6'h2a:6'h2a];
  assign T195 = T209 | T196;
  assign T196 = T208 ? T197 : 64'h0;
  assign T197 = {R203, R198};
  assign T519 = reset ? 6'h0 : T199;
  assign T199 = T202 ? T200 : R198;
  assign T200 = T201[3'h5:1'h0];
  assign T201 = T520 + 7'h1;
  assign T520 = {1'h0, R198};
  assign T202 = io_uarch_counters_11 != 1'h0;
  assign T521 = reset ? 58'h0 : T204;
  assign T204 = T206 ? T205 : R203;
  assign T205 = R203 + 58'h1;
  assign T206 = T202 & T207;
  assign T207 = T201[3'h6:3'h6];
  assign T208 = T10[6'h29:6'h29];
  assign T209 = T223 | T210;
  assign T210 = T222 ? T211 : 64'h0;
  assign T211 = {R217, R212};
  assign T522 = reset ? 6'h0 : T213;
  assign T213 = T216 ? T214 : R212;
  assign T214 = T215[3'h5:1'h0];
  assign T215 = T523 + 7'h1;
  assign T523 = {1'h0, R212};
  assign T216 = io_uarch_counters_10 != 1'h0;
  assign T524 = reset ? 58'h0 : T218;
  assign T218 = T220 ? T219 : R217;
  assign T219 = R217 + 58'h1;
  assign T220 = T216 & T221;
  assign T221 = T215[3'h6:3'h6];
  assign T222 = T10[6'h28:6'h28];
  assign T223 = T237 | T224;
  assign T224 = T236 ? T225 : 64'h0;
  assign T225 = {R231, R226};
  assign T525 = reset ? 6'h0 : T227;
  assign T227 = T230 ? T228 : R226;
  assign T228 = T229[3'h5:1'h0];
  assign T229 = T526 + 7'h1;
  assign T526 = {1'h0, R226};
  assign T230 = io_uarch_counters_9 != 1'h0;
  assign T527 = reset ? 58'h0 : T232;
  assign T232 = T234 ? T233 : R231;
  assign T233 = R231 + 58'h1;
  assign T234 = T230 & T235;
  assign T235 = T229[3'h6:3'h6];
  assign T236 = T10[6'h27:6'h27];
  assign T237 = T251 | T238;
  assign T238 = T250 ? T239 : 64'h0;
  assign T239 = {R245, R240};
  assign T528 = reset ? 6'h0 : T241;
  assign T241 = T244 ? T242 : R240;
  assign T242 = T243[3'h5:1'h0];
  assign T243 = T529 + 7'h1;
  assign T529 = {1'h0, R240};
  assign T244 = io_uarch_counters_8 != 1'h0;
  assign T530 = reset ? 58'h0 : T246;
  assign T246 = T248 ? T247 : R245;
  assign T247 = R245 + 58'h1;
  assign T248 = T244 & T249;
  assign T249 = T243[3'h6:3'h6];
  assign T250 = T10[6'h26:6'h26];
  assign T251 = T265 | T252;
  assign T252 = T264 ? T253 : 64'h0;
  assign T253 = {R259, R254};
  assign T531 = reset ? 6'h0 : T255;
  assign T255 = T258 ? T256 : R254;
  assign T256 = T257[3'h5:1'h0];
  assign T257 = T532 + 7'h1;
  assign T532 = {1'h0, R254};
  assign T258 = io_uarch_counters_7 != 1'h0;
  assign T533 = reset ? 58'h0 : T260;
  assign T260 = T262 ? T261 : R259;
  assign T261 = R259 + 58'h1;
  assign T262 = T258 & T263;
  assign T263 = T257[3'h6:3'h6];
  assign T264 = T10[6'h25:6'h25];
  assign T265 = T279 | T266;
  assign T266 = T278 ? T267 : 64'h0;
  assign T267 = {R273, R268};
  assign T534 = reset ? 6'h0 : T269;
  assign T269 = T272 ? T270 : R268;
  assign T270 = T271[3'h5:1'h0];
  assign T271 = T535 + 7'h1;
  assign T535 = {1'h0, R268};
  assign T272 = io_uarch_counters_6 != 1'h0;
  assign T536 = reset ? 58'h0 : T274;
  assign T274 = T276 ? T275 : R273;
  assign T275 = R273 + 58'h1;
  assign T276 = T272 & T277;
  assign T277 = T271[3'h6:3'h6];
  assign T278 = T10[6'h24:6'h24];
  assign T279 = T293 | T280;
  assign T280 = T292 ? T281 : 64'h0;
  assign T281 = {R287, R282};
  assign T537 = reset ? 6'h0 : T283;
  assign T283 = T286 ? T284 : R282;
  assign T284 = T285[3'h5:1'h0];
  assign T285 = T538 + 7'h1;
  assign T538 = {1'h0, R282};
  assign T286 = io_uarch_counters_5 != 1'h0;
  assign T539 = reset ? 58'h0 : T288;
  assign T288 = T290 ? T289 : R287;
  assign T289 = R287 + 58'h1;
  assign T290 = T286 & T291;
  assign T291 = T285[3'h6:3'h6];
  assign T292 = T10[6'h23:6'h23];
  assign T293 = T307 | T294;
  assign T294 = T306 ? T295 : 64'h0;
  assign T295 = {R301, R296};
  assign T540 = reset ? 6'h0 : T297;
  assign T297 = T300 ? T298 : R296;
  assign T298 = T299[3'h5:1'h0];
  assign T299 = T541 + 7'h1;
  assign T541 = {1'h0, R296};
  assign T300 = io_uarch_counters_4 != 1'h0;
  assign T542 = reset ? 58'h0 : T302;
  assign T302 = T304 ? T303 : R301;
  assign T303 = R301 + 58'h1;
  assign T304 = T300 & T305;
  assign T305 = T299[3'h6:3'h6];
  assign T306 = T10[6'h22:6'h22];
  assign T307 = T321 | T308;
  assign T308 = T320 ? T309 : 64'h0;
  assign T309 = {R315, R310};
  assign T543 = reset ? 6'h0 : T311;
  assign T311 = T314 ? T312 : R310;
  assign T312 = T313[3'h5:1'h0];
  assign T313 = T544 + 7'h1;
  assign T544 = {1'h0, R310};
  assign T314 = io_uarch_counters_3 != 1'h0;
  assign T545 = reset ? 58'h0 : T316;
  assign T316 = T318 ? T317 : R315;
  assign T317 = R315 + 58'h1;
  assign T318 = T314 & T319;
  assign T319 = T313[3'h6:3'h6];
  assign T320 = T10[6'h21:6'h21];
  assign T321 = T335 | T322;
  assign T322 = T334 ? T323 : 64'h0;
  assign T323 = {R329, R324};
  assign T546 = reset ? 6'h0 : T325;
  assign T325 = T328 ? T326 : R324;
  assign T326 = T327[3'h5:1'h0];
  assign T327 = T547 + 7'h1;
  assign T547 = {1'h0, R324};
  assign T328 = io_uarch_counters_2 != 1'h0;
  assign T548 = reset ? 58'h0 : T330;
  assign T330 = T332 ? T331 : R329;
  assign T331 = R329 + 58'h1;
  assign T332 = T328 & T333;
  assign T333 = T327[3'h6:3'h6];
  assign T334 = T10[6'h20:6'h20];
  assign T335 = T349 | T336;
  assign T336 = T348 ? T337 : 64'h0;
  assign T337 = {R343, R338};
  assign T549 = reset ? 6'h0 : T339;
  assign T339 = T342 ? T340 : R338;
  assign T340 = T341[3'h5:1'h0];
  assign T341 = T550 + 7'h1;
  assign T550 = {1'h0, R338};
  assign T342 = io_uarch_counters_1 != 1'h0;
  assign T551 = reset ? 58'h0 : T344;
  assign T344 = T346 ? T345 : R343;
  assign T345 = R343 + 58'h1;
  assign T346 = T342 & T347;
  assign T347 = T341[3'h6:3'h6];
  assign T348 = T10[5'h1f:5'h1f];
  assign T349 = T363 | T350;
  assign T350 = T362 ? T351 : 64'h0;
  assign T351 = {R357, R352};
  assign T552 = reset ? 6'h0 : T353;
  assign T353 = T356 ? T354 : R352;
  assign T354 = T355[3'h5:1'h0];
  assign T355 = T553 + 7'h1;
  assign T553 = {1'h0, R352};
  assign T356 = io_uarch_counters_0 != 1'h0;
  assign T554 = reset ? 58'h0 : T358;
  assign T358 = T360 ? T359 : R357;
  assign T359 = R357 + 58'h1;
  assign T360 = T356 & T361;
  assign T361 = T355[3'h6:3'h6];
  assign T362 = T10[5'h1e:5'h1e];
  assign T363 = T365 | T364;
  assign T364 = T137 ? reg_cfgd : 64'h0;
  assign T365 = T367 | T366;
  assign T366 = T133 ? reg_cfga : 64'h0;
  assign T367 = T369 | T368;
  assign T368 = T120 ? reg_fromhost : 64'h0;
  assign T369 = T381 | T370;
  assign T370 = T380 ? reg_tohost : 64'h0;
  assign T555 = reset ? 64'h0 : T371;
  assign T371 = T376 ? wdata : T372;
  assign T372 = T373 ? 64'h0 : reg_tohost;
  assign T373 = T374 & T380;
  assign T374 = host_pcr_req_fire & T375;
  assign T375 = host_pcr_bits_rw ^ 1'h1;
  assign T376 = T379 & T377;
  assign T377 = T378 | host_pcr_req_fire;
  assign T378 = reg_tohost == 64'h0;
  assign T379 = wen & T380;
  assign T380 = T10[5'h15:5'h15];
  assign T381 = T387 | T556;
  assign T556 = {63'h0, T382};
  assign T382 = T386 ? reg_stats : 1'h0;
  assign T557 = reset ? 1'h0 : T383;
  assign T383 = T385 ? T384 : reg_stats;
  assign T384 = wdata[1'h0:1'h0];
  assign T385 = wen & T386;
  assign T386 = T10[2'h3:2'h3];
  assign T387 = T389 | T558;
  assign T558 = {62'h0, T388};
  assign T388 = T111 ? 2'h2 : 2'h0;
  assign T389 = T392 | T559;
  assign T559 = {62'h0, T390};
  assign T390 = T391 ? 2'h2 : 2'h0;
  assign T391 = T10[5'h12:5'h12];
  assign T392 = T394 | T560;
  assign T560 = {62'h0, T393};
  assign T393 = T37 ? 2'h2 : 2'h0;
  assign T394 = T397 | T561;
  assign T561 = {62'h0, T395};
  assign T395 = T396 ? 2'h2 : 2'h0;
  assign T396 = T10[5'h10:5'h10];
  assign T397 = T400 | T562;
  assign T562 = {63'h0, T398};
  assign T398 = T399 ? io_host_id : 1'h0;
  assign T399 = T10[4'hf:4'hf];
  assign T400 = T414 | T563;
  assign T563 = {32'h0, T401};
  assign T401 = T69 ? T402 : 32'h0;
  assign T402 = T403;
  assign T403 = {T409, T404};
  assign T404 = {T407, T405};
  assign T405 = {io_status_ei, T406};
  assign T406 = {io_status_ps, io_status_s};
  assign T407 = {io_status_u64, T408};
  assign T408 = {io_status_ef, io_status_pei};
  assign T409 = {T412, T410};
  assign T410 = {io_status_er, T411};
  assign T411 = {io_status_vm, io_status_s64};
  assign T412 = {io_status_ip, T413};
  assign T413 = {io_status_im, io_status_zero};
  assign T414 = T418 | T415;
  assign T415 = T417 ? reg_cause : 64'h0;
  assign T416 = io_exception ? io_cause : reg_cause;
  assign T417 = T10[4'hd:4'hd];
  assign T418 = T420 | T564;
  assign T564 = {21'h0, T419};
  assign T419 = T52 ? reg_evec : 43'h0;
  assign T420 = T422 | T565;
  assign T565 = {32'h0, T421};
  assign T421 = T129 ? reg_compare : 32'h0;
  assign T422 = T424 | T423;
  assign T423 = T27 ? T19 : 64'h0;
  assign T424 = T425 | 64'h0;
  assign T425 = T428 | T566;
  assign T566 = {32'h0, T426};
  assign T426 = T58 ? read_ptbr : 32'h0;
  assign read_ptbr = T427 << 4'hd;
  assign T427 = reg_ptbr[5'h1f:4'hd];
  assign T428 = T441 | T567;
  assign T567 = {21'h0, T429};
  assign T429 = T440 ? reg_badvaddr : 43'h0;
  assign T568 = T430[6'h2a:1'h0];
  assign T430 = io_badvaddr_wen ? T431 : T569;
  assign T569 = {1'h0, reg_badvaddr};
  assign T431 = T432;
  assign T432 = {T434, T433};
  assign T433 = io_rw_wdata[6'h2a:1'h0];
  assign T434 = T438 ? T437 : T435;
  assign T435 = T436 != 21'h0;
  assign T436 = io_rw_wdata[6'h3f:6'h2b];
  assign T437 = T436 == 21'h1fffff;
  assign T438 = $signed(T439) < $signed(1'h0);
  assign T439 = T433;
  assign T440 = T10[3'h7:3'h7];
  assign T441 = T443 | T570;
  assign T570 = {20'h0, T442};
  assign T442 = T46 ? reg_epc : 44'h0;
  assign T443 = T448 | T444;
  assign T444 = T447 ? reg_sup1 : 64'h0;
  assign T445 = T446 ? wdata : reg_sup1;
  assign T446 = wen & T447;
  assign T447 = T10[3'h5:3'h5];
  assign T448 = T453 | T449;
  assign T449 = T452 ? reg_sup0 : 64'h0;
  assign T450 = T451 ? wdata : reg_sup0;
  assign T451 = wen & T452;
  assign T452 = T10[3'h4:3'h4];
  assign T453 = T467 | T454;
  assign T454 = T466 ? T455 : 64'h0;
  assign T455 = {R461, R456};
  assign T571 = reset ? 6'h0 : T457;
  assign T457 = T460 ? T458 : R456;
  assign T458 = T459[3'h5:1'h0];
  assign T459 = T572 + 7'h1;
  assign T572 = {1'h0, R456};
  assign T460 = io_retire != 1'h0;
  assign T573 = reset ? 58'h0 : T462;
  assign T462 = T464 ? T463 : R461;
  assign T463 = R461 + 58'h1;
  assign T464 = T460 & T465;
  assign T465 = T459[3'h6:3'h6];
  assign T466 = T10[5'h1d:5'h1d];
  assign T467 = T470 | T468;
  assign T468 = T469 ? T19 : 64'h0;
  assign T469 = T10[5'h1c:5'h1c];
  assign T470 = T574 | T471;
  assign T471 = T472 ? T19 : 64'h0;
  assign T472 = T10[5'h1b:5'h1b];
  assign T574 = {56'h0, T473};
  assign T473 = T577 | T474;
  assign T474 = T18 ? T475 : 8'h0;
  assign T475 = {reg_frm, reg_fflags};
  assign T575 = T476[3'h4:1'h0];
  assign T476 = T17 ? wdata : T477;
  assign T477 = T480 ? wdata : T576;
  assign T576 = {59'h0, T478};
  assign T478 = io_fcsr_flags_valid ? T479 : reg_fflags;
  assign T479 = reg_fflags | io_fcsr_flags_bits;
  assign T480 = wen & T481;
  assign T481 = T10[1'h0:1'h0];
  assign T577 = {3'h0, T482};
  assign T482 = T484 | T578;
  assign T578 = {2'h0, T483};
  assign T483 = T9 ? reg_frm : 3'h0;
  assign T484 = T481 ? reg_fflags : 5'h0;
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T579;
  assign T579 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T485;
  assign T485 = cpu_req_valid & T391;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T486 = T488 ? 1'h0 : T487;
  assign T487 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T488 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T489;
  assign T489 = T491 & T490;
  assign T490 = host_pcr_rep_valid ^ 1'h1;
  assign T491 = host_pcr_req_valid ^ 1'h1;
  ManagementMachine temac_manage(.clk(clk), .reset(reset),
       //.io_stall_out(  )
       .io_write_to_cfga( T132 ),
       .io_cfgd_in( reg_cfgd ),
       .io_s_axi_awvalid( temac_manage_io_s_axi_awvalid ),
       .io_s_axi_awready( io_temac_s_axi_awready ),
       .io_s_axi_wvalid( temac_manage_io_s_axi_wvalid ),
       .io_s_axi_wready( io_temac_s_axi_wready ),
       .io_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_s_axi_bready( temac_manage_io_s_axi_bready ),
       .io_s_axi_arvalid( temac_manage_io_s_axi_arvalid ),
       //.io_s_axi_arready(  )
       .io_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_s_axi_rready( temac_manage_io_s_axi_rready )
  );

  always @(posedge clk) begin
    if(reset) begin
      reg_cfgd <= 64'h0;
    end else if(T136) begin
      reg_cfgd <= wdata;
    end
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T4) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T4) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(T4) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T4) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    reg_frm <= T492;
    if(reset) begin
      R20 <= 6'h0;
    end else if(T26) begin
      R20 <= T24;
    end else begin
      R20 <= T22;
    end
    if(reset) begin
      R28 <= 58'h0;
    end else if(T26) begin
      R28 <= T33;
    end else if(T32) begin
      R28 <= T31;
    end
    if(T45) begin
      reg_epc <= T43;
    end else if(io_exception) begin
      reg_epc <= T42;
    end
    if(T51) begin
      reg_evec <= T49;
    end
    if(T57) begin
      reg_ptbr <= T54;
    end
    if(reset) begin
      reg_status_s <= 1'h1;
    end else if(T68) begin
      reg_status_s <= T67;
    end else if(io_sret) begin
      reg_status_s <= reg_status_ps;
    end else if(io_exception) begin
      reg_status_s <= 1'h1;
    end
    if(reset) begin
      reg_status_ps <= 1'h0;
    end else if(T68) begin
      reg_status_ps <= T66;
    end else if(io_exception) begin
      reg_status_ps <= reg_status_s;
    end
    if(reset) begin
      reg_status_ei <= 1'h0;
    end else if(T68) begin
      reg_status_ei <= T78;
    end else if(io_sret) begin
      reg_status_ei <= reg_status_pei;
    end else if(io_exception) begin
      reg_status_ei <= 1'h0;
    end
    if(reset) begin
      reg_status_pei <= 1'h0;
    end else if(T68) begin
      reg_status_pei <= T77;
    end else if(io_exception) begin
      reg_status_pei <= reg_status_ei;
    end
    if(reset) begin
      reg_status_ef <= 1'h0;
    end else if(T68) begin
      reg_status_ef <= T81;
    end
    if(reset) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= T85;
    end
    if(reset) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= T89;
    end
    if(reset) begin
      reg_status_vm <= 1'h0;
    end else if(T68) begin
      reg_status_vm <= T92;
    end
    if(reset) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= T96;
    end
    if(reset) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= T100;
    end
    if(reset) begin
      reg_status_im <= 8'h0;
    end else if(T68) begin
      reg_status_im <= T103;
    end
    if(reset) begin
      r_irq_ipi <= 1'h1;
    end else if(io_host_ipi_rep_valid) begin
      r_irq_ipi <= 1'h1;
    end else if(T110) begin
      r_irq_ipi <= T109;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T115) begin
      reg_fromhost <= wdata;
    end
    if(reset) begin
      r_irq_timer <= 1'h0;
    end else if(T128) begin
      r_irq_timer <= 1'h0;
    end else if(T123) begin
      r_irq_timer <= 1'h1;
    end
    if(T128) begin
      reg_compare <= T125;
    end
    if(reset) begin
      reg_cfga <= 64'h0;
    end else if(T132) begin
      reg_cfga <= wdata;
    end
    if(reset) begin
      R142 <= 6'h0;
    end else if(T146) begin
      R142 <= T144;
    end
    if(reset) begin
      R147 <= 58'h0;
    end else if(T150) begin
      R147 <= T149;
    end
    if(reset) begin
      R156 <= 6'h0;
    end else if(T160) begin
      R156 <= T158;
    end
    if(reset) begin
      R161 <= 58'h0;
    end else if(T164) begin
      R161 <= T163;
    end
    if(reset) begin
      R170 <= 6'h0;
    end else if(T174) begin
      R170 <= T172;
    end
    if(reset) begin
      R175 <= 58'h0;
    end else if(T178) begin
      R175 <= T177;
    end
    if(reset) begin
      R184 <= 6'h0;
    end else if(T188) begin
      R184 <= T186;
    end
    if(reset) begin
      R189 <= 58'h0;
    end else if(T192) begin
      R189 <= T191;
    end
    if(reset) begin
      R198 <= 6'h0;
    end else if(T202) begin
      R198 <= T200;
    end
    if(reset) begin
      R203 <= 58'h0;
    end else if(T206) begin
      R203 <= T205;
    end
    if(reset) begin
      R212 <= 6'h0;
    end else if(T216) begin
      R212 <= T214;
    end
    if(reset) begin
      R217 <= 58'h0;
    end else if(T220) begin
      R217 <= T219;
    end
    if(reset) begin
      R226 <= 6'h0;
    end else if(T230) begin
      R226 <= T228;
    end
    if(reset) begin
      R231 <= 58'h0;
    end else if(T234) begin
      R231 <= T233;
    end
    if(reset) begin
      R240 <= 6'h0;
    end else if(T244) begin
      R240 <= T242;
    end
    if(reset) begin
      R245 <= 58'h0;
    end else if(T248) begin
      R245 <= T247;
    end
    if(reset) begin
      R254 <= 6'h0;
    end else if(T258) begin
      R254 <= T256;
    end
    if(reset) begin
      R259 <= 58'h0;
    end else if(T262) begin
      R259 <= T261;
    end
    if(reset) begin
      R268 <= 6'h0;
    end else if(T272) begin
      R268 <= T270;
    end
    if(reset) begin
      R273 <= 58'h0;
    end else if(T276) begin
      R273 <= T275;
    end
    if(reset) begin
      R282 <= 6'h0;
    end else if(T286) begin
      R282 <= T284;
    end
    if(reset) begin
      R287 <= 58'h0;
    end else if(T290) begin
      R287 <= T289;
    end
    if(reset) begin
      R296 <= 6'h0;
    end else if(T300) begin
      R296 <= T298;
    end
    if(reset) begin
      R301 <= 58'h0;
    end else if(T304) begin
      R301 <= T303;
    end
    if(reset) begin
      R310 <= 6'h0;
    end else if(T314) begin
      R310 <= T312;
    end
    if(reset) begin
      R315 <= 58'h0;
    end else if(T318) begin
      R315 <= T317;
    end
    if(reset) begin
      R324 <= 6'h0;
    end else if(T328) begin
      R324 <= T326;
    end
    if(reset) begin
      R329 <= 58'h0;
    end else if(T332) begin
      R329 <= T331;
    end
    if(reset) begin
      R338 <= 6'h0;
    end else if(T342) begin
      R338 <= T340;
    end
    if(reset) begin
      R343 <= 58'h0;
    end else if(T346) begin
      R343 <= T345;
    end
    if(reset) begin
      R352 <= 6'h0;
    end else if(T356) begin
      R352 <= T354;
    end
    if(reset) begin
      R357 <= 58'h0;
    end else if(T360) begin
      R357 <= T359;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T376) begin
      reg_tohost <= wdata;
    end else if(T373) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T385) begin
      reg_stats <= T384;
    end
    if(io_exception) begin
      reg_cause <= io_cause;
    end
    reg_badvaddr <= T568;
    if(T446) begin
      reg_sup1 <= wdata;
    end
    if(T451) begin
      reg_sup0 <= wdata;
    end
    if(reset) begin
      R456 <= 6'h0;
    end else if(T460) begin
      R456 <= T458;
    end
    if(reset) begin
      R461 <= 58'h0;
    end else if(T464) begin
      R461 <= T463;
    end
    reg_fflags <= T575;
    if(T488) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module Datapath(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [2:0] io_ctrl_sel_pc,
    input  io_ctrl_killd,
    input  io_ctrl_ren_1,
    input  io_ctrl_ren_0,
    input [2:0] io_ctrl_sel_alu2,
    input [1:0] io_ctrl_sel_alu1,
    input [2:0] io_ctrl_sel_imm,
    input  io_ctrl_fn_dw,
    input [3:0] io_ctrl_fn_alu,
    input  io_ctrl_div_mul_val,
    input  io_ctrl_div_mul_kill,
    //input  io_ctrl_div_val
    //input  io_ctrl_div_kill
    input [2:0] io_ctrl_csr,
    input  io_ctrl_sret,
    input  io_ctrl_mem_load,
    input  io_ctrl_wb_load,
    input  io_ctrl_ex_fp_val,
    input  io_ctrl_mem_fp_val,
    input  io_ctrl_ex_wen,
    input  io_ctrl_ex_valid,
    input  io_ctrl_mem_jalr,
    input  io_ctrl_mem_branch,
    input  io_ctrl_mem_wen,
    input  io_ctrl_wb_wen,
    input [2:0] io_ctrl_ex_mem_type,
    input  io_ctrl_ex_rs2_val,
    input  io_ctrl_ex_rocc_val,
    input  io_ctrl_mem_rocc_val,
    input  io_ctrl_bypass_1,
    input  io_ctrl_bypass_0,
    input [1:0] io_ctrl_bypass_src_1,
    input [1:0] io_ctrl_bypass_src_0,
    input  io_ctrl_ll_ready,
    input  io_ctrl_retire,
    input  io_ctrl_exception,
    input [63:0] io_ctrl_cause,
    input  io_ctrl_badvaddr_wen,
    output[31:0] io_ctrl_inst,
    //output io_ctrl_jalr_eq
    output io_ctrl_mem_br_taken,
    output io_ctrl_mem_misprediction,
    output io_ctrl_div_mul_rdy,
    output io_ctrl_ll_wen,
    output[4:0] io_ctrl_ll_waddr,
    output[4:0] io_ctrl_ex_waddr,
    output io_ctrl_mem_rs1_ra,
    output[4:0] io_ctrl_mem_waddr,
    output[4:0] io_ctrl_wb_waddr,
    output[7:0] io_ctrl_status_ip,
    output[7:0] io_ctrl_status_im,
    output[6:0] io_ctrl_status_zero,
    output io_ctrl_status_er,
    output io_ctrl_status_vm,
    output io_ctrl_status_s64,
    output io_ctrl_status_u64,
    output io_ctrl_status_ef,
    output io_ctrl_status_pei,
    output io_ctrl_status_ei,
    output io_ctrl_status_ps,
    output io_ctrl_status_s,
    output io_ctrl_fp_sboard_clr,
    output[4:0] io_ctrl_fp_sboard_clra,
    output io_ctrl_csr_replay,
    input  io_dmem_req_ready,
    //output io_dmem_req_valid
    //output io_dmem_req_bits_kill
    //output[2:0] io_dmem_req_bits_typ
    //output io_dmem_req_bits_phys
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    //output[4:0] io_dmem_req_bits_cmd
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    //output io_imem_req_valid
    output[43:0] io_imem_req_bits_pc,
    //output io_imem_resp_ready
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    //output io_imem_btb_update_valid
    //output io_imem_btb_update_bits_prediction_valid
    //output io_imem_btb_update_bits_prediction_bits_taken
    //output[42:0] io_imem_btb_update_bits_prediction_bits_target
    //output[5:0] io_imem_btb_update_bits_prediction_bits_entry
    //output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history
    //output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    //output io_imem_btb_update_bits_taken
    //output io_imem_btb_update_bits_isJump
    //output io_imem_btb_update_bits_isCall
    //output io_imem_btb_update_bits_isReturn
    //output io_imem_btb_update_bits_mispredict
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    //output io_imem_invalidate
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  reg  ex_reg_kill;
  wire T7;
  reg  mem_reg_kill;
  wire[31:0] T8;
  wire[63:0] T9;
  reg [63:0] R10;
  reg [63:0] R11;
  wire[63:0] ex_rs_1;
  wire[63:0] T12;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[63:0] id_rs_1;
  wire[63:0] T16;
  wire[63:0] T17;
  reg [63:0] T18 [30:0];
  wire[63:0] T19;
  wire T20;
  wire T21;
  wire[4:0] T22;
  wire T23;
  wire T24;
  wire[4:0] wb_waddr;
  wire wb_wen;
  wire[4:0] T25;
  wire[4:0] T26;
  wire[4:0] T27;
  wire[63:0] wb_wdata;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  reg [63:0] wb_reg_wdata;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] mem_int_wdata;
  reg [63:0] mem_reg_wdata;
  wire[63:0] T33;
  wire[63:0] T200;
  wire[44:0] mem_br_target;
  wire[44:0] T34;
  wire[44:0] T35;
  reg [43:0] mem_reg_pc;
  wire[43:0] T36;
  reg [43:0] ex_reg_pc;
  wire[43:0] T37;
  wire[44:0] T201;
  wire[21:0] T38;
  wire[21:0] T39;
  wire[21:0] T40;
  wire[21:0] T41;
  wire[11:0] T42;
  wire[4:0] T43;
  wire[3:0] T44;
  wire[6:0] T45;
  wire[5:0] T46;
  wire T47;
  wire T48;
  wire[9:0] T49;
  wire[8:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[21:0] T202;
  wire[14:0] T58;
  wire[14:0] T59;
  wire[11:0] T60;
  wire[4:0] T61;
  wire[3:0] T62;
  wire[6:0] T63;
  wire[5:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire[6:0] T203;
  wire T204;
  wire T71;
  wire[22:0] T205;
  wire T206;
  wire[18:0] T207;
  wire T208;
  wire T72;
  wire T73;
  wire[63:0] ll_wdata;
  wire T74;
  wire dmem_resp_xpu;
  wire T75;
  wire T76;
  wire dmem_resp_valid;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T81;
  wire[61:0] T82;
  wire T83;
  wire T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] T209;
  wire bypass_0;
  wire[63:0] bypass_1;
  wire T87;
  wire[1:0] T88;
  wire[63:0] T89;
  wire[63:0] bypass_2;
  wire[63:0] bypass_3;
  wire T90;
  wire T91;
  reg  ex_reg_rs_bypass_1;
  wire T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire[63:0] T95;
  reg [63:0] R96;
  reg [63:0] R97;
  wire[63:0] ex_rs_0;
  wire[63:0] T98;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire[63:0] id_rs_0;
  wire[63:0] T102;
  wire[63:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T110;
  wire[61:0] T111;
  wire T112;
  wire T113;
  wire[63:0] T114;
  wire[63:0] T115;
  wire[63:0] T210;
  wire T116;
  wire[1:0] T117;
  wire[63:0] T118;
  wire T119;
  wire T120;
  reg  ex_reg_rs_bypass_0;
  wire T121;
  wire[4:0] T122;
  wire[4:0] T123;
  wire T124;
  wire[63:0] T125;
  wire[4:0] T126;
  wire[4:0] T127;
  wire[43:0] T128;
  reg [43:0] wb_reg_pc;
  wire[43:0] T129;
  wire T130;
  wire[32:0] T131;
  wire[32:0] T132;
  wire T133;
  wire[1135:0] T134;
  wire[63:0] T223;
  wire[63:0] T224;
  wire[63:0] T225;
  wire[63:0] T226;
  wire T227;
  wire[63:0] T228;
  wire T229;
  wire[1:0] T230;
  wire[11:0] T231;
  wire T232;
  wire T193;
  wire dmem_resp_replay;
  reg  ex_reg_ctrl_fn_dw;
  wire T233;
  wire T234;
  reg [3:0] ex_reg_ctrl_fn_alu;
  wire[3:0] T235;
  wire[63:0] ex_op1;
  wire[63:0] T236;
  wire[43:0] T237;
  wire[43:0] T238;
  wire T239;
  reg [1:0] ex_reg_sel_alu1;
  wire[1:0] T240;
  wire[19:0] T241;
  wire T242;
  wire[63:0] T243;
  wire T244;
  wire[63:0] T245;
  wire[63:0] ex_op2;
  wire[63:0] T246;
  wire[31:0] T247;
  wire[31:0] T248;
  wire[3:0] T249;
  wire T250;
  reg [2:0] ex_reg_sel_alu2;
  wire[2:0] T251;
  wire[27:0] T252;
  wire T253;
  wire[31:0] ex_imm;
  wire[31:0] T254;
  wire[11:0] T255;
  wire[4:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  reg [2:0] ex_reg_sel_imm;
  wire[2:0] T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[3:0] T270;
  wire[3:0] T271;
  wire T272;
  wire[3:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[6:0] T278;
  wire[5:0] T279;
  wire[5:0] T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[19:0] T298;
  wire[18:0] T299;
  wire[7:0] T300;
  wire[7:0] T301;
  wire[7:0] T302;
  wire[7:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[10:0] T307;
  wire[10:0] T308;
  wire[10:0] T309;
  wire[10:0] T310;
  wire T311;
  wire T312;
  wire[31:0] T313;
  wire T314;
  wire[63:0] T315;
  wire T316;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T135;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T136;
  wire[6:0] T137;
  wire[4:0] T138;
  wire T139;
  wire T140;
  wire T141;
  wire[4:0] T142;
  wire[4:0] T143;
  wire[6:0] T144;
  wire[4:0] T211;
  wire[6:0] dmem_resp_waddr;
  wire[7:0] T145;
  wire T146;
  wire dmem_resp_fpu;
  wire T147;
  wire[42:0] T212;
  wire[42:0] T213;
  wire[42:0] T214;
  wire[43:0] T215;
  wire[44:0] T148;
  wire[44:0] T149;
  wire[44:0] T216;
  wire[43:0] T150;
  wire T151;
  wire[44:0] mem_npc;
  wire[44:0] T217;
  wire[43:0] T152;
  wire[42:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[1:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[21:0] T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire[7:0] T218;
  wire[5:0] T168;
  wire[63:0] T169;
  wire[43:0] T170;
  wire[43:0] T171;
  wire[42:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire[1:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire[21:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[4:0] T219;
  wire T186;
  wire[4:0] T187;
  wire[4:0] T188;
  wire T189;
  wire[4:0] T190;
  wire[4:0] T191;
  wire[4:0] T220;
  wire[6:0] T192;
  wire[6:0] T221;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire[44:0] T222;
  wire T199;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;
  wire pcr_io_host_pcr_req_ready;
  wire pcr_io_host_pcr_rep_valid;
  wire[63:0] pcr_io_host_pcr_rep_bits;
  wire pcr_io_host_ipi_req_valid;
  wire pcr_io_host_ipi_req_bits;
  wire pcr_io_host_ipi_rep_ready;
  wire pcr_io_host_debug_stats_pcr;
  wire[63:0] pcr_io_rw_rdata;
  wire pcr_io_temac_rx_axis_fifo_tready;
  wire[7:0] pcr_io_temac_tx_axis_fifo_tdata;
  wire pcr_io_temac_tx_axis_fifo_tvalid;
  wire pcr_io_temac_tx_axis_fifo_tlast;
  wire[11:0] pcr_io_temac_s_axi_awaddr;
  wire pcr_io_temac_s_axi_awvalid;
  wire[31:0] pcr_io_temac_s_axi_wdata;
  wire pcr_io_temac_s_axi_wvalid;
  wire pcr_io_temac_s_axi_bready;
  wire[11:0] pcr_io_temac_s_axi_araddr;
  wire pcr_io_temac_s_axi_arvalid;
  wire pcr_io_temac_s_axi_rready;
  wire[7:0] pcr_io_status_ip;
  wire[7:0] pcr_io_status_im;
  wire[6:0] pcr_io_status_zero;
  wire pcr_io_status_er;
  wire pcr_io_status_vm;
  wire pcr_io_status_s64;
  wire pcr_io_status_u64;
  wire pcr_io_status_ef;
  wire pcr_io_status_pei;
  wire pcr_io_status_ei;
  wire pcr_io_status_ps;
  wire pcr_io_status_s;
  wire[31:0] pcr_io_ptbr;
  wire[43:0] pcr_io_evec;
  wire pcr_io_fatc;
  wire pcr_io_replay;
  wire[63:0] pcr_io_time;
  wire[2:0] pcr_io_fcsr_rm;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_kill = {1{$random}};
    mem_reg_kill = {1{$random}};
    R10 = {2{$random}};
    R11 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T18[initvar] = {2{$random}};
    wb_reg_wdata = {2{$random}};
    mem_reg_wdata = {2{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R96 = {2{$random}};
    R97 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    ex_reg_ctrl_fn_dw = {1{$random}};
    ex_reg_ctrl_fn_alu = {1{$random}};
    ex_reg_sel_alu1 = {1{$random}};
    ex_reg_sel_alu2 = {1{$random}};
    ex_reg_sel_imm = {1{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
  end
`endif

  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T7 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T6 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data : ex_reg_inst;
  assign T5 = io_ctrl_killd ^ 1'h1;
  assign T6 = ex_reg_kill ^ 1'h1;
  assign T7 = mem_reg_kill ^ 1'h1;
  assign T8 = wb_reg_inst;
  assign T9 = R10;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T85 : T12;
  assign T12 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T13 = T80 ? io_ctrl_bypass_src_1 : T14;
  assign T14 = T79 ? T15 : ex_reg_rs_lsb_1;
  assign T15 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T16;
  assign T16 = T77 ? wb_wdata : T17;
  assign T17 = T18[T26];
  assign T20 = T23 & T21;
  assign T21 = T22 < 5'h1f;
  assign T22 = T25[3'h4:1'h0];
  assign T23 = wb_wen & T24;
  assign T24 = wb_waddr != 5'h0;
  assign wb_waddr = io_ctrl_ll_wen ? io_ctrl_ll_waddr : io_ctrl_wb_waddr;
  assign wb_wen = io_ctrl_ll_wen | io_ctrl_wb_wen;
  assign T25 = ~ wb_waddr;
  assign T26 = ~ T27;
  assign T27 = io_imem_resp_bits_data[5'h18:5'h14];
  assign wb_wdata = T28;
  assign T28 = T74 ? io_dmem_resp_bits_data_subword : T29;
  assign T29 = io_ctrl_ll_wen ? ll_wdata : T30;
  assign T30 = T73 ? pcr_io_rw_rdata : wb_reg_wdata;
  assign T31 = T7 ? T32 : wb_reg_wdata;
  assign T32 = T72 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = io_ctrl_mem_jalr ? T200 : mem_reg_wdata;
  assign T33 = T6 ? alu_io_out : mem_reg_wdata;
  assign T200 = {T207, mem_br_target};
  assign mem_br_target = T201 + T34;
  assign T34 = T35;
  assign T35 = {1'h0, mem_reg_pc};
  assign T36 = T6 ? ex_reg_pc : mem_reg_pc;
  assign T37 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T201 = {T205, T38};
  assign T38 = T71 ? T202 : T39;
  assign T39 = T55 ? T40 : 22'h4;
  assign T40 = T41;
  assign T41 = {T49, T42};
  assign T42 = {T45, T43};
  assign T43 = {T44, 1'h0};
  assign T44 = mem_reg_inst[5'h18:5'h15];
  assign T45 = {T47, T46};
  assign T46 = mem_reg_inst[5'h1e:5'h19];
  assign T47 = T48;
  assign T48 = mem_reg_inst[5'h14:5'h14];
  assign T49 = {T53, T50};
  assign T50 = {T53, T51};
  assign T51 = T52;
  assign T52 = mem_reg_inst[5'h13:4'hc];
  assign T53 = T54;
  assign T54 = mem_reg_inst[5'h1f:5'h1f];
  assign T55 = T57 & T56;
  assign T56 = io_ctrl_mem_branch ^ 1'h1;
  assign T57 = io_ctrl_mem_jalr ^ 1'h1;
  assign T202 = {T203, T58};
  assign T58 = T59;
  assign T59 = {T67, T60};
  assign T60 = {T63, T61};
  assign T61 = {T62, 1'h0};
  assign T62 = mem_reg_inst[4'hb:4'h8];
  assign T63 = {T65, T64};
  assign T64 = mem_reg_inst[5'h1e:5'h19];
  assign T65 = T66;
  assign T66 = mem_reg_inst[3'h7:3'h7];
  assign T67 = {T69, T68};
  assign T68 = {T69, T69};
  assign T69 = T70;
  assign T70 = mem_reg_inst[5'h1f:5'h1f];
  assign T203 = T204 ? 7'h7f : 7'h0;
  assign T204 = T58[4'he:4'he];
  assign T71 = io_ctrl_mem_branch & io_ctrl_mem_br_taken;
  assign T205 = T206 ? 23'h7fffff : 23'h0;
  assign T206 = T38[5'h15:5'h15];
  assign T207 = T208 ? 19'h7ffff : 19'h0;
  assign T208 = mem_br_target[6'h2c:6'h2c];
  assign T72 = io_ctrl_mem_fp_val & io_ctrl_mem_wen;
  assign T73 = io_ctrl_csr != 3'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign T74 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_xpu = T75 ^ 1'h1;
  assign T75 = T76;
  assign T76 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T77 = T23 & T78;
  assign T78 = wb_waddr == T27;
  assign T79 = T5 & io_ctrl_ren_1;
  assign T80 = T5 & io_ctrl_bypass_1;
  assign T81 = T83 ? T82 : ex_reg_rs_msb_1;
  assign T82 = id_rs_1 >> 2'h2;
  assign T83 = T79 & T84;
  assign T84 = io_ctrl_bypass_1 ^ 1'h1;
  assign T85 = T91 ? T89 : T86;
  assign T86 = T87 ? bypass_1 : T209;
  assign T209 = {63'h0, bypass_0};
  assign bypass_0 = 1'h0;
  assign bypass_1 = mem_reg_wdata;
  assign T87 = T88[1'h0:1'h0];
  assign T88 = ex_reg_rs_lsb_1;
  assign T89 = T90 ? bypass_3 : bypass_2;
  assign bypass_2 = wb_reg_wdata;
  assign bypass_3 = io_dmem_resp_bits_data;
  assign T90 = T88[1'h0:1'h0];
  assign T91 = T88[1'h1:1'h1];
  assign T92 = T5 ? io_ctrl_bypass_1 : ex_reg_rs_bypass_1;
  assign T93 = T94;
  assign T94 = wb_reg_inst[5'h18:5'h14];
  assign T95 = R96;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T114 : T98;
  assign T98 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T99 = T109 ? io_ctrl_bypass_src_0 : T100;
  assign T100 = T108 ? T101 : ex_reg_rs_lsb_0;
  assign T101 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T102;
  assign T102 = T106 ? wb_wdata : T103;
  assign T103 = T18[T104];
  assign T104 = ~ T105;
  assign T105 = io_imem_resp_bits_data[5'h13:4'hf];
  assign T106 = T23 & T107;
  assign T107 = wb_waddr == T105;
  assign T108 = T5 & io_ctrl_ren_0;
  assign T109 = T5 & io_ctrl_bypass_0;
  assign T110 = T112 ? T111 : ex_reg_rs_msb_0;
  assign T111 = id_rs_0 >> 2'h2;
  assign T112 = T108 & T113;
  assign T113 = io_ctrl_bypass_0 ^ 1'h1;
  assign T114 = T120 ? T118 : T115;
  assign T115 = T116 ? bypass_1 : T210;
  assign T210 = {63'h0, bypass_0};
  assign T116 = T117[1'h0:1'h0];
  assign T117 = ex_reg_rs_lsb_0;
  assign T118 = T119 ? bypass_3 : bypass_2;
  assign T119 = T117[1'h0:1'h0];
  assign T120 = T117[1'h1:1'h1];
  assign T121 = T5 ? io_ctrl_bypass_0 : ex_reg_rs_bypass_0;
  assign T122 = T123;
  assign T123 = wb_reg_inst[5'h13:4'hf];
  assign T124 = wb_wen;
  assign T125 = wb_wdata;
  assign T126 = T127;
  assign T127 = wb_wen ? wb_waddr : 5'h0;
  assign T128 = wb_reg_pc;
  assign T129 = T7 ? mem_reg_pc : wb_reg_pc;
  assign T130 = io_ctrl_retire;
  assign T131 = T132;
  assign T132 = pcr_io_time[6'h20:1'h0];
  assign T133 = io_host_id;
  assign T223 = T229 ? T228 : T224;
  assign T224 = T227 ? T225 : wb_reg_wdata;
  assign T225 = pcr_io_rw_rdata & T226;
  assign T226 = ~ wb_reg_wdata;
  assign T227 = io_ctrl_csr == 3'h3;
  assign T228 = pcr_io_rw_rdata | wb_reg_wdata;
  assign T229 = io_ctrl_csr == 3'h2;
  assign T230 = io_ctrl_csr[1'h1:1'h0];
  assign T231 = wb_reg_inst[5'h1f:5'h14];
  assign T232 = T193 ? 1'h0 : io_ctrl_ll_ready;
  assign T193 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T233 = T5 ? T234 : ex_reg_ctrl_fn_dw;
  assign T234 = io_ctrl_fn_dw;
  assign T235 = T5 ? io_ctrl_fn_alu : ex_reg_ctrl_fn_alu;
  assign ex_op1 = T244 ? T243 : T236;
  assign T236 = {T241, T237};
  assign T237 = T239 ? T238 : 44'h0;
  assign T238 = ex_reg_pc;
  assign T239 = ex_reg_sel_alu1 == 2'h2;
  assign T240 = T5 ? io_ctrl_sel_alu1 : ex_reg_sel_alu1;
  assign T241 = T242 ? 20'hfffff : 20'h0;
  assign T242 = T237[6'h2b:6'h2b];
  assign T243 = ex_rs_0;
  assign T244 = ex_reg_sel_alu1 == 2'h1;
  assign T245 = ex_op2;
  assign ex_op2 = T316 ? T315 : T246;
  assign T246 = {T313, T247};
  assign T247 = T312 ? ex_imm : T248;
  assign T248 = {T252, T249};
  assign T249 = T250 ? 4'h4 : 4'h0;
  assign T250 = ex_reg_sel_alu2 == 3'h1;
  assign T251 = T5 ? io_ctrl_sel_alu2 : ex_reg_sel_alu2;
  assign T252 = T253 ? 28'hfffffff : 28'h0;
  assign T253 = T249[2'h3:2'h3];
  assign ex_imm = T254;
  assign T254 = {T298, T255};
  assign T255 = {T278, T256};
  assign T256 = {T267, T257};
  assign T257 = T266 ? T265 : T258;
  assign T258 = T264 ? T263 : T259;
  assign T259 = T261 ? T260 : 1'h0;
  assign T260 = ex_reg_inst[4'hf:4'hf];
  assign T261 = ex_reg_sel_imm == 3'h5;
  assign T262 = T5 ? io_ctrl_sel_imm : ex_reg_sel_imm;
  assign T263 = ex_reg_inst[5'h14:5'h14];
  assign T264 = ex_reg_sel_imm == 3'h4;
  assign T265 = ex_reg_inst[3'h7:3'h7];
  assign T266 = ex_reg_sel_imm == 3'h0;
  assign T267 = T277 ? 4'h0 : T268;
  assign T268 = T274 ? T273 : T269;
  assign T269 = T272 ? T271 : T270;
  assign T270 = ex_reg_inst[5'h18:5'h15];
  assign T271 = ex_reg_inst[5'h13:5'h10];
  assign T272 = ex_reg_sel_imm == 3'h5;
  assign T273 = ex_reg_inst[4'hb:4'h8];
  assign T274 = T276 | T275;
  assign T275 = ex_reg_sel_imm == 3'h1;
  assign T276 = ex_reg_sel_imm == 3'h0;
  assign T277 = ex_reg_sel_imm == 3'h2;
  assign T278 = {T284, T279};
  assign T279 = T281 ? 6'h0 : T280;
  assign T280 = ex_reg_inst[5'h1e:5'h19];
  assign T281 = T283 | T282;
  assign T282 = ex_reg_sel_imm == 3'h5;
  assign T283 = ex_reg_sel_imm == 3'h2;
  assign T284 = T295 ? 1'h0 : T285;
  assign T285 = T294 ? T292 : T286;
  assign T286 = T291 ? T289 : T287;
  assign T287 = T288;
  assign T288 = ex_reg_inst[5'h1f:5'h1f];
  assign T289 = T290;
  assign T290 = ex_reg_inst[3'h7:3'h7];
  assign T291 = ex_reg_sel_imm == 3'h1;
  assign T292 = T293;
  assign T293 = ex_reg_inst[5'h14:5'h14];
  assign T294 = ex_reg_sel_imm == 3'h3;
  assign T295 = T297 | T296;
  assign T296 = ex_reg_sel_imm == 3'h5;
  assign T297 = ex_reg_sel_imm == 3'h2;
  assign T298 = {T287, T299};
  assign T299 = {T307, T300};
  assign T300 = T304 ? T303 : T301;
  assign T301 = T302;
  assign T302 = ex_reg_inst[5'h13:4'hc];
  assign T303 = T287 ? 8'hff : 8'h0;
  assign T304 = T306 & T305;
  assign T305 = ex_reg_sel_imm != 3'h3;
  assign T306 = ex_reg_sel_imm != 3'h2;
  assign T307 = T311 ? T309 : T308;
  assign T308 = T287 ? 11'h7ff : 11'h0;
  assign T309 = T310;
  assign T310 = ex_reg_inst[5'h1e:5'h14];
  assign T311 = ex_reg_sel_imm == 3'h2;
  assign T312 = ex_reg_sel_alu2 == 3'h3;
  assign T313 = T314 ? 32'hffffffff : 32'h0;
  assign T314 = T247[5'h1f:5'h1f];
  assign T315 = ex_rs_1;
  assign T316 = ex_reg_sel_alu2 == 3'h2;
  assign io_temac_s_axi_rready = pcr_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = pcr_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = pcr_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = pcr_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = pcr_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = pcr_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = pcr_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = pcr_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = pcr_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = pcr_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = pcr_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = pcr_io_temac_rx_axis_fifo_tready;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T135 = io_ctrl_mem_rocc_val ? mem_reg_rs2 : wb_reg_rs2;
  assign T136 = io_ctrl_ex_rs2_val ? ex_rs_1 : mem_reg_rs2;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_inst_opcode = T137;
  assign T137 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T138;
  assign T138 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T139;
  assign T139 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T140;
  assign T140 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T141;
  assign T141 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T142;
  assign T142 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T143;
  assign T143 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T144;
  assign T144 = wb_reg_inst[5'h1f:5'h19];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = T211;
  assign T211 = dmem_resp_waddr[3'h4:1'h0];
  assign dmem_resp_waddr = T145 >> 1'h1;
  assign T145 = io_dmem_resp_bits_tag;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T146;
  assign T146 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T147;
  assign T147 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = pcr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data;
  assign io_imem_btb_update_bits_returnAddr = T212;
  assign T212 = mem_int_wdata[6'h2a:1'h0];
  assign io_imem_btb_update_bits_target = T213;
  assign T213 = io_imem_req_bits_pc[6'h2a:1'h0];
  assign io_imem_btb_update_bits_pc = T214;
  assign T214 = mem_reg_pc[6'h2a:1'h0];
  assign io_imem_req_bits_pc = T215;
  assign T215 = T148[6'h2b:1'h0];
  assign T148 = T149;
  assign T149 = T167 ? mem_npc : T216;
  assign T216 = {1'h0, T150};
  assign T150 = T151 ? pcr_io_evec : wb_reg_pc;
  assign T151 = io_ctrl_sel_pc == 3'h3;
  assign mem_npc = io_ctrl_mem_jalr ? T217 : mem_br_target;
  assign T217 = {1'h0, T152};
  assign T152 = {T154, T153};
  assign T153 = mem_reg_wdata[6'h2a:1'h0];
  assign T154 = T164 ? T163 : T155;
  assign T155 = T159 ? T158 : T156;
  assign T156 = T157[1'h0:1'h0];
  assign T157 = mem_reg_wdata[6'h2b:6'h2a];
  assign T158 = T157 == 2'h3;
  assign T159 = T162 | T160;
  assign T160 = T161 == 22'h3ffffe;
  assign T161 = mem_reg_wdata >> 6'h2a;
  assign T162 = T161 == 22'h3fffff;
  assign T163 = T157 != 2'h0;
  assign T164 = T166 | T165;
  assign T165 = T161 == 22'h1;
  assign T166 = T161 == 22'h0;
  assign T167 = io_ctrl_sel_pc == 3'h1;
  assign io_ptw_status_s = pcr_io_status_s;
  assign io_ptw_status_ps = pcr_io_status_ps;
  assign io_ptw_status_ei = pcr_io_status_ei;
  assign io_ptw_status_pei = pcr_io_status_pei;
  assign io_ptw_status_ef = pcr_io_status_ef;
  assign io_ptw_status_u64 = pcr_io_status_u64;
  assign io_ptw_status_s64 = pcr_io_status_s64;
  assign io_ptw_status_vm = pcr_io_status_vm;
  assign io_ptw_status_er = pcr_io_status_er;
  assign io_ptw_status_zero = pcr_io_status_zero;
  assign io_ptw_status_im = pcr_io_status_im;
  assign io_ptw_status_ip = pcr_io_status_ip;
  assign io_ptw_sret = io_ctrl_sret;
  assign io_ptw_invalidate = pcr_io_fatc;
  assign io_ptw_ptbr = pcr_io_ptbr;
  assign io_dmem_req_bits_tag = T218;
  assign T218 = {2'h0, T168};
  assign T168 = {io_ctrl_ex_waddr, io_ctrl_ex_fp_val};
  assign io_dmem_req_bits_data = T169;
  assign T169 = io_ctrl_mem_fp_val ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_addr = T170;
  assign T170 = T171;
  assign T171 = {T173, T172};
  assign T172 = alu_io_adder_out[6'h2a:1'h0];
  assign T173 = T183 ? T182 : T174;
  assign T174 = T178 ? T177 : T175;
  assign T175 = T176[1'h0:1'h0];
  assign T176 = alu_io_adder_out[6'h2b:6'h2a];
  assign T177 = T176 == 2'h3;
  assign T178 = T181 | T179;
  assign T179 = T180 == 22'h3ffffe;
  assign T180 = ex_rs_0 >> 6'h2a;
  assign T181 = T180 == 22'h3fffff;
  assign T182 = T176 != 2'h0;
  assign T183 = T185 | T184;
  assign T184 = T180 == 22'h1;
  assign T185 = T180 == 22'h0;
  assign io_ctrl_csr_replay = pcr_io_replay;
  assign io_ctrl_fp_sboard_clra = T219;
  assign T219 = dmem_resp_waddr[3'h4:1'h0];
  assign io_ctrl_fp_sboard_clr = T186;
  assign T186 = dmem_resp_replay & dmem_resp_fpu;
  assign io_ctrl_status_s = pcr_io_status_s;
  assign io_ctrl_status_ps = pcr_io_status_ps;
  assign io_ctrl_status_ei = pcr_io_status_ei;
  assign io_ctrl_status_pei = pcr_io_status_pei;
  assign io_ctrl_status_ef = pcr_io_status_ef;
  assign io_ctrl_status_u64 = pcr_io_status_u64;
  assign io_ctrl_status_s64 = pcr_io_status_s64;
  assign io_ctrl_status_vm = pcr_io_status_vm;
  assign io_ctrl_status_er = pcr_io_status_er;
  assign io_ctrl_status_zero = pcr_io_status_zero;
  assign io_ctrl_status_im = pcr_io_status_im;
  assign io_ctrl_status_ip = pcr_io_status_ip;
  assign io_ctrl_wb_waddr = T187;
  assign T187 = wb_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_waddr = T188;
  assign T188 = mem_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_rs1_ra = T189;
  assign T189 = T190 == 5'h1;
  assign T190 = mem_reg_inst[5'h13:4'hf];
  assign io_ctrl_ex_waddr = T191;
  assign T191 = ex_reg_inst[4'hb:3'h7];
  assign io_ctrl_ll_waddr = T220;
  assign T220 = T192[3'h4:1'h0];
  assign T192 = T193 ? dmem_resp_waddr : T221;
  assign T221 = {2'h0, div_io_resp_bits_tag};
  assign io_ctrl_ll_wen = T194;
  assign T194 = T193 ? 1'h1 : T195;
  assign T195 = T232 & div_io_resp_valid;
  assign io_ctrl_div_mul_rdy = div_io_req_ready;
  assign io_ctrl_mem_misprediction = T196;
  assign T196 = T198 | T197;
  assign T197 = io_ctrl_ex_valid ^ 1'h1;
  assign T198 = mem_npc != T222;
  assign T222 = {1'h0, ex_reg_pc};
  assign io_ctrl_mem_br_taken = T199;
  assign T199 = mem_reg_wdata[1'h0:1'h0];
  assign io_ctrl_inst = io_imem_resp_bits_data;
  assign io_host_debug_stats_pcr = pcr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = pcr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = pcr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = pcr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = pcr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = pcr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = pcr_io_host_pcr_req_ready;
  ALU alu(
       .io_dw( ex_reg_ctrl_fn_dw ),
       .io_fn( ex_reg_ctrl_fn_alu ),
       .io_in2( T245 ),
       .io_in1( ex_op1 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( io_ctrl_div_mul_val ),
       .io_req_bits_fn( ex_reg_ctrl_fn_alu ),
       .io_req_bits_dw( ex_reg_ctrl_fn_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( io_ctrl_ex_waddr ),
       .io_kill( io_ctrl_div_mul_kill ),
       .io_resp_ready( T232 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );
  CSRFile pcr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( pcr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( pcr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( pcr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( pcr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( pcr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( pcr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( pcr_io_host_debug_stats_pcr ),
       .io_rw_addr( T231 ),
       .io_rw_cmd( T230 ),
       .io_rw_rdata( pcr_io_rw_rdata ),
       .io_rw_wdata( T223 ),
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( pcr_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( pcr_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( pcr_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( pcr_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( pcr_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( pcr_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( pcr_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( pcr_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( pcr_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( pcr_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( pcr_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( pcr_io_temac_s_axi_rready ),
       .io_status_ip( pcr_io_status_ip ),
       .io_status_im( pcr_io_status_im ),
       .io_status_zero( pcr_io_status_zero ),
       .io_status_er( pcr_io_status_er ),
       .io_status_vm( pcr_io_status_vm ),
       .io_status_s64( pcr_io_status_s64 ),
       .io_status_u64( pcr_io_status_u64 ),
       .io_status_ef( pcr_io_status_ef ),
       .io_status_pei( pcr_io_status_pei ),
       .io_status_ei( pcr_io_status_ei ),
       .io_status_ps( pcr_io_status_ps ),
       .io_status_s( pcr_io_status_s ),
       .io_ptbr( pcr_io_ptbr ),
       .io_evec( pcr_io_evec ),
       .io_exception( io_ctrl_exception ),
       .io_retire( io_ctrl_retire ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( io_ctrl_cause ),
       .io_badvaddr_wen( io_ctrl_badvaddr_wen ),
       .io_pc( wb_reg_pc ),
       .io_sret( io_ctrl_sret ),
       .io_fatc( pcr_io_fatc ),
       .io_replay( pcr_io_replay ),
       .io_time( pcr_io_time ),
       .io_fcsr_rm( pcr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );

  always @(posedge clk) begin
    if(T7) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T6) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data;
    end
    ex_reg_kill <= io_ctrl_killd;
    mem_reg_kill <= ex_reg_kill;
    R10 <= R11;
    if(ex_reg_rs_bypass_1) begin
      R11 <= T85;
    end else begin
      R11 <= T12;
    end
    if(T80) begin
      ex_reg_rs_lsb_1 <= io_ctrl_bypass_src_1;
    end else if(T79) begin
      ex_reg_rs_lsb_1 <= T15;
    end
    if (T20)
      T18[T25] <= wb_wdata;
    if(T7) begin
      wb_reg_wdata <= T32;
    end
    if(T6) begin
      mem_reg_wdata <= alu_io_out;
    end
    if(T6) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T83) begin
      ex_reg_rs_msb_1 <= T82;
    end
    if(T5) begin
      ex_reg_rs_bypass_1 <= io_ctrl_bypass_1;
    end
    R96 <= R97;
    if(ex_reg_rs_bypass_0) begin
      R97 <= T114;
    end else begin
      R97 <= T98;
    end
    if(T109) begin
      ex_reg_rs_lsb_0 <= io_ctrl_bypass_src_0;
    end else if(T108) begin
      ex_reg_rs_lsb_0 <= T101;
    end
    if(T112) begin
      ex_reg_rs_msb_0 <= T111;
    end
    if(T5) begin
      ex_reg_rs_bypass_0 <= io_ctrl_bypass_0;
    end
    if(T7) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if(T5) begin
      ex_reg_ctrl_fn_dw <= T234;
    end
    if(T5) begin
      ex_reg_ctrl_fn_alu <= io_ctrl_fn_alu;
    end
    if(T5) begin
      ex_reg_sel_alu1 <= io_ctrl_sel_alu1;
    end
    if(T5) begin
      ex_reg_sel_alu2 <= io_ctrl_sel_alu2;
    end
    if(T5) begin
      ex_reg_sel_imm <= io_ctrl_sel_imm;
    end
    if(io_ctrl_mem_rocc_val) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(io_ctrl_ex_rs2_val) begin
      mem_reg_rs2 <= ex_rs_1;
    end
`ifndef SYNTHESIS
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T133, T131, T130, T128, T126, T125, T124, T122, T95, T93, T9, T8, T1);
`endif
  end
endmodule

module FPUDecoder(
    input [31:0] io_inst,
    output[4:0] io_sigs_cmd,
    output io_sigs_ldst,
    output io_sigs_wen,
    output io_sigs_ren1,
    output io_sigs_ren2,
    output io_sigs_ren3,
    output io_sigs_swap23,
    output io_sigs_single,
    output io_sigs_fromint,
    output io_sigs_toint,
    output io_sigs_fastpipe,
    output io_sigs_fma,
    output io_sigs_round
);

  wire T0;
  wire T1;
  wire[31:0] T2;
  wire T3;
  wire T4;
  wire[31:0] T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  wire T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire T16;
  wire[31:0] T17;
  wire T18;
  wire T19;
  wire[31:0] T20;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire[31:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire T41;
  wire[31:0] T42;
  wire T43;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire[31:0] T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire[31:0] T55;
  wire T56;
  wire T57;
  wire[31:0] T58;
  wire T59;
  wire T60;
  wire[31:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[31:0] T65;
  wire T66;
  wire T67;
  wire[31:0] T68;
  wire T69;
  wire T70;
  wire[31:0] T71;
  wire T72;
  wire T73;
  wire[31:0] T74;
  wire T75;
  wire T76;
  wire[31:0] T77;
  wire T78;
  wire T79;
  wire[31:0] T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[31:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire[31:0] T114;
  wire[4:0] T115;
  wire[3:0] T116;
  wire[2:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire[31:0] T121;
  wire T122;
  wire[31:0] T123;
  wire T124;
  wire T125;
  wire[31:0] T126;
  wire T127;
  wire[31:0] T128;
  wire T129;
  wire T130;
  wire[31:0] T131;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire T135;
  wire[31:0] T136;
  wire T137;
  wire[31:0] T138;


  assign io_sigs_round = T0;
  assign T0 = T3 | T1;
  assign T1 = T2 == 32'he0000053;
  assign T2 = io_inst & 32'hedf0707f;
  assign T3 = T6 | T4;
  assign T4 = T5 == 32'he0000053;
  assign T5 = io_inst & 32'hfdf0607f;
  assign T6 = T9 | T7;
  assign T7 = T8 == 32'hc0000053;
  assign T8 = io_inst & 32'hedc0007f;
  assign T9 = T12 | T10;
  assign T10 = T11 == 32'h42000053;
  assign T11 = io_inst & 32'h7ff0007f;
  assign T12 = T15 | T13;
  assign T13 = T14 == 32'h40100053;
  assign T14 = io_inst & 32'h7ff0007f;
  assign T15 = T18 | T16;
  assign T16 = T17 == 32'h53;
  assign T17 = io_inst & 32'hec00007f;
  assign T18 = T21 | T19;
  assign T19 = T20 == 32'h53;
  assign T20 = io_inst & 32'hf400007f;
  assign T21 = T22 == 32'h43;
  assign T22 = io_inst & 32'h4000073;
  assign io_sigs_fma = T23;
  assign T23 = T24 | T16;
  assign T24 = T21 | T19;
  assign io_sigs_fastpipe = T25;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h42000053;
  assign T27 = io_inst & 32'hfff0007f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h40100053;
  assign T30 = io_inst & 32'hfff0007f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h20000053;
  assign T33 = io_inst & 32'hf400607f;
  assign T34 = T35 == 32'h20000053;
  assign T35 = io_inst & 32'hfc00507f;
  assign io_sigs_toint = T36;
  assign T36 = T37 | T4;
  assign T37 = T40 | T38;
  assign T38 = T39 == 32'hc0000053;
  assign T39 = io_inst & 32'hfdc0007f;
  assign T40 = T43 | T41;
  assign T41 = T42 == 32'ha0000053;
  assign T42 = io_inst & 32'hfc00507f;
  assign T43 = T46 | T44;
  assign T44 = T45 == 32'ha0000053;
  assign T45 = io_inst & 32'hfc00607f;
  assign T46 = T47 == 32'h2027;
  assign T47 = io_inst & 32'h607f;
  assign io_sigs_fromint = T48;
  assign T48 = T51 | T49;
  assign T49 = T50 == 32'hf0000053;
  assign T50 = io_inst & 32'hfdf0707f;
  assign T51 = T52 == 32'hd0000053;
  assign T52 = io_inst & 32'hfdc0007f;
  assign io_sigs_single = T53;
  assign T53 = T56 | T54;
  assign T54 = T55 == 32'he0000053;
  assign T55 = io_inst & 32'heff0707f;
  assign T56 = T59 | T57;
  assign T57 = T58 == 32'he0000053;
  assign T58 = io_inst & 32'hfff0607f;
  assign T59 = T62 | T60;
  assign T60 = T61 == 32'hc0000053;
  assign T61 = io_inst & 32'hefc0007f;
  assign T62 = T63 | T13;
  assign T63 = T66 | T64;
  assign T64 = T65 == 32'h20000053;
  assign T65 = io_inst & 32'h7e00507f;
  assign T66 = T69 | T67;
  assign T67 = T68 == 32'h20000053;
  assign T68 = io_inst & 32'h7e00607f;
  assign T69 = T72 | T70;
  assign T70 = T71 == 32'h20000053;
  assign T71 = io_inst & 32'hf600607f;
  assign T72 = T75 | T73;
  assign T73 = T74 == 32'h2007;
  assign T74 = io_inst & 32'h705f;
  assign T75 = T78 | T76;
  assign T76 = T77 == 32'h53;
  assign T77 = io_inst & 32'hee00007f;
  assign T78 = T81 | T79;
  assign T79 = T80 == 32'h53;
  assign T80 = io_inst & 32'hf600007f;
  assign T81 = T82 == 32'h43;
  assign T82 = io_inst & 32'h6000073;
  assign io_sigs_swap23 = T19;
  assign io_sigs_ren3 = T21;
  assign io_sigs_ren2 = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h20000053;
  assign T85 = io_inst & 32'h7c00507f;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h20000053;
  assign T88 = io_inst & 32'h7c00607f;
  assign T89 = T90 | T32;
  assign T90 = T91 | T46;
  assign T91 = T92 | T16;
  assign T92 = T21 | T19;
  assign io_sigs_ren1 = T93;
  assign T93 = T94 | T4;
  assign T94 = T95 | T38;
  assign T95 = T96 | T10;
  assign T96 = T97 | T13;
  assign T97 = T98 | T84;
  assign T98 = T99 | T87;
  assign T99 = T100 | T32;
  assign T100 = T101 | T16;
  assign T101 = T21 | T19;
  assign io_sigs_wen = T102;
  assign T102 = T103 | T49;
  assign T103 = T104 | T51;
  assign T104 = T105 | T26;
  assign T105 = T106 | T29;
  assign T106 = T107 | T32;
  assign T107 = T108 | T34;
  assign T108 = T111 | T109;
  assign T109 = T110 == 32'h2007;
  assign T110 = io_inst & 32'h607f;
  assign T111 = T112 | T16;
  assign T112 = T21 | T19;
  assign io_sigs_ldst = T113;
  assign T113 = T114 == 32'h2007;
  assign T114 = io_inst & 32'h605f;
  assign io_sigs_cmd = T115;
  assign T115 = {T137, T116};
  assign T116 = {T134, T117};
  assign T117 = {T129, T118};
  assign T118 = {T124, T119};
  assign T119 = T122 | T120;
  assign T120 = T121 == 32'h8000010;
  assign T121 = io_inst & 32'h8000010;
  assign T122 = T123 == 32'h4;
  assign T123 = io_inst & 32'h4;
  assign T124 = T127 | T125;
  assign T125 = T126 == 32'h10000010;
  assign T126 = io_inst & 32'h10000010;
  assign T127 = T128 == 32'h8;
  assign T128 = io_inst & 32'h8;
  assign T129 = T132 | T130;
  assign T130 = T131 == 32'h20000000;
  assign T131 = io_inst & 32'h20000000;
  assign T132 = T133 == 32'h0;
  assign T133 = io_inst & 32'h40;
  assign T134 = T132 | T135;
  assign T135 = T136 == 32'h40000000;
  assign T136 = io_inst & 32'h40000000;
  assign T137 = T138 == 32'h0;
  assign T138 = io_inst & 32'h10;
endmodule

module mulAddSubRecodedFloatN_0(
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[27:0] T4;
  wire[27:0] T529;
  wire[25:0] T5;
  wire[26:0] roundMask;
  wire[26:0] T6;
  wire[24:0] T7;
  wire[24:0] T530;
  wire T8;
  wire[24:0] T9;
  wire[8:0] T10;
  wire T11;
  wire[8:0] T12;
  wire[24:0] T13;
  wire[1024:0] T14;
  wire[9:0] T15;
  wire[9:0] sExpX3_13;
  wire[10:0] sExpX3;
  wire[10:0] T531;
  wire[6:0] estNormDist;
  wire[6:0] T16;
  wire[6:0] estNormNeg_dist;
  wire[6:0] T17;
  wire[6:0] T18;
  wire[6:0] T19;
  wire[6:0] T20;
  wire[6:0] T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[6:0] T24;
  wire[6:0] T25;
  wire[6:0] T26;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[6:0] T29;
  wire[6:0] T30;
  wire[6:0] T31;
  wire[6:0] T32;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[6:0] T40;
  wire[6:0] T41;
  wire[6:0] T42;
  wire[6:0] T43;
  wire[6:0] T44;
  wire[6:0] T45;
  wire[6:0] T46;
  wire[6:0] T47;
  wire[6:0] T48;
  wire[6:0] T49;
  wire[6:0] T50;
  wire[6:0] T51;
  wire[6:0] T52;
  wire[6:0] T53;
  wire[6:0] T54;
  wire[6:0] T55;
  wire[6:0] T56;
  wire[6:0] T57;
  wire[6:0] T58;
  wire[6:0] T59;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire T65;
  wire[50:0] T66;
  wire[50:0] T67;
  wire[49:0] T68;
  wire[49:0] T69;
  wire[74:0] sigSum;
  wire[74:0] alignedNegSigC;
  wire[75:0] T70;
  wire T71;
  wire doSubMags;
  wire opSignC;
  wire T72;
  wire T73;
  wire signProd;
  wire T74;
  wire T75;
  wire signB;
  wire signA;
  wire T76;
  wire[23:0] T77;
  wire[23:0] CExtraMask;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[6:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[5:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[3:0] T89;
  wire[7:0] T90;
  wire[23:0] T91;
  wire[128:0] T92;
  wire[6:0] CAlignDist;
  wire[10:0] T93;
  wire[10:0] T94;
  wire[10:0] sNatCAlignDist;
  wire[10:0] T532;
  wire[8:0] expC;
  wire[10:0] sExpAlignedProd;
  wire[10:0] T95;
  wire[10:0] T533;
  wire[8:0] expA;
  wire[10:0] T96;
  wire[7:0] T97;
  wire[8:0] expB;
  wire[2:0] T98;
  wire[2:0] T534;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire CAlignDist_floor;
  wire T103;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T104;
  wire isZeroA;
  wire[2:0] T105;
  wire[7:0] T106;
  wire[7:0] T535;
  wire[3:0] T107;
  wire[7:0] T108;
  wire[7:0] T536;
  wire[5:0] T109;
  wire[7:0] T110;
  wire[7:0] T537;
  wire[6:0] T111;
  wire[15:0] T112;
  wire[15:0] T113;
  wire[15:0] T114;
  wire[14:0] T115;
  wire[15:0] T116;
  wire[15:0] T117;
  wire[15:0] T118;
  wire[13:0] T119;
  wire[15:0] T120;
  wire[15:0] T121;
  wire[15:0] T122;
  wire[11:0] T123;
  wire[15:0] T124;
  wire[15:0] T125;
  wire[15:0] T126;
  wire[7:0] T127;
  wire[15:0] T128;
  wire[15:0] T129;
  wire[15:0] T538;
  wire[7:0] T130;
  wire[15:0] T131;
  wire[15:0] T539;
  wire[11:0] T132;
  wire[15:0] T133;
  wire[15:0] T540;
  wire[13:0] T134;
  wire[15:0] T135;
  wire[15:0] T541;
  wire[14:0] T136;
  wire[23:0] sigC;
  wire[22:0] fractC;
  wire T137;
  wire isZeroC;
  wire[2:0] T138;
  wire[74:0] T139;
  wire[74:0] T140;
  wire[74:0] T141;
  wire[73:0] T142;
  wire[49:0] T143;
  wire[49:0] T542;
  wire[23:0] negSigC;
  wire[23:0] T144;
  wire[74:0] T543;
  wire[48:0] T145;
  wire[47:0] T146;
  wire[23:0] sigB;
  wire[22:0] fractB;
  wire T147;
  wire[23:0] sigA;
  wire[22:0] fractA;
  wire T148;
  wire[50:0] T544;
  wire[49:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire notCDom_signSigSum;
  wire[6:0] CDom_estNormDist;
  wire[6:0] T545;
  wire[4:0] T198;
  wire[6:0] T199;
  wire T200;
  wire CAlignDist_0;
  wire T201;
  wire[9:0] T202;
  wire isCDominant;
  wire T203;
  wire T204;
  wire[9:0] T205;
  wire T206;
  wire[10:0] sExpSum;
  wire[10:0] T546;
  wire[7:0] T207;
  wire[7:0] T208;
  wire[7:0] T209;
  wire[6:0] T210;
  wire[7:0] T211;
  wire[7:0] T212;
  wire[7:0] T213;
  wire[5:0] T214;
  wire[7:0] T215;
  wire[7:0] T216;
  wire[7:0] T217;
  wire[3:0] T218;
  wire[7:0] T219;
  wire[7:0] T220;
  wire[7:0] T547;
  wire[3:0] T221;
  wire[7:0] T222;
  wire[7:0] T548;
  wire[5:0] T223;
  wire[7:0] T224;
  wire[7:0] T549;
  wire[6:0] T225;
  wire[15:0] T226;
  wire[15:0] T227;
  wire[15:0] T228;
  wire[14:0] T229;
  wire[15:0] T230;
  wire[15:0] T231;
  wire[15:0] T232;
  wire[13:0] T233;
  wire[15:0] T234;
  wire[15:0] T235;
  wire[15:0] T236;
  wire[11:0] T237;
  wire[15:0] T238;
  wire[15:0] T239;
  wire[15:0] T240;
  wire[7:0] T241;
  wire[15:0] T242;
  wire[15:0] T243;
  wire[15:0] T550;
  wire[7:0] T244;
  wire[15:0] T245;
  wire[15:0] T551;
  wire[11:0] T246;
  wire[15:0] T247;
  wire[15:0] T552;
  wire[13:0] T248;
  wire[15:0] T249;
  wire[15:0] T553;
  wire[14:0] T250;
  wire[26:0] T251;
  wire[26:0] T554;
  wire T252;
  wire[27:0] sigX3;
  wire[42:0] T253;
  wire T254;
  wire T255;
  wire[15:0] T256;
  wire[15:0] absSigSumExtraMask;
  wire[14:0] T257;
  wire[6:0] T258;
  wire[2:0] T259;
  wire T260;
  wire[2:0] T261;
  wire[6:0] T262;
  wire[14:0] T263;
  wire[16:0] T264;
  wire[3:0] normTo2ShiftDist;
  wire[3:0] estNormDist_5;
  wire[3:0] T265;
  wire[1:0] T266;
  wire T267;
  wire[1:0] T268;
  wire T269;
  wire[3:0] T270;
  wire[1:0] T271;
  wire T272;
  wire[1:0] T273;
  wire[3:0] T274;
  wire T275;
  wire[1:0] T276;
  wire T277;
  wire[1:0] T278;
  wire T279;
  wire[7:0] T280;
  wire[7:0] T281;
  wire[7:0] T282;
  wire[6:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[7:0] T286;
  wire[5:0] T287;
  wire[7:0] T288;
  wire[7:0] T289;
  wire[7:0] T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T293;
  wire[7:0] T555;
  wire[3:0] T294;
  wire[7:0] T295;
  wire[7:0] T556;
  wire[5:0] T296;
  wire[7:0] T297;
  wire[7:0] T557;
  wire[6:0] T298;
  wire[15:0] T299;
  wire[42:0] cFirstNormAbsSigSum;
  wire[42:0] T558;
  wire[41:0] T300;
  wire[41:0] notCDom_pos_firstNormAbsSigSum;
  wire[41:0] T301;
  wire[41:0] T302;
  wire[31:0] T303;
  wire[31:0] T559;
  wire[9:0] T304;
  wire[41:0] T560;
  wire[33:0] T305;
  wire T306;
  wire T307;
  wire[1:0] firstReduceSigSum;
  wire T308;
  wire[17:0] T309;
  wire T310;
  wire[15:0] T311;
  wire T312;
  wire T313;
  wire[1:0] firstReduceNotSigSum;
  wire T314;
  wire[17:0] T315;
  wire[74:0] notSigSum;
  wire T316;
  wire[15:0] T317;
  wire[32:0] T318;
  wire T319;
  wire[41:0] T320;
  wire[41:0] T321;
  wire[41:0] T322;
  wire[15:0] T323;
  wire[15:0] T561;
  wire[25:0] T324;
  wire T325;
  wire T326;
  wire[41:0] CDom_firstNormAbsSigSum;
  wire[41:0] T327;
  wire[41:0] T328;
  wire[41:0] T329;
  wire T330;
  wire[40:0] T331;
  wire[41:0] T562;
  wire T332;
  wire T333;
  wire T334;
  wire[41:0] T335;
  wire[41:0] T336;
  wire[41:0] T337;
  wire T338;
  wire[40:0] T339;
  wire[41:0] T563;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[41:0] T344;
  wire[41:0] T345;
  wire[41:0] T346;
  wire T347;
  wire[40:0] T348;
  wire[41:0] T564;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire[41:0] T353;
  wire[41:0] T354;
  wire T355;
  wire[40:0] T356;
  wire[41:0] T565;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire[42:0] T362;
  wire[42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[42:0] T363;
  wire[42:0] T364;
  wire[10:0] T365;
  wire[42:0] T566;
  wire[32:0] T366;
  wire T367;
  wire[31:0] T368;
  wire T369;
  wire[42:0] T370;
  wire[42:0] T567;
  wire[41:0] T371;
  wire[42:0] T372;
  wire[26:0] T373;
  wire T374;
  wire T375;
  wire[42:0] T568;
  wire T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[41:0] T380;
  wire[41:0] T381;
  wire roundPosBit;
  wire[27:0] T382;
  wire[27:0] T569;
  wire[26:0] roundPosMask;
  wire[26:0] T570;
  wire[25:0] T383;
  wire[25:0] T384;
  wire T385;
  wire allRound;
  wire allRoundExtra;
  wire[27:0] T386;
  wire[27:0] T571;
  wire[25:0] T387;
  wire[27:0] T388;
  wire doIncrSig;
  wire T389;
  wire T390;
  wire T391;
  wire commonCase;
  wire T392;
  wire notSpecial_addZeros;
  wire T393;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T394;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T395;
  wire isSpecialA;
  wire[1:0] T396;
  wire underflow;
  wire underflowY;
  wire T397;
  wire T398;
  wire[9:0] T572;
  wire[7:0] T399;
  wire sigX3Shift1;
  wire[1:0] T400;
  wire T401;
  wire overflow;
  wire overflowY;
  wire[2:0] T402;
  wire[10:0] sExpY;
  wire[10:0] T403;
  wire[10:0] T404;
  wire T405;
  wire[1:0] T406;
  wire[25:0] sigY3;
  wire[25:0] T407;
  wire[25:0] T408;
  wire[25:0] T409;
  wire[25:0] T410;
  wire[25:0] roundUp_sigY3;
  wire[25:0] T411;
  wire[25:0] T412;
  wire[27:0] T413;
  wire[27:0] T573;
  wire roundEven;
  wire T414;
  wire T415;
  wire T416;
  wire roundingMode_nearest_even;
  wire T417;
  wire T418;
  wire T419;
  wire[25:0] T420;
  wire[25:0] T421;
  wire roundUp;
  wire T422;
  wire T423;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T424;
  wire doNegSignSum;
  wire T425;
  wire T426;
  wire T427;
  wire isZeroY;
  wire[2:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire[25:0] T442;
  wire[25:0] T443;
  wire[27:0] T444;
  wire[27:0] T574;
  wire[26:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[10:0] T449;
  wire[10:0] T450;
  wire T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire[1:0] T455;
  wire invalid;
  wire notSigNaN_invalid;
  wire T456;
  wire T457;
  wire isInfC;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire isInfB;
  wire T462;
  wire T463;
  wire isInfA;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire isNaNB;
  wire T468;
  wire T469;
  wire isNaNA;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire isSigNaNC;
  wire T475;
  wire T476;
  wire isNaNC;
  wire T477;
  wire T478;
  wire isSigNaNB;
  wire T479;
  wire T480;
  wire isSigNaNA;
  wire T481;
  wire T482;
  wire[32:0] T483;
  wire[31:0] T484;
  wire[22:0] fractOut;
  wire[22:0] T485;
  wire[22:0] T575;
  wire T486;
  wire isSatOut;
  wire T487;
  wire overflowY_roundMagUp;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire isNaNOut;
  wire T492;
  wire T493;
  wire[22:0] fractY;
  wire[22:0] T494;
  wire[22:0] T495;
  wire[8:0] expOut;
  wire[8:0] T496;
  wire[8:0] T497;
  wire[8:0] T498;
  wire notNaN_isInfOut;
  wire T499;
  wire T500;
  wire T501;
  wire[8:0] T502;
  wire[8:0] T503;
  wire[8:0] T504;
  wire[8:0] T505;
  wire[8:0] T506;
  wire[8:0] T507;
  wire[8:0] T508;
  wire[8:0] T509;
  wire[8:0] T510;
  wire[8:0] T511;
  wire[8:0] T512;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T513;
  wire[8:0] T514;
  wire T515;
  wire T516;
  wire[8:0] expY;
  wire signOut;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;


  assign io_exceptionFlags = T0;
  assign T0 = {T455, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T385 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 28'h0;
  assign T4 = sigX3 & T529;
  assign T529 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T251 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T530;
  assign T530 = {24'h0, T8};
  assign T8 = sigX3[5'h1a:5'h1a];
  assign T9 = {T226, T10};
  assign T10 = {T207, T11};
  assign T11 = T12[4'h8:4'h8];
  assign T12 = T13[5'h18:5'h10];
  assign T13 = T14[8'h83:7'h6b];
  assign T14 = $signed(1025'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T15;
  assign T15 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'h9:1'h0];
  assign sExpX3 = sExpSum - T531;
  assign T531 = {4'h0, estNormDist};
  assign estNormDist = isCDominant ? CDom_estNormDist : T16;
  assign T16 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = T197 ? 7'h18 : T17;
  assign T17 = T196 ? 7'h19 : T18;
  assign T18 = T195 ? 7'h1a : T19;
  assign T19 = T194 ? 7'h1b : T20;
  assign T20 = T193 ? 7'h1c : T21;
  assign T21 = T192 ? 7'h1d : T22;
  assign T22 = T191 ? 7'h1e : T23;
  assign T23 = T190 ? 7'h1f : T24;
  assign T24 = T189 ? 7'h20 : T25;
  assign T25 = T188 ? 7'h21 : T26;
  assign T26 = T187 ? 7'h22 : T27;
  assign T27 = T186 ? 7'h23 : T28;
  assign T28 = T185 ? 7'h24 : T29;
  assign T29 = T184 ? 7'h25 : T30;
  assign T30 = T183 ? 7'h26 : T31;
  assign T31 = T182 ? 7'h27 : T32;
  assign T32 = T181 ? 7'h28 : T33;
  assign T33 = T180 ? 7'h29 : T34;
  assign T34 = T179 ? 7'h2a : T35;
  assign T35 = T178 ? 7'h2b : T36;
  assign T36 = T177 ? 7'h2c : T37;
  assign T37 = T176 ? 7'h2d : T38;
  assign T38 = T175 ? 7'h2e : T39;
  assign T39 = T174 ? 7'h2f : T40;
  assign T40 = T173 ? 7'h30 : T41;
  assign T41 = T172 ? 7'h31 : T42;
  assign T42 = T171 ? 7'h32 : T43;
  assign T43 = T170 ? 7'h33 : T44;
  assign T44 = T169 ? 7'h34 : T45;
  assign T45 = T168 ? 7'h35 : T46;
  assign T46 = T167 ? 7'h36 : T47;
  assign T47 = T166 ? 7'h37 : T48;
  assign T48 = T165 ? 7'h38 : T49;
  assign T49 = T164 ? 7'h39 : T50;
  assign T50 = T163 ? 7'h3a : T51;
  assign T51 = T162 ? 7'h3b : T52;
  assign T52 = T161 ? 7'h3c : T53;
  assign T53 = T160 ? 7'h3d : T54;
  assign T54 = T159 ? 7'h3e : T55;
  assign T55 = T158 ? 7'h3f : T56;
  assign T56 = T157 ? 7'h40 : T57;
  assign T57 = T156 ? 7'h41 : T58;
  assign T58 = T155 ? 7'h42 : T59;
  assign T59 = T154 ? 7'h43 : T60;
  assign T60 = T153 ? 7'h44 : T61;
  assign T61 = T152 ? 7'h45 : T62;
  assign T62 = T151 ? 7'h46 : T63;
  assign T63 = T150 ? 7'h47 : T64;
  assign T64 = T65 ? 7'h48 : 7'h49;
  assign T65 = T66[1'h1:1'h1];
  assign T66 = T544 ^ T67;
  assign T67 = T68 << 1'h1;
  assign T68 = 50'h0 | T69;
  assign T69 = sigSum[6'h32:1'h1];
  assign sigSum = T543 + alignedNegSigC;
  assign alignedNegSigC = T70[7'h4a:1'h0];
  assign T70 = {T139, T71};
  assign T71 = T76 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T73 ^ T72;
  assign T72 = io_op[1'h0:1'h0];
  assign T73 = io_c[6'h20:6'h20];
  assign signProd = T75 ^ T74;
  assign T74 = io_op[1'h1:1'h1];
  assign T75 = signA ^ signB;
  assign signB = io_b[6'h20:6'h20];
  assign signA = io_a[6'h20:6'h20];
  assign T76 = T77 != 24'h0;
  assign T77 = sigC & CExtraMask;
  assign CExtraMask = {T112, T78};
  assign T78 = T110 | T79;
  assign T79 = T80 & 8'haa;
  assign T80 = T81 << 1'h1;
  assign T81 = T82[3'h6:1'h0];
  assign T82 = T108 | T83;
  assign T83 = T84 & 8'hcc;
  assign T84 = T85 << 2'h2;
  assign T85 = T86[3'h5:1'h0];
  assign T86 = T106 | T87;
  assign T87 = T88 & 8'hf0;
  assign T88 = T89 << 3'h4;
  assign T89 = T90[2'h3:1'h0];
  assign T90 = T91[5'h17:5'h10];
  assign T91 = T92[7'h4d:6'h36];
  assign T92 = $signed(129'h100000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = T93[3'h6:1'h0];
  assign T93 = CAlignDist_floor ? 11'h0 : T94;
  assign T94 = T101 ? sNatCAlignDist : 11'h4a;
  assign sNatCAlignDist = sExpAlignedProd - T532;
  assign T532 = {2'h0, expC};
  assign expC = io_c[5'h1f:5'h17];
  assign sExpAlignedProd = T95 + 11'h1b;
  assign T95 = T96 + T533;
  assign T533 = {2'h0, expA};
  assign expA = io_a[5'h1f:5'h17];
  assign T96 = {T98, T97};
  assign T97 = expB[3'h7:1'h0];
  assign expB = io_b[5'h1f:5'h17];
  assign T98 = 3'h0 - T534;
  assign T534 = {2'h0, T99};
  assign T99 = T100 ^ 1'h1;
  assign T100 = expB[4'h8:4'h8];
  assign T101 = T102 < 10'h4a;
  assign T102 = sNatCAlignDist[4'h9:1'h0];
  assign CAlignDist_floor = isZeroProd | T103;
  assign T103 = sNatCAlignDist[4'ha:4'ha];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T104 == 3'h0;
  assign T104 = expB[4'h8:3'h6];
  assign isZeroA = T105 == 3'h0;
  assign T105 = expA[4'h8:3'h6];
  assign T106 = T535 & 8'hf;
  assign T535 = {4'h0, T107};
  assign T107 = T90 >> 3'h4;
  assign T108 = T536 & 8'h33;
  assign T536 = {2'h0, T109};
  assign T109 = T86 >> 2'h2;
  assign T110 = T537 & 8'h55;
  assign T537 = {1'h0, T111};
  assign T111 = T82 >> 1'h1;
  assign T112 = T135 | T113;
  assign T113 = T114 & 16'haaaa;
  assign T114 = T115 << 1'h1;
  assign T115 = T116[4'he:1'h0];
  assign T116 = T133 | T117;
  assign T117 = T118 & 16'hcccc;
  assign T118 = T119 << 2'h2;
  assign T119 = T120[4'hd:1'h0];
  assign T120 = T131 | T121;
  assign T121 = T122 & 16'hf0f0;
  assign T122 = T123 << 3'h4;
  assign T123 = T124[4'hb:1'h0];
  assign T124 = T129 | T125;
  assign T125 = T126 & 16'hff00;
  assign T126 = T127 << 4'h8;
  assign T127 = T128[3'h7:1'h0];
  assign T128 = T91[4'hf:1'h0];
  assign T129 = T538 & 16'hff;
  assign T538 = {8'h0, T130};
  assign T130 = T128 >> 4'h8;
  assign T131 = T539 & 16'hf0f;
  assign T539 = {4'h0, T132};
  assign T132 = T124 >> 3'h4;
  assign T133 = T540 & 16'h3333;
  assign T540 = {2'h0, T134};
  assign T134 = T120 >> 2'h2;
  assign T135 = T541 & 16'h5555;
  assign T541 = {1'h0, T136};
  assign T136 = T116 >> 1'h1;
  assign sigC = {T137, fractC};
  assign fractC = io_c[5'h16:1'h0];
  assign T137 = isZeroC ^ 1'h1;
  assign isZeroC = T138 == 3'h0;
  assign T138 = expC[4'h8:3'h6];
  assign T139 = $signed(T140) >>> CAlignDist;
  assign T140 = T141;
  assign T141 = {doSubMags, T142};
  assign T142 = {negSigC, T143};
  assign T143 = 50'h0 - T542;
  assign T542 = {49'h0, doSubMags};
  assign negSigC = doSubMags ? T144 : sigC;
  assign T144 = ~ sigC;
  assign T543 = {26'h0, T145};
  assign T145 = T146 << 1'h1;
  assign T146 = sigA * sigB;
  assign sigB = {T147, fractB};
  assign fractB = io_b[5'h16:1'h0];
  assign T147 = isZeroB ^ 1'h1;
  assign sigA = {T148, fractA};
  assign fractA = io_a[5'h16:1'h0];
  assign T148 = isZeroA ^ 1'h1;
  assign T544 = {1'h0, T149};
  assign T149 = 50'h0 ^ T69;
  assign T150 = T66[2'h2:2'h2];
  assign T151 = T66[2'h3:2'h3];
  assign T152 = T66[3'h4:3'h4];
  assign T153 = T66[3'h5:3'h5];
  assign T154 = T66[3'h6:3'h6];
  assign T155 = T66[3'h7:3'h7];
  assign T156 = T66[4'h8:4'h8];
  assign T157 = T66[4'h9:4'h9];
  assign T158 = T66[4'ha:4'ha];
  assign T159 = T66[4'hb:4'hb];
  assign T160 = T66[4'hc:4'hc];
  assign T161 = T66[4'hd:4'hd];
  assign T162 = T66[4'he:4'he];
  assign T163 = T66[4'hf:4'hf];
  assign T164 = T66[5'h10:5'h10];
  assign T165 = T66[5'h11:5'h11];
  assign T166 = T66[5'h12:5'h12];
  assign T167 = T66[5'h13:5'h13];
  assign T168 = T66[5'h14:5'h14];
  assign T169 = T66[5'h15:5'h15];
  assign T170 = T66[5'h16:5'h16];
  assign T171 = T66[5'h17:5'h17];
  assign T172 = T66[5'h18:5'h18];
  assign T173 = T66[5'h19:5'h19];
  assign T174 = T66[5'h1a:5'h1a];
  assign T175 = T66[5'h1b:5'h1b];
  assign T176 = T66[5'h1c:5'h1c];
  assign T177 = T66[5'h1d:5'h1d];
  assign T178 = T66[5'h1e:5'h1e];
  assign T179 = T66[5'h1f:5'h1f];
  assign T180 = T66[6'h20:6'h20];
  assign T181 = T66[6'h21:6'h21];
  assign T182 = T66[6'h22:6'h22];
  assign T183 = T66[6'h23:6'h23];
  assign T184 = T66[6'h24:6'h24];
  assign T185 = T66[6'h25:6'h25];
  assign T186 = T66[6'h26:6'h26];
  assign T187 = T66[6'h27:6'h27];
  assign T188 = T66[6'h28:6'h28];
  assign T189 = T66[6'h29:6'h29];
  assign T190 = T66[6'h2a:6'h2a];
  assign T191 = T66[6'h2b:6'h2b];
  assign T192 = T66[6'h2c:6'h2c];
  assign T193 = T66[6'h2d:6'h2d];
  assign T194 = T66[6'h2e:6'h2e];
  assign T195 = T66[6'h2f:6'h2f];
  assign T196 = T66[6'h30:6'h30];
  assign T197 = T66[6'h31:6'h31];
  assign notCDom_signSigSum = sigSum[6'h33:6'h33];
  assign CDom_estNormDist = T200 ? CAlignDist : T545;
  assign T545 = {2'h0, T198};
  assign T198 = T199[3'h4:1'h0];
  assign T199 = CAlignDist - 7'h1;
  assign T200 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T201;
  assign T201 = T202 == 10'h0;
  assign T202 = sNatCAlignDist[4'h9:1'h0];
  assign isCDominant = T206 & T203;
  assign T203 = CAlignDist_floor | T204;
  assign T204 = T205 < 10'h19;
  assign T205 = sNatCAlignDist[4'h9:1'h0];
  assign T206 = isZeroC ^ 1'h1;
  assign sExpSum = CAlignDist_floor ? T546 : sExpAlignedProd;
  assign T546 = {2'h0, expC};
  assign T207 = T224 | T208;
  assign T208 = T209 & 8'haa;
  assign T209 = T210 << 1'h1;
  assign T210 = T211[3'h6:1'h0];
  assign T211 = T222 | T212;
  assign T212 = T213 & 8'hcc;
  assign T213 = T214 << 2'h2;
  assign T214 = T215[3'h5:1'h0];
  assign T215 = T220 | T216;
  assign T216 = T217 & 8'hf0;
  assign T217 = T218 << 3'h4;
  assign T218 = T219[2'h3:1'h0];
  assign T219 = T12[3'h7:1'h0];
  assign T220 = T547 & 8'hf;
  assign T547 = {4'h0, T221};
  assign T221 = T219 >> 3'h4;
  assign T222 = T548 & 8'h33;
  assign T548 = {2'h0, T223};
  assign T223 = T215 >> 2'h2;
  assign T224 = T549 & 8'h55;
  assign T549 = {1'h0, T225};
  assign T225 = T211 >> 1'h1;
  assign T226 = T249 | T227;
  assign T227 = T228 & 16'haaaa;
  assign T228 = T229 << 1'h1;
  assign T229 = T230[4'he:1'h0];
  assign T230 = T247 | T231;
  assign T231 = T232 & 16'hcccc;
  assign T232 = T233 << 2'h2;
  assign T233 = T234[4'hd:1'h0];
  assign T234 = T245 | T235;
  assign T235 = T236 & 16'hf0f0;
  assign T236 = T237 << 3'h4;
  assign T237 = T238[4'hb:1'h0];
  assign T238 = T243 | T239;
  assign T239 = T240 & 16'hff00;
  assign T240 = T241 << 4'h8;
  assign T241 = T242[3'h7:1'h0];
  assign T242 = T13[4'hf:1'h0];
  assign T243 = T550 & 16'hff;
  assign T550 = {8'h0, T244};
  assign T244 = T242 >> 4'h8;
  assign T245 = T551 & 16'hf0f;
  assign T551 = {4'h0, T246};
  assign T246 = T238 >> 3'h4;
  assign T247 = T552 & 16'h3333;
  assign T552 = {2'h0, T248};
  assign T248 = T234 >> 2'h2;
  assign T249 = T553 & 16'h5555;
  assign T553 = {1'h0, T250};
  assign T250 = T230 >> 1'h1;
  assign T251 = 27'h0 - T554;
  assign T554 = {26'h0, T252};
  assign T252 = sExpX3[4'ha:4'ha];
  assign sigX3 = T253[5'h1b:1'h0];
  assign T253 = {T380, T254};
  assign T254 = doIncrSig ? T376 : T255;
  assign T255 = T256 != 16'h0;
  assign T256 = T299 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T257, 1'h1};
  assign T257 = {T280, T258};
  assign T258 = {T270, T259};
  assign T259 = {T266, T260};
  assign T260 = T261[2'h2:2'h2];
  assign T261 = T262[3'h6:3'h4];
  assign T262 = T263[4'he:4'h8];
  assign T263 = T264[4'hf:1'h1];
  assign T264 = $signed(17'h10000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T265;
  assign T265 = estNormDist[2'h3:1'h0];
  assign T266 = {T269, T267};
  assign T267 = T268[1'h1:1'h1];
  assign T268 = T261[1'h1:1'h0];
  assign T269 = T268[1'h0:1'h0];
  assign T270 = {T276, T271};
  assign T271 = {T275, T272};
  assign T272 = T273[1'h1:1'h1];
  assign T273 = T274[2'h3:2'h2];
  assign T274 = T262[2'h3:1'h0];
  assign T275 = T273[1'h0:1'h0];
  assign T276 = {T279, T277};
  assign T277 = T278[1'h1:1'h1];
  assign T278 = T274[1'h1:1'h0];
  assign T279 = T278[1'h0:1'h0];
  assign T280 = T297 | T281;
  assign T281 = T282 & 8'haa;
  assign T282 = T283 << 1'h1;
  assign T283 = T284[3'h6:1'h0];
  assign T284 = T295 | T285;
  assign T285 = T286 & 8'hcc;
  assign T286 = T287 << 2'h2;
  assign T287 = T288[3'h5:1'h0];
  assign T288 = T293 | T289;
  assign T289 = T290 & 8'hf0;
  assign T290 = T291 << 3'h4;
  assign T291 = T292[2'h3:1'h0];
  assign T292 = T263[3'h7:1'h0];
  assign T293 = T555 & 8'hf;
  assign T555 = {4'h0, T294};
  assign T294 = T292 >> 3'h4;
  assign T295 = T556 & 8'h33;
  assign T556 = {2'h0, T296};
  assign T296 = T288 >> 2'h2;
  assign T297 = T557 & 8'h55;
  assign T557 = {1'h0, T298};
  assign T298 = T284 >> 1'h1;
  assign T299 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T362 : T558;
  assign T558 = {1'h0, T300};
  assign T300 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T326 ? T320 : T301;
  assign T301 = T319 ? T560 : T302;
  assign T302 = {T304, T303};
  assign T303 = 32'h0 - T559;
  assign T559 = {31'h0, doSubMags};
  assign T304 = sigSum[4'ha:1'h1];
  assign T560 = {8'h0, T305};
  assign T305 = {T318, T306};
  assign T306 = doSubMags ? T312 : T307;
  assign T307 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T310, T308};
  assign T308 = T309 != 18'h0;
  assign T309 = sigSum[5'h11:1'h0];
  assign T310 = T311 != 16'h0;
  assign T311 = sigSum[6'h21:5'h12];
  assign T312 = ~ T313;
  assign T313 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T316, T314};
  assign T314 = T315 != 18'h0;
  assign T315 = notSigSum[5'h11:1'h0];
  assign notSigSum = ~ sigSum;
  assign T316 = T317 != 16'h0;
  assign T317 = notSigSum[6'h21:5'h12];
  assign T318 = sigSum[6'h32:5'h12];
  assign T319 = estNormNeg_dist[3'h4:3'h4];
  assign T320 = T325 ? T322 : T321;
  assign T321 = sigSum[6'h2a:1'h1];
  assign T322 = {T324, T323};
  assign T323 = 16'h0 - T561;
  assign T561 = {15'h0, doSubMags};
  assign T324 = sigSum[5'h1a:1'h1];
  assign T325 = estNormNeg_dist[3'h4:3'h4];
  assign T326 = estNormNeg_dist[3'h5:3'h5];
  assign CDom_firstNormAbsSigSum = T327;
  assign T327 = T335 | T328;
  assign T328 = T562 & T329;
  assign T329 = {T331, T330};
  assign T330 = firstReduceNotSigSum[1'h0:1'h0];
  assign T331 = notSigSum[6'h3a:5'h12];
  assign T562 = T332 ? 42'h3ffffffffff : 42'h0;
  assign T332 = T333;
  assign T333 = doSubMags & T334;
  assign T334 = CDom_estNormDist[3'h4:3'h4];
  assign T335 = T344 | T336;
  assign T336 = T563 & T337;
  assign T337 = {T339, T338};
  assign T338 = firstReduceNotSigSum != 2'h0;
  assign T339 = notSigSum[7'h4a:6'h22];
  assign T563 = T340 ? 42'h3ffffffffff : 42'h0;
  assign T340 = T341;
  assign T341 = doSubMags & T342;
  assign T342 = ~ T343;
  assign T343 = CDom_estNormDist[3'h4:3'h4];
  assign T344 = T353 | T345;
  assign T345 = T564 & T346;
  assign T346 = {T348, T347};
  assign T347 = firstReduceSigSum[1'h0:1'h0];
  assign T348 = sigSum[6'h3a:5'h12];
  assign T564 = T349 ? 42'h3ffffffffff : 42'h0;
  assign T349 = T350;
  assign T350 = T352 & T351;
  assign T351 = CDom_estNormDist[3'h4:3'h4];
  assign T352 = ~ doSubMags;
  assign T353 = T565 & T354;
  assign T354 = {T356, T355};
  assign T355 = firstReduceSigSum != 2'h0;
  assign T356 = sigSum[7'h4a:6'h22];
  assign T565 = T357 ? 42'h3ffffffffff : 42'h0;
  assign T357 = T358;
  assign T358 = T361 & T359;
  assign T359 = ~ T360;
  assign T360 = CDom_estNormDist[3'h4:3'h4];
  assign T361 = ~ doSubMags;
  assign T362 = isCDominant ? T568 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T375 ? T370 : T363;
  assign T363 = T369 ? T566 : T364;
  assign T364 = T365 << 6'h20;
  assign T365 = notSigSum[4'hb:1'h1];
  assign T566 = {10'h0, T366};
  assign T366 = {T368, T367};
  assign T367 = firstReduceNotSigSum[1'h0:1'h0];
  assign T368 = notSigSum[6'h31:5'h12];
  assign T369 = estNormNeg_dist[3'h4:3'h4];
  assign T370 = T374 ? T372 : T567;
  assign T567 = {1'h0, T371};
  assign T371 = notSigSum[6'h2a:1'h1];
  assign T372 = T373 << 5'h10;
  assign T373 = notSigSum[5'h1b:1'h1];
  assign T374 = estNormNeg_dist[3'h4:3'h4];
  assign T375 = estNormNeg_dist[3'h5:3'h5];
  assign T568 = {1'h0, CDom_firstNormAbsSigSum};
  assign T376 = T377 == 16'h0;
  assign T377 = T378 & absSigSumExtraMask;
  assign T378 = ~ T379;
  assign T379 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign T380 = T381 >> normTo2ShiftDist;
  assign T381 = cFirstNormAbsSigSum[6'h2a:1'h1];
  assign roundPosBit = T382 != 28'h0;
  assign T382 = sigX3 & T569;
  assign T569 = {1'h0, roundPosMask};
  assign roundPosMask = T570 & roundMask;
  assign T570 = {1'h0, T383};
  assign T383 = ~ T384;
  assign T384 = roundMask >> 1'h1;
  assign T385 = ~ allRound;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T386 == 28'h0;
  assign T386 = T388 & T571;
  assign T571 = {2'h0, T387};
  assign T387 = roundMask >> 1'h1;
  assign T388 = ~ sigX3;
  assign doIncrSig = T389 & doSubMags;
  assign T389 = T391 & T390;
  assign T390 = ~ notCDom_signSigSum;
  assign T391 = ~ isCDominant;
  assign commonCase = T393 & T392;
  assign T392 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T393 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T394 == 2'h3;
  assign T394 = expC[4'h8:3'h7];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T395 == 2'h3;
  assign T395 = expB[4'h8:3'h7];
  assign isSpecialA = T396 == 2'h3;
  assign T396 = expA[4'h8:3'h7];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T397;
  assign T397 = T401 | T398;
  assign T398 = sExpX3_13 <= T572;
  assign T572 = {2'h0, T399};
  assign T399 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign sigX3Shift1 = T400 == 2'h0;
  assign T400 = sigX3[5'h1b:5'h1a];
  assign T401 = sExpX3[4'ha:4'ha];
  assign overflow = commonCase & overflowY;
  assign overflowY = T402 == 3'h3;
  assign T402 = sExpY[4'h9:3'h7];
  assign sExpY = T449 | T403;
  assign T403 = T405 ? T404 : 11'h0;
  assign T404 = sExpX3 - 11'h1;
  assign T405 = T406 == 2'h0;
  assign T406 = sigY3[5'h19:5'h18];
  assign sigY3 = T420 | T407;
  assign T407 = roundEven ? T408 : 26'h0;
  assign T408 = roundUp_sigY3 & T409;
  assign T409 = ~ T410;
  assign T410 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T411[5'h19:1'h0];
  assign T411 = T412 + 26'h1;
  assign T412 = T413 >> 2'h2;
  assign T413 = sigX3 | T573;
  assign T573 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T417 : T414;
  assign T414 = T416 & T415;
  assign T415 = ~ anyRoundExtra;
  assign T416 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T417 = T418 & allRoundExtra;
  assign T418 = roundingMode_nearest_even & T419;
  assign T419 = ~ roundPosBit;
  assign T420 = T442 | T421;
  assign T421 = roundUp ? roundUp_sigY3 : 26'h0;
  assign roundUp = T429 | T422;
  assign T422 = T423 & 1'h1;
  assign T423 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T427 & T424;
  assign T424 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T425 : notCDom_signSigSum;
  assign T425 = doSubMags & T426;
  assign T426 = ~ isZeroC;
  assign T427 = ~ isZeroY;
  assign isZeroY = T428 == 3'h0;
  assign T428 = sigX3[5'h1b:5'h19];
  assign T429 = T432 | T430;
  assign T430 = T431 & roundPosBit;
  assign T431 = doIncrSig & roundingMode_nearest_even;
  assign T432 = T434 | T433;
  assign T433 = doIncrSig & allRound;
  assign T434 = T438 | T435;
  assign T435 = T436 & anyRound;
  assign T436 = T437 & roundDirectUp;
  assign T437 = ~ doIncrSig;
  assign T438 = T439 & anyRoundExtra;
  assign T439 = T440 & roundPosBit;
  assign T440 = T441 & roundingMode_nearest_even;
  assign T441 = ~ doIncrSig;
  assign T442 = T446 ? T443 : 26'h0;
  assign T443 = T444 >> 2'h2;
  assign T444 = sigX3 & T574;
  assign T574 = {1'h0, T445};
  assign T445 = ~ roundMask;
  assign T446 = T448 & T447;
  assign T447 = ~ roundEven;
  assign T448 = ~ roundUp;
  assign T449 = T452 | T450;
  assign T450 = T451 ? sExpX3 : 11'h0;
  assign T451 = sigY3[5'h18:5'h18];
  assign T452 = T454 ? T453 : 11'h0;
  assign T453 = sExpX3 + 11'h1;
  assign T454 = sigY3[5'h19:5'h19];
  assign T455 = {invalid, 1'h0};
  assign invalid = T474 | notSigNaN_invalid;
  assign notSigNaN_invalid = T471 | T456;
  assign T456 = T457 & doSubMags;
  assign T457 = T460 & isInfC;
  assign isInfC = isSpecialC & T458;
  assign T458 = T459 ^ 1'h1;
  assign T459 = expC[3'h6:3'h6];
  assign T460 = T466 & T461;
  assign T461 = isInfA | isInfB;
  assign isInfB = isSpecialB & T462;
  assign T462 = T463 ^ 1'h1;
  assign T463 = expB[3'h6:3'h6];
  assign isInfA = isSpecialA & T464;
  assign T464 = T465 ^ 1'h1;
  assign T465 = expA[3'h6:3'h6];
  assign T466 = T469 & T467;
  assign T467 = ~ isNaNB;
  assign isNaNB = isSpecialB & T468;
  assign T468 = expB[3'h6:3'h6];
  assign T469 = ~ isNaNA;
  assign isNaNA = isSpecialA & T470;
  assign T470 = expA[3'h6:3'h6];
  assign T471 = T473 | T472;
  assign T472 = isZeroA & isInfB;
  assign T473 = isInfA & isZeroB;
  assign T474 = T478 | isSigNaNC;
  assign isSigNaNC = isNaNC & T475;
  assign T475 = T476 ^ 1'h1;
  assign T476 = fractC[5'h16:5'h16];
  assign isNaNC = isSpecialC & T477;
  assign T477 = expC[3'h6:3'h6];
  assign T478 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T479;
  assign T479 = T480 ^ 1'h1;
  assign T480 = fractB[5'h16:5'h16];
  assign isSigNaNA = isNaNA & T481;
  assign T481 = T482 ^ 1'h1;
  assign T482 = fractA[5'h16:5'h16];
  assign io_out = T483;
  assign T483 = {signOut, T484};
  assign T484 = {expOut, fractOut};
  assign fractOut = fractY | T485;
  assign T485 = 23'h0 - T575;
  assign T575 = {22'h0, T486};
  assign T486 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T487;
  assign T487 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T490 | T488;
  assign T488 = roundingMode_max & T489;
  assign T489 = ~ signY;
  assign T490 = roundingMode_nearest_even | T491;
  assign T491 = roundingMode_min & signY;
  assign isNaNOut = T492 | notSigNaN_invalid;
  assign T492 = T493 | isNaNC;
  assign T493 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T495 : T494;
  assign T494 = sigY3[5'h17:1'h1];
  assign T495 = sigY3[5'h16:1'h0];
  assign expOut = T497 | T496;
  assign T496 = isNaNOut ? 9'h1c0 : 9'h0;
  assign T497 = T502 | T498;
  assign T498 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign notNaN_isInfOut = T500 | T499;
  assign T499 = overflow & overflowY_roundMagUp;
  assign T500 = T501 | isInfC;
  assign T501 = isInfA | isInfB;
  assign T502 = T504 | T503;
  assign T503 = isSatOut ? 9'h17f : 9'h0;
  assign T504 = T507 & T505;
  assign T505 = ~ T506;
  assign T506 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T507 = T510 & T508;
  assign T508 = ~ T509;
  assign T509 = isSatOut ? 9'h80 : 9'h0;
  assign T510 = expY & T511;
  assign T511 = ~ T512;
  assign T512 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign notSpecial_isZeroOut = T516 | totalUnderflowY;
  assign totalUnderflowY = T515 | T513;
  assign T513 = T514 < 9'h6b;
  assign T514 = sExpY[4'h8:1'h0];
  assign T515 = sExpY[4'h9:4'h9];
  assign T516 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'h8:1'h0];
  assign signOut = T518 | T517;
  assign T517 = commonCase & signY;
  assign T518 = T522 | T519;
  assign T519 = T520 & opSignC;
  assign T520 = T521 & isSpecialC;
  assign T521 = mulSpecial ^ 1'h1;
  assign T522 = T526 | T523;
  assign T523 = T524 & signProd;
  assign T524 = mulSpecial & T525;
  assign T525 = isSpecialC ^ 1'h1;
  assign T526 = T527 | isNaNOut;
  assign T527 = T528 & opSignC;
  assign T528 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_0(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T7;
  reg [2:0] in_rm;
  wire[2:0] T8;
  wire[32:0] T9;
  reg [64:0] in_in3;
  wire[64:0] T10;
  wire[64:0] T11;
  wire[64:0] T12;
  wire[32:0] zero;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[32:0] T19;
  reg [64:0] in_in2;
  wire[64:0] T20;
  wire[64:0] T21;
  wire T22;
  wire[32:0] T23;
  reg [64:0] in_in1;
  wire[64:0] T24;
  wire[1:0] T25;
  reg [4:0] in_cmd;
  wire[4:0] T26;
  wire[4:0] T27;
  wire[4:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg [4:0] R0;
  wire[4:0] T1;
  wire[4:0] res_exc;
  reg  valid;
  reg [64:0] R2;
  wire[64:0] T3;
  wire[64:0] res_data;
  wire[64:0] T5;
  reg  R4;
  wire T6;
  wire[32:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R0 = {1{$random}};
    valid = {1{$random}};
    R2 = {3{$random}};
    R4 = {1{$random}};
  end
`endif

  assign T7 = in_rm[1'h1:1'h0];
  assign T8 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T9 = in_in3[6'h20:1'h0];
  assign T10 = T16 ? T12 : T11;
  assign T11 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T12 = {32'h0, zero};
  assign zero = T13 << 6'h20;
  assign T13 = T15 ^ T14;
  assign T14 = io_in_bits_in2[6'h20:6'h20];
  assign T15 = io_in_bits_in1[6'h20:6'h20];
  assign T16 = io_in_valid & T17;
  assign T17 = T18 ^ 1'h1;
  assign T18 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T19 = in_in2[6'h20:1'h0];
  assign T20 = T22 ? 65'h80000000 : T21;
  assign T21 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T22 = io_in_valid & io_in_bits_swap23;
  assign T23 = in_in1[6'h20:1'h0];
  assign T24 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T25 = in_cmd[1'h1:1'h0];
  assign T26 = io_in_valid ? T28 : T27;
  assign T27 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T28 = {3'h0, T29};
  assign T29 = {T31, T30};
  assign T30 = io_in_bits_cmd[1'h0:1'h0];
  assign T31 = T33 & T32;
  assign T32 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T33 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R0;
  assign T1 = valid ? res_exc : R0;
  assign res_exc = fma_io_exceptionFlags;
  assign io_out_bits_data = R2;
  assign T3 = valid ? res_data : R2;
  assign res_data = T5;
  assign T5 = {32'h0, fma_io_out};
  assign io_out_valid = R4;
  assign T6 = reset ? 1'h0 : valid;
  mulAddSubRecodedFloatN_0 fma(
       .io_op( T25 ),
       .io_a( T23 ),
       .io_b( T19 ),
       .io_c( T9 ),
       .io_roundingMode( T7 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T16) begin
      in_in3 <= T12;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T22) begin
      in_in2 <= 65'h80000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T28;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(valid) begin
      R0 <= res_exc;
    end
    valid <= io_in_valid;
    if(valid) begin
      R2 <= res_data;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else begin
      R4 <= valid;
    end
  end
endmodule

module mulAddSubRecodedFloatN_1(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[56:0] T4;
  wire[56:0] T744;
  wire[54:0] T5;
  wire[55:0] roundMask;
  wire[55:0] T6;
  wire[53:0] T7;
  wire[53:0] T745;
  wire T8;
  wire[53:0] T9;
  wire[21:0] T10;
  wire[5:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[5:0] T15;
  wire[21:0] T16;
  wire[53:0] T17;
  wire[8192:0] T18;
  wire[12:0] T19;
  wire[12:0] sExpX3_13;
  wire[13:0] sExpX3;
  wire[13:0] T746;
  wire[7:0] estNormDist;
  wire[7:0] T20;
  wire[7:0] estNormNeg_dist;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[7:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[7:0] T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[7:0] T58;
  wire[7:0] T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire[7:0] T75;
  wire[7:0] T76;
  wire[7:0] T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire[7:0] T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T119;
  wire[7:0] T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire T127;
  wire[108:0] T128;
  wire[108:0] T129;
  wire[107:0] T130;
  wire[107:0] T131;
  wire[161:0] sigSum;
  wire[161:0] alignedNegSigC;
  wire[162:0] T132;
  wire T133;
  wire doSubMags;
  wire opSignC;
  wire T134;
  wire T135;
  wire signProd;
  wire T136;
  wire T137;
  wire signB;
  wire signA;
  wire T138;
  wire[52:0] T139;
  wire[52:0] CExtraMask;
  wire[20:0] T140;
  wire[4:0] T141;
  wire T142;
  wire[4:0] T143;
  wire[20:0] T144;
  wire[52:0] T145;
  wire[256:0] T146;
  wire[7:0] CAlignDist;
  wire[13:0] T147;
  wire[13:0] T148;
  wire[13:0] sNatCAlignDist;
  wire[13:0] T747;
  wire[11:0] expC;
  wire[13:0] sExpAlignedProd;
  wire[13:0] T149;
  wire[13:0] T748;
  wire[11:0] expA;
  wire[13:0] T150;
  wire[10:0] T151;
  wire[11:0] expB;
  wire[2:0] T152;
  wire[2:0] T749;
  wire T153;
  wire T154;
  wire T155;
  wire[12:0] T156;
  wire CAlignDist_floor;
  wire T157;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T158;
  wire isZeroA;
  wire[2:0] T159;
  wire[3:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[1:0] T163;
  wire[3:0] T164;
  wire T165;
  wire[1:0] T166;
  wire T167;
  wire[1:0] T168;
  wire T169;
  wire[15:0] T170;
  wire[15:0] T171;
  wire[15:0] T172;
  wire[14:0] T173;
  wire[15:0] T174;
  wire[15:0] T175;
  wire[15:0] T176;
  wire[13:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[15:0] T180;
  wire[11:0] T181;
  wire[15:0] T182;
  wire[15:0] T183;
  wire[15:0] T184;
  wire[7:0] T185;
  wire[15:0] T186;
  wire[15:0] T187;
  wire[15:0] T750;
  wire[7:0] T188;
  wire[15:0] T189;
  wire[15:0] T751;
  wire[11:0] T190;
  wire[15:0] T191;
  wire[15:0] T752;
  wire[13:0] T192;
  wire[15:0] T193;
  wire[15:0] T753;
  wire[14:0] T194;
  wire[31:0] T195;
  wire[31:0] T196;
  wire[31:0] T197;
  wire[30:0] T198;
  wire[31:0] T199;
  wire[31:0] T200;
  wire[31:0] T201;
  wire[29:0] T202;
  wire[31:0] T203;
  wire[31:0] T204;
  wire[31:0] T205;
  wire[27:0] T206;
  wire[31:0] T207;
  wire[31:0] T208;
  wire[31:0] T209;
  wire[23:0] T210;
  wire[31:0] T211;
  wire[31:0] T212;
  wire[31:0] T213;
  wire[15:0] T214;
  wire[31:0] T215;
  wire[31:0] T216;
  wire[31:0] T754;
  wire[15:0] T217;
  wire[31:0] T218;
  wire[31:0] T755;
  wire[23:0] T219;
  wire[31:0] T220;
  wire[31:0] T756;
  wire[27:0] T221;
  wire[31:0] T222;
  wire[31:0] T757;
  wire[29:0] T223;
  wire[31:0] T224;
  wire[31:0] T758;
  wire[30:0] T225;
  wire[52:0] sigC;
  wire[51:0] fractC;
  wire T226;
  wire isZeroC;
  wire[2:0] T227;
  wire[161:0] T228;
  wire[161:0] T229;
  wire[161:0] T230;
  wire[160:0] T231;
  wire[107:0] T232;
  wire[107:0] T759;
  wire[52:0] negSigC;
  wire[52:0] T233;
  wire[161:0] T760;
  wire[106:0] T234;
  wire[105:0] T235;
  wire[52:0] sigB;
  wire[51:0] fractB;
  wire T236;
  wire[52:0] sigA;
  wire[51:0] fractA;
  wire T237;
  wire[108:0] T761;
  wire[107:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire notCDom_signSigSum;
  wire[7:0] CDom_estNormDist;
  wire[7:0] T762;
  wire[5:0] T345;
  wire[7:0] T346;
  wire T347;
  wire CAlignDist_0;
  wire T348;
  wire[12:0] T349;
  wire isCDominant;
  wire T350;
  wire T351;
  wire[12:0] T352;
  wire T353;
  wire[13:0] sExpSum;
  wire[13:0] T763;
  wire T354;
  wire[3:0] T355;
  wire[1:0] T356;
  wire T357;
  wire[1:0] T358;
  wire[3:0] T359;
  wire T360;
  wire[1:0] T361;
  wire T362;
  wire[1:0] T363;
  wire T364;
  wire[15:0] T365;
  wire[15:0] T366;
  wire[15:0] T367;
  wire[14:0] T368;
  wire[15:0] T369;
  wire[15:0] T370;
  wire[15:0] T371;
  wire[13:0] T372;
  wire[15:0] T373;
  wire[15:0] T374;
  wire[15:0] T375;
  wire[11:0] T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[7:0] T380;
  wire[15:0] T381;
  wire[15:0] T382;
  wire[15:0] T764;
  wire[7:0] T383;
  wire[15:0] T384;
  wire[15:0] T765;
  wire[11:0] T385;
  wire[15:0] T386;
  wire[15:0] T766;
  wire[13:0] T387;
  wire[15:0] T388;
  wire[15:0] T767;
  wire[14:0] T389;
  wire[31:0] T390;
  wire[31:0] T391;
  wire[31:0] T392;
  wire[30:0] T393;
  wire[31:0] T394;
  wire[31:0] T395;
  wire[31:0] T396;
  wire[29:0] T397;
  wire[31:0] T398;
  wire[31:0] T399;
  wire[31:0] T400;
  wire[27:0] T401;
  wire[31:0] T402;
  wire[31:0] T403;
  wire[31:0] T404;
  wire[23:0] T405;
  wire[31:0] T406;
  wire[31:0] T407;
  wire[31:0] T408;
  wire[15:0] T409;
  wire[31:0] T410;
  wire[31:0] T411;
  wire[31:0] T768;
  wire[15:0] T412;
  wire[31:0] T413;
  wire[31:0] T769;
  wire[23:0] T414;
  wire[31:0] T415;
  wire[31:0] T770;
  wire[27:0] T416;
  wire[31:0] T417;
  wire[31:0] T771;
  wire[29:0] T418;
  wire[31:0] T419;
  wire[31:0] T772;
  wire[30:0] T420;
  wire[55:0] T421;
  wire[55:0] T773;
  wire T422;
  wire[56:0] sigX3;
  wire[87:0] T423;
  wire T424;
  wire T425;
  wire[31:0] T426;
  wire[31:0] absSigSumExtraMask;
  wire[30:0] T427;
  wire[14:0] T428;
  wire[6:0] T429;
  wire[2:0] T430;
  wire T431;
  wire[2:0] T432;
  wire[6:0] T433;
  wire[14:0] T434;
  wire[30:0] T435;
  wire[32:0] T436;
  wire[4:0] normTo2ShiftDist;
  wire[4:0] estNormDist_5;
  wire[4:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[1:0] T440;
  wire T441;
  wire[3:0] T442;
  wire[1:0] T443;
  wire T444;
  wire[1:0] T445;
  wire[3:0] T446;
  wire T447;
  wire[1:0] T448;
  wire T449;
  wire[1:0] T450;
  wire T451;
  wire[7:0] T452;
  wire[7:0] T453;
  wire[7:0] T454;
  wire[6:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[5:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[3:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T774;
  wire[3:0] T466;
  wire[7:0] T467;
  wire[7:0] T775;
  wire[5:0] T468;
  wire[7:0] T469;
  wire[7:0] T776;
  wire[6:0] T470;
  wire[15:0] T471;
  wire[15:0] T472;
  wire[15:0] T473;
  wire[14:0] T474;
  wire[15:0] T475;
  wire[15:0] T476;
  wire[15:0] T477;
  wire[13:0] T478;
  wire[15:0] T479;
  wire[15:0] T480;
  wire[15:0] T481;
  wire[11:0] T482;
  wire[15:0] T483;
  wire[15:0] T484;
  wire[15:0] T485;
  wire[7:0] T486;
  wire[15:0] T487;
  wire[15:0] T488;
  wire[15:0] T777;
  wire[7:0] T489;
  wire[15:0] T490;
  wire[15:0] T778;
  wire[11:0] T491;
  wire[15:0] T492;
  wire[15:0] T779;
  wire[13:0] T493;
  wire[15:0] T494;
  wire[15:0] T780;
  wire[14:0] T495;
  wire[31:0] T496;
  wire[87:0] cFirstNormAbsSigSum;
  wire[87:0] T781;
  wire[86:0] T497;
  wire[86:0] notCDom_pos_firstNormAbsSigSum;
  wire[86:0] T498;
  wire[86:0] T499;
  wire[53:0] T500;
  wire[53:0] T782;
  wire[32:0] T501;
  wire[86:0] T502;
  wire[86:0] T503;
  wire[85:0] T504;
  wire[85:0] T783;
  wire T505;
  wire[86:0] T784;
  wire[65:0] T506;
  wire T507;
  wire T508;
  wire[1:0] firstReduceSigSum;
  wire T509;
  wire[43:0] T510;
  wire T511;
  wire[31:0] T512;
  wire T513;
  wire T514;
  wire[1:0] firstReduceNotSigSum;
  wire T515;
  wire[43:0] T516;
  wire[161:0] notSigSum;
  wire T517;
  wire[31:0] T518;
  wire[64:0] T519;
  wire T520;
  wire T521;
  wire[86:0] T522;
  wire[86:0] T523;
  wire T524;
  wire T525;
  wire[10:0] T526;
  wire T527;
  wire[10:0] T528;
  wire[85:0] T529;
  wire[86:0] T530;
  wire[21:0] T531;
  wire[21:0] T785;
  wire[64:0] T532;
  wire T533;
  wire T534;
  wire[86:0] CDom_firstNormAbsSigSum;
  wire[86:0] T535;
  wire[86:0] T536;
  wire[86:0] T537;
  wire T538;
  wire[85:0] T539;
  wire[86:0] T786;
  wire T540;
  wire T541;
  wire T542;
  wire[86:0] T543;
  wire[86:0] T544;
  wire[86:0] T545;
  wire T546;
  wire[85:0] T547;
  wire[86:0] T787;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire[86:0] T552;
  wire[86:0] T553;
  wire[86:0] T554;
  wire T555;
  wire[85:0] T556;
  wire[86:0] T788;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire[86:0] T561;
  wire[86:0] T562;
  wire T563;
  wire[85:0] T564;
  wire[86:0] T789;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire[87:0] T570;
  wire[87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[87:0] T571;
  wire[87:0] T572;
  wire[33:0] T573;
  wire[87:0] T574;
  wire[87:0] T575;
  wire[1:0] T576;
  wire[87:0] T790;
  wire[64:0] T577;
  wire T578;
  wire[63:0] T579;
  wire T580;
  wire T581;
  wire[87:0] T582;
  wire[87:0] T583;
  wire T584;
  wire[10:0] T585;
  wire[86:0] T586;
  wire[87:0] T587;
  wire[65:0] T588;
  wire T589;
  wire T590;
  wire[87:0] T791;
  wire T591;
  wire[31:0] T592;
  wire[31:0] T593;
  wire[31:0] T594;
  wire[86:0] T595;
  wire[86:0] T596;
  wire roundPosBit;
  wire[56:0] T597;
  wire[56:0] T792;
  wire[55:0] roundPosMask;
  wire[55:0] T793;
  wire[54:0] T598;
  wire[54:0] T599;
  wire T600;
  wire allRound;
  wire allRoundExtra;
  wire[56:0] T601;
  wire[56:0] T794;
  wire[54:0] T602;
  wire[56:0] T603;
  wire doIncrSig;
  wire T604;
  wire T605;
  wire T606;
  wire commonCase;
  wire T607;
  wire notSpecial_addZeros;
  wire T608;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T609;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T610;
  wire isSpecialA;
  wire[1:0] T611;
  wire underflow;
  wire underflowY;
  wire T612;
  wire T613;
  wire[12:0] T795;
  wire[10:0] T614;
  wire sigX3Shift1;
  wire[1:0] T615;
  wire T616;
  wire overflow;
  wire overflowY;
  wire[2:0] T617;
  wire[13:0] sExpY;
  wire[13:0] T618;
  wire[13:0] T619;
  wire T620;
  wire[1:0] T621;
  wire[54:0] sigY3;
  wire[54:0] T622;
  wire[54:0] T623;
  wire[54:0] T624;
  wire[54:0] T625;
  wire[54:0] roundUp_sigY3;
  wire[54:0] T626;
  wire[54:0] T627;
  wire[56:0] T628;
  wire[56:0] T796;
  wire roundEven;
  wire T629;
  wire T630;
  wire T631;
  wire roundingMode_nearest_even;
  wire T632;
  wire T633;
  wire T634;
  wire[54:0] T635;
  wire[54:0] T636;
  wire roundUp;
  wire T637;
  wire T638;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T639;
  wire doNegSignSum;
  wire T640;
  wire T641;
  wire T642;
  wire isZeroY;
  wire[2:0] T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire[54:0] T657;
  wire[54:0] T658;
  wire[56:0] T659;
  wire[56:0] T797;
  wire[55:0] T660;
  wire T661;
  wire T662;
  wire T663;
  wire[13:0] T664;
  wire[13:0] T665;
  wire T666;
  wire[13:0] T667;
  wire[13:0] T668;
  wire T669;
  wire[1:0] T670;
  wire invalid;
  wire notSigNaN_invalid;
  wire T671;
  wire T672;
  wire isInfC;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire isInfB;
  wire T677;
  wire T678;
  wire isInfA;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire isNaNB;
  wire T683;
  wire T684;
  wire isNaNA;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire isSigNaNC;
  wire T690;
  wire T691;
  wire isNaNC;
  wire T692;
  wire T693;
  wire isSigNaNB;
  wire T694;
  wire T695;
  wire isSigNaNA;
  wire T696;
  wire T697;
  wire[64:0] T698;
  wire[63:0] T699;
  wire[51:0] fractOut;
  wire[51:0] T700;
  wire[51:0] T798;
  wire T701;
  wire isSatOut;
  wire T702;
  wire overflowY_roundMagUp;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire isNaNOut;
  wire T707;
  wire T708;
  wire[51:0] fractY;
  wire[51:0] T709;
  wire[51:0] T710;
  wire[11:0] expOut;
  wire[11:0] T711;
  wire[11:0] T712;
  wire[11:0] T713;
  wire notNaN_isInfOut;
  wire T714;
  wire T715;
  wire T716;
  wire[11:0] T717;
  wire[11:0] T718;
  wire[11:0] T719;
  wire[11:0] T720;
  wire[11:0] T721;
  wire[11:0] T722;
  wire[11:0] T723;
  wire[11:0] T724;
  wire[11:0] T725;
  wire[11:0] T726;
  wire[11:0] T727;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T728;
  wire[11:0] T729;
  wire T730;
  wire T731;
  wire[11:0] expY;
  wire signOut;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;


  assign io_exceptionFlags = T0;
  assign T0 = {T670, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T600 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 57'h0;
  assign T4 = sigX3 & T744;
  assign T744 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T421 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T745;
  assign T745 = {53'h0, T8};
  assign T8 = sigX3[6'h37:6'h37];
  assign T9 = {T390, T10};
  assign T10 = {T365, T11};
  assign T11 = {T355, T12};
  assign T12 = {T354, T13};
  assign T13 = T14[1'h1:1'h1];
  assign T14 = T15[3'h5:3'h4];
  assign T15 = T16[5'h15:5'h10];
  assign T16 = T17[6'h35:6'h20];
  assign T17 = T18[11'h403:10'h3ce];
  assign T18 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T19;
  assign T19 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'hc:1'h0];
  assign sExpX3 = sExpSum - T746;
  assign T746 = {6'h0, estNormDist};
  assign estNormDist = isCDominant ? CDom_estNormDist : T20;
  assign T20 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = T344 ? 8'h35 : T21;
  assign T21 = T343 ? 8'h36 : T22;
  assign T22 = T342 ? 8'h37 : T23;
  assign T23 = T341 ? 8'h38 : T24;
  assign T24 = T340 ? 8'h39 : T25;
  assign T25 = T339 ? 8'h3a : T26;
  assign T26 = T338 ? 8'h3b : T27;
  assign T27 = T337 ? 8'h3c : T28;
  assign T28 = T336 ? 8'h3d : T29;
  assign T29 = T335 ? 8'h3e : T30;
  assign T30 = T334 ? 8'h3f : T31;
  assign T31 = T333 ? 8'h40 : T32;
  assign T32 = T332 ? 8'h41 : T33;
  assign T33 = T331 ? 8'h42 : T34;
  assign T34 = T330 ? 8'h43 : T35;
  assign T35 = T329 ? 8'h44 : T36;
  assign T36 = T328 ? 8'h45 : T37;
  assign T37 = T327 ? 8'h46 : T38;
  assign T38 = T326 ? 8'h47 : T39;
  assign T39 = T325 ? 8'h48 : T40;
  assign T40 = T324 ? 8'h49 : T41;
  assign T41 = T323 ? 8'h4a : T42;
  assign T42 = T322 ? 8'h4b : T43;
  assign T43 = T321 ? 8'h4c : T44;
  assign T44 = T320 ? 8'h4d : T45;
  assign T45 = T319 ? 8'h4e : T46;
  assign T46 = T318 ? 8'h4f : T47;
  assign T47 = T317 ? 8'h50 : T48;
  assign T48 = T316 ? 8'h51 : T49;
  assign T49 = T315 ? 8'h52 : T50;
  assign T50 = T314 ? 8'h53 : T51;
  assign T51 = T313 ? 8'h54 : T52;
  assign T52 = T312 ? 8'h55 : T53;
  assign T53 = T311 ? 8'h56 : T54;
  assign T54 = T310 ? 8'h57 : T55;
  assign T55 = T309 ? 8'h58 : T56;
  assign T56 = T308 ? 8'h59 : T57;
  assign T57 = T307 ? 8'h5a : T58;
  assign T58 = T306 ? 8'h5b : T59;
  assign T59 = T305 ? 8'h5c : T60;
  assign T60 = T304 ? 8'h5d : T61;
  assign T61 = T303 ? 8'h5e : T62;
  assign T62 = T302 ? 8'h5f : T63;
  assign T63 = T301 ? 8'h60 : T64;
  assign T64 = T300 ? 8'h61 : T65;
  assign T65 = T299 ? 8'h62 : T66;
  assign T66 = T298 ? 8'h63 : T67;
  assign T67 = T297 ? 8'h64 : T68;
  assign T68 = T296 ? 8'h65 : T69;
  assign T69 = T295 ? 8'h66 : T70;
  assign T70 = T294 ? 8'h67 : T71;
  assign T71 = T293 ? 8'h68 : T72;
  assign T72 = T292 ? 8'h69 : T73;
  assign T73 = T291 ? 8'h6a : T74;
  assign T74 = T290 ? 8'h6b : T75;
  assign T75 = T289 ? 8'h6c : T76;
  assign T76 = T288 ? 8'h6d : T77;
  assign T77 = T287 ? 8'h6e : T78;
  assign T78 = T286 ? 8'h6f : T79;
  assign T79 = T285 ? 8'h70 : T80;
  assign T80 = T284 ? 8'h71 : T81;
  assign T81 = T283 ? 8'h72 : T82;
  assign T82 = T282 ? 8'h73 : T83;
  assign T83 = T281 ? 8'h74 : T84;
  assign T84 = T280 ? 8'h75 : T85;
  assign T85 = T279 ? 8'h76 : T86;
  assign T86 = T278 ? 8'h77 : T87;
  assign T87 = T277 ? 8'h78 : T88;
  assign T88 = T276 ? 8'h79 : T89;
  assign T89 = T275 ? 8'h7a : T90;
  assign T90 = T274 ? 8'h7b : T91;
  assign T91 = T273 ? 8'h7c : T92;
  assign T92 = T272 ? 8'h7d : T93;
  assign T93 = T271 ? 8'h7e : T94;
  assign T94 = T270 ? 8'h7f : T95;
  assign T95 = T269 ? 8'h80 : T96;
  assign T96 = T268 ? 8'h81 : T97;
  assign T97 = T267 ? 8'h82 : T98;
  assign T98 = T266 ? 8'h83 : T99;
  assign T99 = T265 ? 8'h84 : T100;
  assign T100 = T264 ? 8'h85 : T101;
  assign T101 = T263 ? 8'h86 : T102;
  assign T102 = T262 ? 8'h87 : T103;
  assign T103 = T261 ? 8'h88 : T104;
  assign T104 = T260 ? 8'h89 : T105;
  assign T105 = T259 ? 8'h8a : T106;
  assign T106 = T258 ? 8'h8b : T107;
  assign T107 = T257 ? 8'h8c : T108;
  assign T108 = T256 ? 8'h8d : T109;
  assign T109 = T255 ? 8'h8e : T110;
  assign T110 = T254 ? 8'h8f : T111;
  assign T111 = T253 ? 8'h90 : T112;
  assign T112 = T252 ? 8'h91 : T113;
  assign T113 = T251 ? 8'h92 : T114;
  assign T114 = T250 ? 8'h93 : T115;
  assign T115 = T249 ? 8'h94 : T116;
  assign T116 = T248 ? 8'h95 : T117;
  assign T117 = T247 ? 8'h96 : T118;
  assign T118 = T246 ? 8'h97 : T119;
  assign T119 = T245 ? 8'h98 : T120;
  assign T120 = T244 ? 8'h99 : T121;
  assign T121 = T243 ? 8'h9a : T122;
  assign T122 = T242 ? 8'h9b : T123;
  assign T123 = T241 ? 8'h9c : T124;
  assign T124 = T240 ? 8'h9d : T125;
  assign T125 = T239 ? 8'h9e : T126;
  assign T126 = T127 ? 8'h9f : 8'ha0;
  assign T127 = T128[1'h1:1'h1];
  assign T128 = T761 ^ T129;
  assign T129 = T130 << 1'h1;
  assign T130 = 108'h0 | T131;
  assign T131 = sigSum[7'h6c:1'h1];
  assign sigSum = T760 + alignedNegSigC;
  assign alignedNegSigC = T132[8'ha1:1'h0];
  assign T132 = {T228, T133};
  assign T133 = T138 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T135 ^ T134;
  assign T134 = io_op[1'h0:1'h0];
  assign T135 = io_c[7'h40:7'h40];
  assign signProd = T137 ^ T136;
  assign T136 = io_op[1'h1:1'h1];
  assign T137 = signA ^ signB;
  assign signB = io_b[7'h40:7'h40];
  assign signA = io_a[7'h40:7'h40];
  assign T138 = T139 != 53'h0;
  assign T139 = sigC & CExtraMask;
  assign CExtraMask = {T195, T140};
  assign T140 = {T170, T141};
  assign T141 = {T160, T142};
  assign T142 = T143[3'h4:3'h4];
  assign T143 = T144[5'h14:5'h10];
  assign T144 = T145[6'h34:6'h20];
  assign T145 = T146[8'h93:7'h5f];
  assign T146 = $signed(257'h10000000000000000000000000000000000000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = T147[3'h7:1'h0];
  assign T147 = CAlignDist_floor ? 14'h0 : T148;
  assign T148 = T155 ? sNatCAlignDist : 14'ha1;
  assign sNatCAlignDist = sExpAlignedProd - T747;
  assign T747 = {2'h0, expC};
  assign expC = io_c[6'h3f:6'h34];
  assign sExpAlignedProd = T149 + 14'h38;
  assign T149 = T150 + T748;
  assign T748 = {2'h0, expA};
  assign expA = io_a[6'h3f:6'h34];
  assign T150 = {T152, T151};
  assign T151 = expB[4'ha:1'h0];
  assign expB = io_b[6'h3f:6'h34];
  assign T152 = 3'h0 - T749;
  assign T749 = {2'h0, T153};
  assign T153 = T154 ^ 1'h1;
  assign T154 = expB[4'hb:4'hb];
  assign T155 = T156 < 13'ha1;
  assign T156 = sNatCAlignDist[4'hc:1'h0];
  assign CAlignDist_floor = isZeroProd | T157;
  assign T157 = sNatCAlignDist[4'hd:4'hd];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T158 == 3'h0;
  assign T158 = expB[4'hb:4'h9];
  assign isZeroA = T159 == 3'h0;
  assign T159 = expA[4'hb:4'h9];
  assign T160 = {T166, T161};
  assign T161 = {T165, T162};
  assign T162 = T163[1'h1:1'h1];
  assign T163 = T164[2'h3:2'h2];
  assign T164 = T143[2'h3:1'h0];
  assign T165 = T163[1'h0:1'h0];
  assign T166 = {T169, T167};
  assign T167 = T168[1'h1:1'h1];
  assign T168 = T164[1'h1:1'h0];
  assign T169 = T168[1'h0:1'h0];
  assign T170 = T193 | T171;
  assign T171 = T172 & 16'haaaa;
  assign T172 = T173 << 1'h1;
  assign T173 = T174[4'he:1'h0];
  assign T174 = T191 | T175;
  assign T175 = T176 & 16'hcccc;
  assign T176 = T177 << 2'h2;
  assign T177 = T178[4'hd:1'h0];
  assign T178 = T189 | T179;
  assign T179 = T180 & 16'hf0f0;
  assign T180 = T181 << 3'h4;
  assign T181 = T182[4'hb:1'h0];
  assign T182 = T187 | T183;
  assign T183 = T184 & 16'hff00;
  assign T184 = T185 << 4'h8;
  assign T185 = T186[3'h7:1'h0];
  assign T186 = T144[4'hf:1'h0];
  assign T187 = T750 & 16'hff;
  assign T750 = {8'h0, T188};
  assign T188 = T186 >> 4'h8;
  assign T189 = T751 & 16'hf0f;
  assign T751 = {4'h0, T190};
  assign T190 = T182 >> 3'h4;
  assign T191 = T752 & 16'h3333;
  assign T752 = {2'h0, T192};
  assign T192 = T178 >> 2'h2;
  assign T193 = T753 & 16'h5555;
  assign T753 = {1'h0, T194};
  assign T194 = T174 >> 1'h1;
  assign T195 = T224 | T196;
  assign T196 = T197 & 32'haaaaaaaa;
  assign T197 = T198 << 1'h1;
  assign T198 = T199[5'h1e:1'h0];
  assign T199 = T222 | T200;
  assign T200 = T201 & 32'hcccccccc;
  assign T201 = T202 << 2'h2;
  assign T202 = T203[5'h1d:1'h0];
  assign T203 = T220 | T204;
  assign T204 = T205 & 32'hf0f0f0f0;
  assign T205 = T206 << 3'h4;
  assign T206 = T207[5'h1b:1'h0];
  assign T207 = T218 | T208;
  assign T208 = T209 & 32'hff00ff00;
  assign T209 = T210 << 4'h8;
  assign T210 = T211[5'h17:1'h0];
  assign T211 = T216 | T212;
  assign T212 = T213 & 32'hffff0000;
  assign T213 = T214 << 5'h10;
  assign T214 = T215[4'hf:1'h0];
  assign T215 = T145[5'h1f:1'h0];
  assign T216 = T754 & 32'hffff;
  assign T754 = {16'h0, T217};
  assign T217 = T215 >> 5'h10;
  assign T218 = T755 & 32'hff00ff;
  assign T755 = {8'h0, T219};
  assign T219 = T211 >> 4'h8;
  assign T220 = T756 & 32'hf0f0f0f;
  assign T756 = {4'h0, T221};
  assign T221 = T207 >> 3'h4;
  assign T222 = T757 & 32'h33333333;
  assign T757 = {2'h0, T223};
  assign T223 = T203 >> 2'h2;
  assign T224 = T758 & 32'h55555555;
  assign T758 = {1'h0, T225};
  assign T225 = T199 >> 1'h1;
  assign sigC = {T226, fractC};
  assign fractC = io_c[6'h33:1'h0];
  assign T226 = isZeroC ^ 1'h1;
  assign isZeroC = T227 == 3'h0;
  assign T227 = expC[4'hb:4'h9];
  assign T228 = $signed(T229) >>> CAlignDist;
  assign T229 = T230;
  assign T230 = {doSubMags, T231};
  assign T231 = {negSigC, T232};
  assign T232 = 108'h0 - T759;
  assign T759 = {107'h0, doSubMags};
  assign negSigC = doSubMags ? T233 : sigC;
  assign T233 = ~ sigC;
  assign T760 = {55'h0, T234};
  assign T234 = T235 << 1'h1;
  assign T235 = sigA * sigB;
  assign sigB = {T236, fractB};
  assign fractB = io_b[6'h33:1'h0];
  assign T236 = isZeroB ^ 1'h1;
  assign sigA = {T237, fractA};
  assign fractA = io_a[6'h33:1'h0];
  assign T237 = isZeroA ^ 1'h1;
  assign T761 = {1'h0, T238};
  assign T238 = 108'h0 ^ T131;
  assign T239 = T128[2'h2:2'h2];
  assign T240 = T128[2'h3:2'h3];
  assign T241 = T128[3'h4:3'h4];
  assign T242 = T128[3'h5:3'h5];
  assign T243 = T128[3'h6:3'h6];
  assign T244 = T128[3'h7:3'h7];
  assign T245 = T128[4'h8:4'h8];
  assign T246 = T128[4'h9:4'h9];
  assign T247 = T128[4'ha:4'ha];
  assign T248 = T128[4'hb:4'hb];
  assign T249 = T128[4'hc:4'hc];
  assign T250 = T128[4'hd:4'hd];
  assign T251 = T128[4'he:4'he];
  assign T252 = T128[4'hf:4'hf];
  assign T253 = T128[5'h10:5'h10];
  assign T254 = T128[5'h11:5'h11];
  assign T255 = T128[5'h12:5'h12];
  assign T256 = T128[5'h13:5'h13];
  assign T257 = T128[5'h14:5'h14];
  assign T258 = T128[5'h15:5'h15];
  assign T259 = T128[5'h16:5'h16];
  assign T260 = T128[5'h17:5'h17];
  assign T261 = T128[5'h18:5'h18];
  assign T262 = T128[5'h19:5'h19];
  assign T263 = T128[5'h1a:5'h1a];
  assign T264 = T128[5'h1b:5'h1b];
  assign T265 = T128[5'h1c:5'h1c];
  assign T266 = T128[5'h1d:5'h1d];
  assign T267 = T128[5'h1e:5'h1e];
  assign T268 = T128[5'h1f:5'h1f];
  assign T269 = T128[6'h20:6'h20];
  assign T270 = T128[6'h21:6'h21];
  assign T271 = T128[6'h22:6'h22];
  assign T272 = T128[6'h23:6'h23];
  assign T273 = T128[6'h24:6'h24];
  assign T274 = T128[6'h25:6'h25];
  assign T275 = T128[6'h26:6'h26];
  assign T276 = T128[6'h27:6'h27];
  assign T277 = T128[6'h28:6'h28];
  assign T278 = T128[6'h29:6'h29];
  assign T279 = T128[6'h2a:6'h2a];
  assign T280 = T128[6'h2b:6'h2b];
  assign T281 = T128[6'h2c:6'h2c];
  assign T282 = T128[6'h2d:6'h2d];
  assign T283 = T128[6'h2e:6'h2e];
  assign T284 = T128[6'h2f:6'h2f];
  assign T285 = T128[6'h30:6'h30];
  assign T286 = T128[6'h31:6'h31];
  assign T287 = T128[6'h32:6'h32];
  assign T288 = T128[6'h33:6'h33];
  assign T289 = T128[6'h34:6'h34];
  assign T290 = T128[6'h35:6'h35];
  assign T291 = T128[6'h36:6'h36];
  assign T292 = T128[6'h37:6'h37];
  assign T293 = T128[6'h38:6'h38];
  assign T294 = T128[6'h39:6'h39];
  assign T295 = T128[6'h3a:6'h3a];
  assign T296 = T128[6'h3b:6'h3b];
  assign T297 = T128[6'h3c:6'h3c];
  assign T298 = T128[6'h3d:6'h3d];
  assign T299 = T128[6'h3e:6'h3e];
  assign T300 = T128[6'h3f:6'h3f];
  assign T301 = T128[7'h40:7'h40];
  assign T302 = T128[7'h41:7'h41];
  assign T303 = T128[7'h42:7'h42];
  assign T304 = T128[7'h43:7'h43];
  assign T305 = T128[7'h44:7'h44];
  assign T306 = T128[7'h45:7'h45];
  assign T307 = T128[7'h46:7'h46];
  assign T308 = T128[7'h47:7'h47];
  assign T309 = T128[7'h48:7'h48];
  assign T310 = T128[7'h49:7'h49];
  assign T311 = T128[7'h4a:7'h4a];
  assign T312 = T128[7'h4b:7'h4b];
  assign T313 = T128[7'h4c:7'h4c];
  assign T314 = T128[7'h4d:7'h4d];
  assign T315 = T128[7'h4e:7'h4e];
  assign T316 = T128[7'h4f:7'h4f];
  assign T317 = T128[7'h50:7'h50];
  assign T318 = T128[7'h51:7'h51];
  assign T319 = T128[7'h52:7'h52];
  assign T320 = T128[7'h53:7'h53];
  assign T321 = T128[7'h54:7'h54];
  assign T322 = T128[7'h55:7'h55];
  assign T323 = T128[7'h56:7'h56];
  assign T324 = T128[7'h57:7'h57];
  assign T325 = T128[7'h58:7'h58];
  assign T326 = T128[7'h59:7'h59];
  assign T327 = T128[7'h5a:7'h5a];
  assign T328 = T128[7'h5b:7'h5b];
  assign T329 = T128[7'h5c:7'h5c];
  assign T330 = T128[7'h5d:7'h5d];
  assign T331 = T128[7'h5e:7'h5e];
  assign T332 = T128[7'h5f:7'h5f];
  assign T333 = T128[7'h60:7'h60];
  assign T334 = T128[7'h61:7'h61];
  assign T335 = T128[7'h62:7'h62];
  assign T336 = T128[7'h63:7'h63];
  assign T337 = T128[7'h64:7'h64];
  assign T338 = T128[7'h65:7'h65];
  assign T339 = T128[7'h66:7'h66];
  assign T340 = T128[7'h67:7'h67];
  assign T341 = T128[7'h68:7'h68];
  assign T342 = T128[7'h69:7'h69];
  assign T343 = T128[7'h6a:7'h6a];
  assign T344 = T128[7'h6b:7'h6b];
  assign notCDom_signSigSum = sigSum[7'h6d:7'h6d];
  assign CDom_estNormDist = T347 ? CAlignDist : T762;
  assign T762 = {2'h0, T345};
  assign T345 = T346[3'h5:1'h0];
  assign T346 = CAlignDist - 8'h1;
  assign T347 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T348;
  assign T348 = T349 == 13'h0;
  assign T349 = sNatCAlignDist[4'hc:1'h0];
  assign isCDominant = T353 & T350;
  assign T350 = CAlignDist_floor | T351;
  assign T351 = T352 < 13'h36;
  assign T352 = sNatCAlignDist[4'hc:1'h0];
  assign T353 = isZeroC ^ 1'h1;
  assign sExpSum = CAlignDist_floor ? T763 : sExpAlignedProd;
  assign T763 = {2'h0, expC};
  assign T354 = T14[1'h0:1'h0];
  assign T355 = {T361, T356};
  assign T356 = {T360, T357};
  assign T357 = T358[1'h1:1'h1];
  assign T358 = T359[2'h3:2'h2];
  assign T359 = T15[2'h3:1'h0];
  assign T360 = T358[1'h0:1'h0];
  assign T361 = {T364, T362};
  assign T362 = T363[1'h1:1'h1];
  assign T363 = T359[1'h1:1'h0];
  assign T364 = T363[1'h0:1'h0];
  assign T365 = T388 | T366;
  assign T366 = T367 & 16'haaaa;
  assign T367 = T368 << 1'h1;
  assign T368 = T369[4'he:1'h0];
  assign T369 = T386 | T370;
  assign T370 = T371 & 16'hcccc;
  assign T371 = T372 << 2'h2;
  assign T372 = T373[4'hd:1'h0];
  assign T373 = T384 | T374;
  assign T374 = T375 & 16'hf0f0;
  assign T375 = T376 << 3'h4;
  assign T376 = T377[4'hb:1'h0];
  assign T377 = T382 | T378;
  assign T378 = T379 & 16'hff00;
  assign T379 = T380 << 4'h8;
  assign T380 = T381[3'h7:1'h0];
  assign T381 = T16[4'hf:1'h0];
  assign T382 = T764 & 16'hff;
  assign T764 = {8'h0, T383};
  assign T383 = T381 >> 4'h8;
  assign T384 = T765 & 16'hf0f;
  assign T765 = {4'h0, T385};
  assign T385 = T377 >> 3'h4;
  assign T386 = T766 & 16'h3333;
  assign T766 = {2'h0, T387};
  assign T387 = T373 >> 2'h2;
  assign T388 = T767 & 16'h5555;
  assign T767 = {1'h0, T389};
  assign T389 = T369 >> 1'h1;
  assign T390 = T419 | T391;
  assign T391 = T392 & 32'haaaaaaaa;
  assign T392 = T393 << 1'h1;
  assign T393 = T394[5'h1e:1'h0];
  assign T394 = T417 | T395;
  assign T395 = T396 & 32'hcccccccc;
  assign T396 = T397 << 2'h2;
  assign T397 = T398[5'h1d:1'h0];
  assign T398 = T415 | T399;
  assign T399 = T400 & 32'hf0f0f0f0;
  assign T400 = T401 << 3'h4;
  assign T401 = T402[5'h1b:1'h0];
  assign T402 = T413 | T403;
  assign T403 = T404 & 32'hff00ff00;
  assign T404 = T405 << 4'h8;
  assign T405 = T406[5'h17:1'h0];
  assign T406 = T411 | T407;
  assign T407 = T408 & 32'hffff0000;
  assign T408 = T409 << 5'h10;
  assign T409 = T410[4'hf:1'h0];
  assign T410 = T17[5'h1f:1'h0];
  assign T411 = T768 & 32'hffff;
  assign T768 = {16'h0, T412};
  assign T412 = T410 >> 5'h10;
  assign T413 = T769 & 32'hff00ff;
  assign T769 = {8'h0, T414};
  assign T414 = T406 >> 4'h8;
  assign T415 = T770 & 32'hf0f0f0f;
  assign T770 = {4'h0, T416};
  assign T416 = T402 >> 3'h4;
  assign T417 = T771 & 32'h33333333;
  assign T771 = {2'h0, T418};
  assign T418 = T398 >> 2'h2;
  assign T419 = T772 & 32'h55555555;
  assign T772 = {1'h0, T420};
  assign T420 = T394 >> 1'h1;
  assign T421 = 56'h0 - T773;
  assign T773 = {55'h0, T422};
  assign T422 = sExpX3[4'hd:4'hd];
  assign sigX3 = T423[6'h38:1'h0];
  assign T423 = {T595, T424};
  assign T424 = doIncrSig ? T591 : T425;
  assign T425 = T426 != 32'h0;
  assign T426 = T496 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T427, 1'h1};
  assign T427 = {T471, T428};
  assign T428 = {T452, T429};
  assign T429 = {T442, T430};
  assign T430 = {T438, T431};
  assign T431 = T432[2'h2:2'h2];
  assign T432 = T433[3'h6:3'h4];
  assign T433 = T434[4'he:4'h8];
  assign T434 = T435[5'h1e:5'h10];
  assign T435 = T436[5'h1f:1'h1];
  assign T436 = $signed(33'h100000000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T437;
  assign T437 = estNormDist[3'h4:1'h0];
  assign T438 = {T441, T439};
  assign T439 = T440[1'h1:1'h1];
  assign T440 = T432[1'h1:1'h0];
  assign T441 = T440[1'h0:1'h0];
  assign T442 = {T448, T443};
  assign T443 = {T447, T444};
  assign T444 = T445[1'h1:1'h1];
  assign T445 = T446[2'h3:2'h2];
  assign T446 = T433[2'h3:1'h0];
  assign T447 = T445[1'h0:1'h0];
  assign T448 = {T451, T449};
  assign T449 = T450[1'h1:1'h1];
  assign T450 = T446[1'h1:1'h0];
  assign T451 = T450[1'h0:1'h0];
  assign T452 = T469 | T453;
  assign T453 = T454 & 8'haa;
  assign T454 = T455 << 1'h1;
  assign T455 = T456[3'h6:1'h0];
  assign T456 = T467 | T457;
  assign T457 = T458 & 8'hcc;
  assign T458 = T459 << 2'h2;
  assign T459 = T460[3'h5:1'h0];
  assign T460 = T465 | T461;
  assign T461 = T462 & 8'hf0;
  assign T462 = T463 << 3'h4;
  assign T463 = T464[2'h3:1'h0];
  assign T464 = T434[3'h7:1'h0];
  assign T465 = T774 & 8'hf;
  assign T774 = {4'h0, T466};
  assign T466 = T464 >> 3'h4;
  assign T467 = T775 & 8'h33;
  assign T775 = {2'h0, T468};
  assign T468 = T460 >> 2'h2;
  assign T469 = T776 & 8'h55;
  assign T776 = {1'h0, T470};
  assign T470 = T456 >> 1'h1;
  assign T471 = T494 | T472;
  assign T472 = T473 & 16'haaaa;
  assign T473 = T474 << 1'h1;
  assign T474 = T475[4'he:1'h0];
  assign T475 = T492 | T476;
  assign T476 = T477 & 16'hcccc;
  assign T477 = T478 << 2'h2;
  assign T478 = T479[4'hd:1'h0];
  assign T479 = T490 | T480;
  assign T480 = T481 & 16'hf0f0;
  assign T481 = T482 << 3'h4;
  assign T482 = T483[4'hb:1'h0];
  assign T483 = T488 | T484;
  assign T484 = T485 & 16'hff00;
  assign T485 = T486 << 4'h8;
  assign T486 = T487[3'h7:1'h0];
  assign T487 = T435[4'hf:1'h0];
  assign T488 = T777 & 16'hff;
  assign T777 = {8'h0, T489};
  assign T489 = T487 >> 4'h8;
  assign T490 = T778 & 16'hf0f;
  assign T778 = {4'h0, T491};
  assign T491 = T483 >> 3'h4;
  assign T492 = T779 & 16'h3333;
  assign T779 = {2'h0, T493};
  assign T493 = T479 >> 2'h2;
  assign T494 = T780 & 16'h5555;
  assign T780 = {1'h0, T495};
  assign T495 = T475 >> 1'h1;
  assign T496 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T570 : T781;
  assign T781 = {1'h0, T497};
  assign T497 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T534 ? T522 : T498;
  assign T498 = T521 ? T502 : T499;
  assign T499 = {T501, T500};
  assign T500 = 54'h0 - T782;
  assign T782 = {53'h0, doSubMags};
  assign T501 = sigSum[6'h21:1'h1];
  assign T502 = T520 ? T784 : T503;
  assign T503 = {T505, T504};
  assign T504 = 86'h0 - T783;
  assign T783 = {85'h0, doSubMags};
  assign T505 = sigSum[1'h1:1'h1];
  assign T784 = {21'h0, T506};
  assign T506 = {T519, T507};
  assign T507 = doSubMags ? T513 : T508;
  assign T508 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T511, T509};
  assign T509 = T510 != 44'h0;
  assign T510 = sigSum[6'h2b:1'h0];
  assign T511 = T512 != 32'h0;
  assign T512 = sigSum[7'h4b:6'h2c];
  assign T513 = ~ T514;
  assign T514 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T517, T515};
  assign T515 = T516 != 44'h0;
  assign T516 = notSigSum[6'h2b:1'h0];
  assign notSigSum = ~ sigSum;
  assign T517 = T518 != 32'h0;
  assign T518 = notSigSum[7'h4b:6'h2c];
  assign T519 = sigSum[7'h6c:6'h2c];
  assign T520 = estNormNeg_dist[3'h4:3'h4];
  assign T521 = estNormNeg_dist[3'h5:3'h5];
  assign T522 = T533 ? T530 : T523;
  assign T523 = {T529, T524};
  assign T524 = doSubMags ? T527 : T525;
  assign T525 = T526 != 11'h0;
  assign T526 = sigSum[4'hb:1'h1];
  assign T527 = T528 == 11'h0;
  assign T528 = notSigSum[4'hb:1'h1];
  assign T529 = sigSum[7'h61:4'hc];
  assign T530 = {T532, T531};
  assign T531 = 22'h0 - T785;
  assign T785 = {21'h0, doSubMags};
  assign T532 = sigSum[7'h41:1'h1];
  assign T533 = estNormNeg_dist[3'h5:3'h5];
  assign T534 = estNormNeg_dist[3'h6:3'h6];
  assign CDom_firstNormAbsSigSum = T535;
  assign T535 = T543 | T536;
  assign T536 = T786 & T537;
  assign T537 = {T539, T538};
  assign T538 = firstReduceNotSigSum[1'h0:1'h0];
  assign T539 = notSigSum[8'h81:6'h2c];
  assign T786 = T540 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T540 = T541;
  assign T541 = doSubMags & T542;
  assign T542 = CDom_estNormDist[3'h5:3'h5];
  assign T543 = T552 | T544;
  assign T544 = T787 & T545;
  assign T545 = {T547, T546};
  assign T546 = firstReduceNotSigSum != 2'h0;
  assign T547 = notSigSum[8'ha1:7'h4c];
  assign T787 = T548 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T548 = T549;
  assign T549 = doSubMags & T550;
  assign T550 = ~ T551;
  assign T551 = CDom_estNormDist[3'h5:3'h5];
  assign T552 = T561 | T553;
  assign T553 = T788 & T554;
  assign T554 = {T556, T555};
  assign T555 = firstReduceSigSum[1'h0:1'h0];
  assign T556 = sigSum[8'h81:6'h2c];
  assign T788 = T557 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T557 = T558;
  assign T558 = T560 & T559;
  assign T559 = CDom_estNormDist[3'h5:3'h5];
  assign T560 = ~ doSubMags;
  assign T561 = T789 & T562;
  assign T562 = {T564, T563};
  assign T563 = firstReduceSigSum != 2'h0;
  assign T564 = sigSum[8'ha1:7'h4c];
  assign T789 = T565 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T565 = T566;
  assign T566 = T569 & T567;
  assign T567 = ~ T568;
  assign T568 = CDom_estNormDist[3'h5:3'h5];
  assign T569 = ~ doSubMags;
  assign T570 = isCDominant ? T791 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T590 ? T582 : T571;
  assign T571 = T581 ? T574 : T572;
  assign T572 = T573 << 6'h36;
  assign T573 = notSigSum[6'h22:1'h1];
  assign T574 = T580 ? T790 : T575;
  assign T575 = T576 << 7'h56;
  assign T576 = notSigSum[2'h2:1'h1];
  assign T790 = {23'h0, T577};
  assign T577 = {T579, T578};
  assign T578 = firstReduceNotSigSum[1'h0:1'h0];
  assign T579 = notSigSum[7'h6b:6'h2c];
  assign T580 = estNormNeg_dist[3'h4:3'h4];
  assign T581 = estNormNeg_dist[3'h5:3'h5];
  assign T582 = T589 ? T587 : T583;
  assign T583 = {T586, T584};
  assign T584 = T585 != 11'h0;
  assign T585 = notSigSum[4'hb:1'h1];
  assign T586 = notSigSum[7'h62:4'hc];
  assign T587 = T588 << 5'h16;
  assign T588 = notSigSum[7'h42:1'h1];
  assign T589 = estNormNeg_dist[3'h5:3'h5];
  assign T590 = estNormNeg_dist[3'h6:3'h6];
  assign T791 = {1'h0, CDom_firstNormAbsSigSum};
  assign T591 = T592 == 32'h0;
  assign T592 = T593 & absSigSumExtraMask;
  assign T593 = ~ T594;
  assign T594 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign T595 = T596 >> normTo2ShiftDist;
  assign T596 = cFirstNormAbsSigSum[7'h57:1'h1];
  assign roundPosBit = T597 != 57'h0;
  assign T597 = sigX3 & T792;
  assign T792 = {1'h0, roundPosMask};
  assign roundPosMask = T793 & roundMask;
  assign T793 = {1'h0, T598};
  assign T598 = ~ T599;
  assign T599 = roundMask >> 1'h1;
  assign T600 = ~ allRound;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T601 == 57'h0;
  assign T601 = T603 & T794;
  assign T794 = {2'h0, T602};
  assign T602 = roundMask >> 1'h1;
  assign T603 = ~ sigX3;
  assign doIncrSig = T604 & doSubMags;
  assign T604 = T606 & T605;
  assign T605 = ~ notCDom_signSigSum;
  assign T606 = ~ isCDominant;
  assign commonCase = T608 & T607;
  assign T607 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T608 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T609 == 2'h3;
  assign T609 = expC[4'hb:4'ha];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T610 == 2'h3;
  assign T610 = expB[4'hb:4'ha];
  assign isSpecialA = T611 == 2'h3;
  assign T611 = expA[4'hb:4'ha];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T612;
  assign T612 = T616 | T613;
  assign T613 = sExpX3_13 <= T795;
  assign T795 = {2'h0, T614};
  assign T614 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign sigX3Shift1 = T615 == 2'h0;
  assign T615 = sigX3[6'h38:6'h37];
  assign T616 = sExpX3[4'hd:4'hd];
  assign overflow = commonCase & overflowY;
  assign overflowY = T617 == 3'h3;
  assign T617 = sExpY[4'hc:4'ha];
  assign sExpY = T664 | T618;
  assign T618 = T620 ? T619 : 14'h0;
  assign T619 = sExpX3 - 14'h1;
  assign T620 = T621 == 2'h0;
  assign T621 = sigY3[6'h36:6'h35];
  assign sigY3 = T635 | T622;
  assign T622 = roundEven ? T623 : 55'h0;
  assign T623 = roundUp_sigY3 & T624;
  assign T624 = ~ T625;
  assign T625 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T626[6'h36:1'h0];
  assign T626 = T627 + 55'h1;
  assign T627 = T628 >> 2'h2;
  assign T628 = sigX3 | T796;
  assign T796 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T632 : T629;
  assign T629 = T631 & T630;
  assign T630 = ~ anyRoundExtra;
  assign T631 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T632 = T633 & allRoundExtra;
  assign T633 = roundingMode_nearest_even & T634;
  assign T634 = ~ roundPosBit;
  assign T635 = T657 | T636;
  assign T636 = roundUp ? roundUp_sigY3 : 55'h0;
  assign roundUp = T644 | T637;
  assign T637 = T638 & 1'h1;
  assign T638 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T642 & T639;
  assign T639 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T640 : notCDom_signSigSum;
  assign T640 = doSubMags & T641;
  assign T641 = ~ isZeroC;
  assign T642 = ~ isZeroY;
  assign isZeroY = T643 == 3'h0;
  assign T643 = sigX3[6'h38:6'h36];
  assign T644 = T647 | T645;
  assign T645 = T646 & roundPosBit;
  assign T646 = doIncrSig & roundingMode_nearest_even;
  assign T647 = T649 | T648;
  assign T648 = doIncrSig & allRound;
  assign T649 = T653 | T650;
  assign T650 = T651 & anyRound;
  assign T651 = T652 & roundDirectUp;
  assign T652 = ~ doIncrSig;
  assign T653 = T654 & anyRoundExtra;
  assign T654 = T655 & roundPosBit;
  assign T655 = T656 & roundingMode_nearest_even;
  assign T656 = ~ doIncrSig;
  assign T657 = T661 ? T658 : 55'h0;
  assign T658 = T659 >> 2'h2;
  assign T659 = sigX3 & T797;
  assign T797 = {1'h0, T660};
  assign T660 = ~ roundMask;
  assign T661 = T663 & T662;
  assign T662 = ~ roundEven;
  assign T663 = ~ roundUp;
  assign T664 = T667 | T665;
  assign T665 = T666 ? sExpX3 : 14'h0;
  assign T666 = sigY3[6'h35:6'h35];
  assign T667 = T669 ? T668 : 14'h0;
  assign T668 = sExpX3 + 14'h1;
  assign T669 = sigY3[6'h36:6'h36];
  assign T670 = {invalid, 1'h0};
  assign invalid = T689 | notSigNaN_invalid;
  assign notSigNaN_invalid = T686 | T671;
  assign T671 = T672 & doSubMags;
  assign T672 = T675 & isInfC;
  assign isInfC = isSpecialC & T673;
  assign T673 = T674 ^ 1'h1;
  assign T674 = expC[4'h9:4'h9];
  assign T675 = T681 & T676;
  assign T676 = isInfA | isInfB;
  assign isInfB = isSpecialB & T677;
  assign T677 = T678 ^ 1'h1;
  assign T678 = expB[4'h9:4'h9];
  assign isInfA = isSpecialA & T679;
  assign T679 = T680 ^ 1'h1;
  assign T680 = expA[4'h9:4'h9];
  assign T681 = T684 & T682;
  assign T682 = ~ isNaNB;
  assign isNaNB = isSpecialB & T683;
  assign T683 = expB[4'h9:4'h9];
  assign T684 = ~ isNaNA;
  assign isNaNA = isSpecialA & T685;
  assign T685 = expA[4'h9:4'h9];
  assign T686 = T688 | T687;
  assign T687 = isZeroA & isInfB;
  assign T688 = isInfA & isZeroB;
  assign T689 = T693 | isSigNaNC;
  assign isSigNaNC = isNaNC & T690;
  assign T690 = T691 ^ 1'h1;
  assign T691 = fractC[6'h33:6'h33];
  assign isNaNC = isSpecialC & T692;
  assign T692 = expC[4'h9:4'h9];
  assign T693 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T694;
  assign T694 = T695 ^ 1'h1;
  assign T695 = fractB[6'h33:6'h33];
  assign isSigNaNA = isNaNA & T696;
  assign T696 = T697 ^ 1'h1;
  assign T697 = fractA[6'h33:6'h33];
  assign io_out = T698;
  assign T698 = {signOut, T699};
  assign T699 = {expOut, fractOut};
  assign fractOut = fractY | T700;
  assign T700 = 52'h0 - T798;
  assign T798 = {51'h0, T701};
  assign T701 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T702;
  assign T702 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T705 | T703;
  assign T703 = roundingMode_max & T704;
  assign T704 = ~ signY;
  assign T705 = roundingMode_nearest_even | T706;
  assign T706 = roundingMode_min & signY;
  assign isNaNOut = T707 | notSigNaN_invalid;
  assign T707 = T708 | isNaNC;
  assign T708 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T710 : T709;
  assign T709 = sigY3[6'h34:1'h1];
  assign T710 = sigY3[6'h33:1'h0];
  assign expOut = T712 | T711;
  assign T711 = isNaNOut ? 12'he00 : 12'h0;
  assign T712 = T717 | T713;
  assign T713 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = T715 | T714;
  assign T714 = overflow & overflowY_roundMagUp;
  assign T715 = T716 | isInfC;
  assign T716 = isInfA | isInfB;
  assign T717 = T719 | T718;
  assign T718 = isSatOut ? 12'hbff : 12'h0;
  assign T719 = T722 & T720;
  assign T720 = ~ T721;
  assign T721 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T722 = T725 & T723;
  assign T723 = ~ T724;
  assign T724 = isSatOut ? 12'h400 : 12'h0;
  assign T725 = expY & T726;
  assign T726 = ~ T727;
  assign T727 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign notSpecial_isZeroOut = T731 | totalUnderflowY;
  assign totalUnderflowY = T730 | T728;
  assign T728 = T729 < 12'h3ce;
  assign T729 = sExpY[4'hb:1'h0];
  assign T730 = sExpY[4'hc:4'hc];
  assign T731 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'hb:1'h0];
  assign signOut = T733 | T732;
  assign T732 = commonCase & signY;
  assign T733 = T737 | T734;
  assign T734 = T735 & opSignC;
  assign T735 = T736 & isSpecialC;
  assign T736 = mulSpecial ^ 1'h1;
  assign T737 = T741 | T738;
  assign T738 = T739 & signProd;
  assign T739 = mulSpecial & T740;
  assign T740 = isSpecialC ^ 1'h1;
  assign T741 = T742 | isNaNOut;
  assign T742 = T743 & opSignC;
  assign T743 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_1(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T12;
  reg [2:0] in_rm;
  wire[2:0] T13;
  reg [64:0] in_in3;
  wire[64:0] T14;
  wire[64:0] T15;
  wire[64:0] zero;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg [64:0] in_in2;
  wire[64:0] T22;
  wire[64:0] T23;
  wire T24;
  reg [64:0] in_in1;
  wire[64:0] T25;
  wire[1:0] T26;
  reg [4:0] in_cmd;
  wire[4:0] T27;
  wire[4:0] T28;
  wire[4:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg [4:0] R0;
  wire[4:0] T1;
  reg [4:0] R2;
  wire[4:0] T3;
  wire[4:0] res_exc;
  reg  valid;
  reg  R4;
  wire T10;
  reg [64:0] R5;
  wire[64:0] T6;
  reg [64:0] R7;
  wire[64:0] T8;
  wire[64:0] res_data;
  reg  R9;
  wire T11;
  wire[64:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R0 = {1{$random}};
    R2 = {1{$random}};
    valid = {1{$random}};
    R4 = {1{$random}};
    R5 = {3{$random}};
    R7 = {3{$random}};
    R9 = {1{$random}};
  end
`endif

  assign T12 = in_rm[1'h1:1'h0];
  assign T13 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T14 = T19 ? zero : T15;
  assign T15 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign zero = T16 << 7'h40;
  assign T16 = T18 ^ T17;
  assign T17 = io_in_bits_in2[7'h40:7'h40];
  assign T18 = io_in_bits_in1[7'h40:7'h40];
  assign T19 = io_in_valid & T20;
  assign T20 = T21 ^ 1'h1;
  assign T21 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T22 = T24 ? 65'h8000000000000000 : T23;
  assign T23 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T24 = io_in_valid & io_in_bits_swap23;
  assign T25 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T26 = in_cmd[1'h1:1'h0];
  assign T27 = io_in_valid ? T29 : T28;
  assign T28 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T29 = {3'h0, T30};
  assign T30 = {T32, T31};
  assign T31 = io_in_bits_cmd[1'h0:1'h0];
  assign T32 = T34 & T33;
  assign T33 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T34 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R0;
  assign T1 = R4 ? R2 : R0;
  assign T3 = valid ? res_exc : R2;
  assign res_exc = fma_io_exceptionFlags;
  assign T10 = reset ? 1'h0 : valid;
  assign io_out_bits_data = R5;
  assign T6 = R4 ? R7 : R5;
  assign T8 = valid ? res_data : R7;
  assign res_data = fma_io_out;
  assign io_out_valid = R9;
  assign T11 = reset ? 1'h0 : R4;
  mulAddSubRecodedFloatN_1 fma(
       .io_op( T26 ),
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_c( in_in3 ),
       .io_roundingMode( T12 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T19) begin
      in_in3 <= zero;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T24) begin
      in_in2 <= 65'h8000000000000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T29;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(R4) begin
      R0 <= R2;
    end
    if(valid) begin
      R2 <= res_exc;
    end
    valid <= io_in_valid;
    if(reset) begin
      R4 <= 1'h0;
    end else begin
      R4 <= valid;
    end
    if(R4) begin
      R5 <= R7;
    end
    if(valid) begin
      R7 <= res_data;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else begin
      R9 <= R4;
    end
  end
endmodule

module recodedFloatNCompare(
    input [64:0] io_a,
    input [64:0] io_b,
    output io_a_eq_b,
    output io_a_lt_b,
    output io_a_eq_b_invalid,
    output io_a_lt_b_invalid
);

  wire T0;
  wire isNaNB;
  wire[2:0] codeB;
  wire[11:0] expB;
  wire isNaNA;
  wire[2:0] codeA;
  wire[11:0] expA;
  wire T1;
  wire isSignalingNaNB;
  wire T2;
  wire T3;
  wire[51:0] sigB;
  wire isSignalingNaNA;
  wire T4;
  wire T5;
  wire[51:0] sigA;
  wire T6;
  wire T7;
  wire T8;
  wire magLess;
  wire T9;
  wire T10;
  wire expEqual;
  wire T11;
  wire T12;
  wire T13;
  wire isZeroB;
  wire T14;
  wire isZeroA;
  wire T15;
  wire signA;
  wire T16;
  wire T17;
  wire magEqual;
  wire T18;
  wire T19;
  wire T20;
  wire signB;
  wire T21;
  wire T22;
  wire T23;
  wire signEqual;
  wire T24;
  wire T25;


  assign io_a_lt_b_invalid = T0;
  assign T0 = isNaNA | isNaNB;
  assign isNaNB = codeB == 3'h7;
  assign codeB = expB[4'hb:4'h9];
  assign expB = io_b[6'h3f:6'h34];
  assign isNaNA = codeA == 3'h7;
  assign codeA = expA[4'hb:4'h9];
  assign expA = io_a[6'h3f:6'h34];
  assign io_a_eq_b_invalid = T1;
  assign T1 = isSignalingNaNA | isSignalingNaNB;
  assign isSignalingNaNB = isNaNB & T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = sigB[6'h33:6'h33];
  assign sigB = io_b[6'h33:1'h0];
  assign isSignalingNaNA = isNaNA & T4;
  assign T4 = T5 ^ 1'h1;
  assign T5 = sigA[6'h33:6'h33];
  assign sigA = io_a[6'h33:1'h0];
  assign io_a_lt_b = T6;
  assign T6 = T21 & T7;
  assign T7 = signB ? T16 : T8;
  assign T8 = signA ? T12 : magLess;
  assign magLess = T11 | T9;
  assign T9 = expEqual & T10;
  assign T10 = sigA < sigB;
  assign expEqual = expA == expB;
  assign T11 = expA < expB;
  assign T12 = T13 ^ 1'h1;
  assign T13 = isZeroA & isZeroB;
  assign isZeroB = T14 ^ 1'h1;
  assign T14 = codeB != 3'h0;
  assign isZeroA = T15 ^ 1'h1;
  assign T15 = codeA != 3'h0;
  assign signA = io_a[7'h40:7'h40];
  assign T16 = T19 & T17;
  assign T17 = magEqual ^ 1'h1;
  assign magEqual = expEqual & T18;
  assign T18 = sigA == sigB;
  assign T19 = signA & T20;
  assign T20 = magLess ^ 1'h1;
  assign signB = io_b[7'h40:7'h40];
  assign T21 = io_a_lt_b_invalid ^ 1'h1;
  assign io_a_eq_b = T22;
  assign T22 = T24 & T23;
  assign T23 = isZeroA | signEqual;
  assign signEqual = signA == signB;
  assign T24 = T25 & magEqual;
  assign T25 = isNaNA ^ 1'h1;
endmodule

module FPToInt(input clk,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output io_out_bits_lt,
    output[63:0] io_out_bits_store,
    output[63:0] io_out_bits_toint,
    output[4:0] io_out_bits_exc
);

  reg [64:0] in_in2;
  wire[64:0] T346;
  wire[64:0] T347;
  wire[64:0] T348;
  wire[63:0] T349;
  wire[51:0] T350;
  wire[51:0] T351;
  wire[22:0] T352;
  wire[51:0] T353;
  wire[51:0] T354;
  wire T355;
  wire[2:0] T356;
  wire[11:0] T357;
  wire[11:0] T358;
  wire[11:0] T359;
  wire[11:0] T360;
  wire T361;
  wire[11:0] T362;
  wire[7:0] T363;
  wire T364;
  wire[11:0] T365;
  wire[10:0] T366;
  wire T367;
  wire[11:0] T368;
  wire T369;
  wire T370;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[4:0] T49;
  wire T50;
  wire T51;
  reg [64:0] in_in1;
  wire[64:0] T23;
  wire[64:0] T24;
  wire[64:0] T25;
  wire[63:0] T26;
  wire[51:0] T27;
  wire[51:0] T28;
  wire[22:0] T29;
  wire[51:0] T30;
  wire[51:0] T331;
  wire T31;
  wire[2:0] T32;
  wire[11:0] T33;
  wire[11:0] T34;
  wire[11:0] T35;
  wire[11:0] T36;
  wire T37;
  wire[11:0] T38;
  wire[7:0] T42;
  wire T39;
  wire[11:0] T332;
  wire[10:0] T40;
  wire T41;
  wire[11:0] T333;
  wire T43;
  wire T44;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] dcmp_exc;
  wire T2;
  wire[2:0] T3;
  wire[2:0] T330;
  wire[1:0] T4;
  wire[2:0] T5;
  reg [2:0] in_rm;
  wire[2:0] T6;
  wire T7;
  wire[4:0] T8;
  reg [4:0] in_cmd;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[3:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] T15;
  wire[2:0] T16;
  wire T17;
  wire[50:0] T18;
  wire[115:0] T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire[11:0] T22;
  wire T52;
  wire T53;
  wire[52:0] T54;
  wire[51:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[10:0] T66;
  wire T67;
  wire T68;
  wire[63:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[1:0] T87;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[10:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[1:0] T110;
  reg [1:0] in_typ;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[1:0] T127;
  wire T128;
  wire[4:0] T129;
  wire[63:0] T130;
  wire[63:0] T131;
  wire[63:0] T132;
  wire[63:0] unrec_out;
  wire[63:0] unrec_d;
  wire[62:0] T133;
  wire[51:0] T134;
  wire[51:0] T135;
  wire[51:0] T136;
  wire[52:0] T137;
  wire[5:0] T138;
  wire[5:0] T139;
  wire[11:0] T140;
  wire[52:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[9:0] T145;
  wire T146;
  wire[1:0] T147;
  wire T148;
  wire[2:0] T149;
  wire[51:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire[1:0] T162;
  wire[10:0] T163;
  wire[10:0] T164;
  wire[10:0] T334;
  wire[10:0] T165;
  wire[10:0] T166;
  wire T167;
  wire[63:0] T168;
  wire[31:0] unrec_s;
  wire[30:0] T169;
  wire[22:0] T170;
  wire[22:0] T171;
  wire[22:0] T172;
  wire[23:0] T173;
  wire[4:0] T174;
  wire[4:0] T175;
  wire[8:0] T176;
  wire[23:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire[6:0] T181;
  wire T182;
  wire[1:0] T183;
  wire T184;
  wire[2:0] T185;
  wire[22:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[1:0] T191;
  wire T192;
  wire T193;
  wire[1:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire[1:0] T198;
  wire[7:0] T199;
  wire[7:0] T200;
  wire[7:0] T335;
  wire[7:0] T201;
  wire[7:0] T202;
  wire T203;
  wire[31:0] T204;
  wire[31:0] T336;
  wire T205;
  reg  in_single;
  wire T206;
  wire[63:0] T337;
  wire[9:0] classify_out;
  wire[9:0] classify_d;
  wire[4:0] T207;
  wire[2:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[11:0] T215;
  wire T216;
  wire[1:0] T217;
  wire[2:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[9:0] T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[4:0] T237;
  wire[2:0] T238;
  wire[1:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire[1:0] T246;
  wire T247;
  wire T248;
  wire T249;
  wire[51:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire[9:0] classify_s;
  wire[4:0] T254;
  wire[2:0] T255;
  wire[1:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire[8:0] T262;
  wire T263;
  wire[1:0] T264;
  wire[2:0] T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire[6:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[1:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[4:0] T284;
  wire[2:0] T285;
  wire[1:0] T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[22:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire[63:0] T338;
  wire dcmp_out;
  wire[2:0] T302;
  wire[2:0] T339;
  wire[1:0] T303;
  wire[2:0] T304;
  wire[63:0] T305;
  wire[63:0] T340;
  wire[31:0] T306;
  wire[31:0] T307;
  wire[31:0] T341;
  wire T342;
  wire[63:0] T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] T312;
  wire[63:0] T313;
  wire T314;
  wire[63:0] T315;
  wire[63:0] T316;
  wire[63:0] T317;
  wire[63:0] T343;
  wire[31:0] T318;
  wire T319;
  wire T320;
  wire T321;
  wire[31:0] T344;
  wire T345;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg  valid;
  wire dcmp_io_a_eq_b;
  wire dcmp_io_a_lt_b;
  wire dcmp_io_a_eq_b_invalid;
  wire dcmp_io_a_lt_b_invalid;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_rm = {1{$random}};
    in_cmd = {1{$random}};
    in_typ = {1{$random}};
    in_single = {1{$random}};
    valid = {1{$random}};
  end
`endif

  assign T346 = T45 ? T348 : T347;
  assign T347 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T348 = {T370, T349};
  assign T349 = {T357, T350};
  assign T350 = T353 | T351;
  assign T351 = T352 << 5'h1d;
  assign T352 = io_in_bits_in2[5'h16:1'h0];
  assign T353 = 52'h0 - T354;
  assign T354 = {51'h0, T355};
  assign T355 = T356 == 3'h7;
  assign T356 = io_in_bits_in2[5'h1f:5'h1d];
  assign T357 = T369 ? T368 : T358;
  assign T358 = T367 ? T365 : T359;
  assign T359 = T364 ? T362 : T360;
  assign T360 = T361 ? 12'hc00 : 12'he00;
  assign T361 = T356 < 3'h7;
  assign T362 = {4'h8, T363};
  assign T363 = io_in_bits_in2[5'h1e:5'h17];
  assign T364 = T356 < 3'h6;
  assign T365 = {1'h0, T366};
  assign T366 = {3'h7, T363};
  assign T367 = T356 < 3'h4;
  assign T368 = {4'h0, T363};
  assign T369 = T356 < 3'h1;
  assign T370 = io_in_bits_in2[6'h20:6'h20];
  assign T45 = io_in_valid & T46;
  assign T46 = T50 & T47;
  assign T47 = T48 == 1'h0;
  assign T48 = T49 == 5'hc;
  assign T49 = io_in_bits_cmd & 5'hc;
  assign T50 = io_in_bits_single & T51;
  assign T51 = io_in_bits_ldst ^ 1'h1;
  assign T23 = T45 ? T25 : T24;
  assign T24 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T25 = {T44, T26};
  assign T26 = {T33, T27};
  assign T27 = T30 | T28;
  assign T28 = T29 << 5'h1d;
  assign T29 = io_in_bits_in1[5'h16:1'h0];
  assign T30 = 52'h0 - T331;
  assign T331 = {51'h0, T31};
  assign T31 = T32 == 3'h7;
  assign T32 = io_in_bits_in1[5'h1f:5'h1d];
  assign T33 = T43 ? T333 : T34;
  assign T34 = T41 ? T332 : T35;
  assign T35 = T39 ? T38 : T36;
  assign T36 = T37 ? 12'hc00 : 12'he00;
  assign T37 = T32 < 3'h7;
  assign T38 = {4'h8, T42};
  assign T42 = io_in_bits_in1[5'h1e:5'h17];
  assign T39 = T32 < 3'h6;
  assign T332 = {1'h0, T40};
  assign T40 = {3'h7, T42};
  assign T41 = T32 < 3'h4;
  assign T333 = {4'h0, T42};
  assign T43 = T32 < 3'h1;
  assign T44 = io_in_bits_in1[6'h20:6'h20];
  assign io_out_bits_exc = T0;
  assign T0 = T128 ? T10 : T1;
  assign T1 = T7 ? dcmp_exc : 5'h0;
  assign dcmp_exc = T2 << 3'h4;
  assign T2 = T3 != 3'h0;
  assign T3 = T5 & T330;
  assign T330 = {1'h0, T4};
  assign T4 = {dcmp_io_a_lt_b_invalid, dcmp_io_a_eq_b_invalid};
  assign T5 = ~ in_rm;
  assign T6 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T7 = T8 == 5'h4;
  assign T8 = in_cmd & 5'hc;
  assign T9 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T10 = {T58, T11};
  assign T11 = {3'h0, T12};
  assign T12 = T14 & T13;
  assign T13 = T58 ^ 1'h1;
  assign T14 = T15 != 2'h0;
  assign T15 = T16[1'h1:1'h0];
  assign T16 = {T57, T17};
  assign T17 = T18 != 51'h0;
  assign T18 = T19[6'h32:1'h0];
  assign T19 = T54 << T20;
  assign T20 = T52 ? 6'h0 : T21;
  assign T21 = T22[3'h5:1'h0];
  assign T22 = in_in1[6'h3f:6'h34];
  assign T52 = T53 ^ 1'h1;
  assign T53 = T22[4'hb:4'hb];
  assign T54 = {T56, T55};
  assign T55 = in_in1[6'h33:1'h0];
  assign T56 = T52 ^ 1'h1;
  assign T57 = T19[6'h34:6'h33];
  assign T58 = T126 | T59;
  assign T59 = T125 ? T119 : T60;
  assign T60 = T118 ? T112 : T61;
  assign T61 = T109 ? T103 : T62;
  assign T62 = T52 ? 1'h0 : T63;
  assign T63 = T102 ? T98 : T64;
  assign T64 = T97 ? T67 : T65;
  assign T65 = 11'h40 <= T66;
  assign T66 = T22[4'ha:1'h0];
  assign T67 = T70 | T68;
  assign T68 = T69 != 64'h0;
  assign T69 = T19[7'h73:6'h34];
  assign T70 = T96 | T71;
  assign T71 = T95 ? T84 : T72;
  assign T72 = T83 ? T82 : T73;
  assign T73 = T81 ? T74 : 1'h0;
  assign T74 = T79 & T75;
  assign T75 = T52 ? T76 : T14;
  assign T76 = T77 ^ 1'h1;
  assign T77 = T78 == 3'h0;
  assign T78 = T22[4'hb:4'h9];
  assign T79 = T80 ^ 1'h1;
  assign T80 = in_in1[7'h40:7'h40];
  assign T81 = in_rm == 3'h3;
  assign T82 = T80 & T75;
  assign T83 = in_rm == 3'h2;
  assign T84 = T52 ? T90 : T85;
  assign T85 = T88 | T86;
  assign T86 = T87 == 2'h3;
  assign T87 = T16[1'h1:1'h0];
  assign T88 = T89 == 2'h3;
  assign T89 = T16[2'h2:1'h1];
  assign T90 = T91 & T14;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T94 == 11'h7ff;
  assign T94 = T22[4'ha:1'h0];
  assign T95 = in_rm == 3'h0;
  assign T96 = T80 ^ 1'h1;
  assign T97 = T66 == 11'h3f;
  assign T98 = T101 & T99;
  assign T99 = T71 & T100;
  assign T100 = T69 == 64'hffffffffffffffff;
  assign T101 = T80 ^ 1'h1;
  assign T102 = T66 == 11'h3e;
  assign T103 = T52 ? T108 : T104;
  assign T104 = T80 | T105;
  assign T105 = T107 ? T99 : T106;
  assign T106 = 11'h40 <= T66;
  assign T107 = T66 == 11'h3f;
  assign T108 = T80 & T71;
  assign T109 = T110 == 2'h2;
  assign T110 = in_typ ^ 2'h1;
  assign T111 = io_in_valid ? io_in_bits_typ : in_typ;
  assign T112 = T52 ? 1'h0 : T113;
  assign T113 = T117 ? T98 : T114;
  assign T114 = T116 ? T67 : T115;
  assign T115 = 11'h20 <= T66;
  assign T116 = T66 == 11'h1f;
  assign T117 = T66 == 11'h1e;
  assign T118 = T110 == 2'h1;
  assign T119 = T52 ? T124 : T120;
  assign T120 = T80 | T121;
  assign T121 = T123 ? T99 : T122;
  assign T122 = 11'h20 <= T66;
  assign T123 = T66 == 11'h1f;
  assign T124 = T80 & T71;
  assign T125 = T110 == 2'h0;
  assign T126 = T127 == 2'h3;
  assign T127 = T22[4'hb:4'ha];
  assign T128 = T129 == 5'h8;
  assign T129 = in_cmd & 5'hc;
  assign io_out_bits_toint = T130;
  assign T130 = T128 ? T305 : T131;
  assign T131 = T7 ? T338 : T132;
  assign T132 = T301 ? T337 : unrec_out;
  assign unrec_out = in_single ? T168 : unrec_d;
  assign unrec_d = {T167, T133};
  assign T133 = {T163, T134};
  assign T134 = T151 ? T150 : T135;
  assign T135 = T142 ? T136 : 52'h0;
  assign T136 = T137[6'h33:1'h0];
  assign T137 = T141 >> T138;
  assign T138 = 6'h2 - T139;
  assign T139 = T140[3'h5:1'h0];
  assign T140 = in_in1[6'h3f:6'h34];
  assign T141 = {1'h1, T150};
  assign T142 = T148 | T143;
  assign T143 = T146 & T144;
  assign T144 = T145 < 10'h2;
  assign T145 = T140[4'h9:1'h0];
  assign T146 = T147 == 2'h1;
  assign T147 = T140[4'hb:4'ha];
  assign T148 = T149 == 3'h1;
  assign T149 = T140[4'hb:4'h9];
  assign T150 = in_in1[6'h33:1'h0];
  assign T151 = T156 | T152;
  assign T152 = T154 & T153;
  assign T153 = T140[4'h9:4'h9];
  assign T154 = T155 == 2'h3;
  assign T155 = T140[4'hb:4'ha];
  assign T156 = T159 | T157;
  assign T157 = T158 == 2'h2;
  assign T158 = T140[4'hb:4'ha];
  assign T159 = T161 & T160;
  assign T160 = T144 ^ 1'h1;
  assign T161 = T162 == 2'h1;
  assign T162 = T140[4'hb:4'ha];
  assign T163 = T156 ? T165 : T164;
  assign T164 = 11'h0 - T334;
  assign T334 = {10'h0, T154};
  assign T165 = T166 - 11'h401;
  assign T166 = T140[4'ha:1'h0];
  assign T167 = in_in1[7'h40:7'h40];
  assign T168 = {T204, unrec_s};
  assign unrec_s = {T203, T169};
  assign T169 = {T199, T170};
  assign T170 = T187 ? T186 : T171;
  assign T171 = T178 ? T172 : 23'h0;
  assign T172 = T173[5'h16:1'h0];
  assign T173 = T177 >> T174;
  assign T174 = 5'h2 - T175;
  assign T175 = T176[3'h4:1'h0];
  assign T176 = in_in1[5'h1f:5'h17];
  assign T177 = {1'h1, T186};
  assign T178 = T184 | T179;
  assign T179 = T182 & T180;
  assign T180 = T181 < 7'h2;
  assign T181 = T176[3'h6:1'h0];
  assign T182 = T183 == 2'h1;
  assign T183 = T176[4'h8:3'h7];
  assign T184 = T185 == 3'h1;
  assign T185 = T176[4'h8:3'h6];
  assign T186 = in_in1[5'h16:1'h0];
  assign T187 = T192 | T188;
  assign T188 = T190 & T189;
  assign T189 = T176[3'h6:3'h6];
  assign T190 = T191 == 2'h3;
  assign T191 = T176[4'h8:3'h7];
  assign T192 = T195 | T193;
  assign T193 = T194 == 2'h2;
  assign T194 = T176[4'h8:3'h7];
  assign T195 = T197 & T196;
  assign T196 = T180 ^ 1'h1;
  assign T197 = T198 == 2'h1;
  assign T198 = T176[4'h8:3'h7];
  assign T199 = T192 ? T201 : T200;
  assign T200 = 8'h0 - T335;
  assign T335 = {7'h0, T190};
  assign T201 = T202 - 8'h81;
  assign T202 = T176[3'h7:1'h0];
  assign T203 = in_in1[6'h20:6'h20];
  assign T204 = 32'h0 - T336;
  assign T336 = {31'h0, T205};
  assign T205 = unrec_s[5'h1f:5'h1f];
  assign T206 = io_in_valid ? io_in_bits_single : in_single;
  assign T337 = {54'h0, classify_out};
  assign classify_out = in_single ? classify_s : classify_d;
  assign classify_d = {T237, T207};
  assign T207 = {T232, T208};
  assign T208 = {T227, T209};
  assign T209 = {T219, T210};
  assign T210 = T212 & T211;
  assign T211 = in_in1[7'h40:7'h40];
  assign T212 = T216 & T213;
  assign T213 = T214 ^ 1'h1;
  assign T214 = T215[4'h9:4'h9];
  assign T215 = in_in1[6'h3f:6'h34];
  assign T216 = T217 == 2'h3;
  assign T217 = T218[2'h2:1'h1];
  assign T218 = T215[4'hb:4'h9];
  assign T219 = T220 & T211;
  assign T220 = T222 | T221;
  assign T221 = T217 == 2'h2;
  assign T222 = T226 & T223;
  assign T223 = T224 ^ 1'h1;
  assign T224 = T225 < 10'h2;
  assign T225 = T215[4'h9:1'h0];
  assign T226 = T217 == 2'h1;
  assign T227 = T228 & T211;
  assign T228 = T231 | T229;
  assign T229 = T230 & T224;
  assign T230 = T217 == 2'h1;
  assign T231 = T218 == 3'h1;
  assign T232 = {T235, T233};
  assign T233 = T234 & T211;
  assign T234 = T218 == 3'h0;
  assign T235 = T234 & T236;
  assign T236 = T211 ^ 1'h1;
  assign T237 = {T246, T238};
  assign T238 = {T244, T239};
  assign T239 = {T242, T240};
  assign T240 = T228 & T241;
  assign T241 = T211 ^ 1'h1;
  assign T242 = T220 & T243;
  assign T243 = T211 ^ 1'h1;
  assign T244 = T212 & T245;
  assign T245 = T211 ^ 1'h1;
  assign T246 = {T252, T247};
  assign T247 = T251 & T248;
  assign T248 = T249 ^ 1'h1;
  assign T249 = T250[6'h33:6'h33];
  assign T250 = in_in1[6'h33:1'h0];
  assign T251 = T218 == 3'h7;
  assign T252 = T251 & T253;
  assign T253 = T250[6'h33:6'h33];
  assign classify_s = {T284, T254};
  assign T254 = {T279, T255};
  assign T255 = {T274, T256};
  assign T256 = {T266, T257};
  assign T257 = T259 & T258;
  assign T258 = in_in1[6'h20:6'h20];
  assign T259 = T263 & T260;
  assign T260 = T261 ^ 1'h1;
  assign T261 = T262[3'h6:3'h6];
  assign T262 = in_in1[5'h1f:5'h17];
  assign T263 = T264 == 2'h3;
  assign T264 = T265[2'h2:1'h1];
  assign T265 = T262[4'h8:3'h6];
  assign T266 = T267 & T258;
  assign T267 = T269 | T268;
  assign T268 = T264 == 2'h2;
  assign T269 = T273 & T270;
  assign T270 = T271 ^ 1'h1;
  assign T271 = T272 < 7'h2;
  assign T272 = T262[3'h6:1'h0];
  assign T273 = T264 == 2'h1;
  assign T274 = T275 & T258;
  assign T275 = T278 | T276;
  assign T276 = T277 & T271;
  assign T277 = T264 == 2'h1;
  assign T278 = T265 == 3'h1;
  assign T279 = {T282, T280};
  assign T280 = T281 & T258;
  assign T281 = T265 == 3'h0;
  assign T282 = T281 & T283;
  assign T283 = T258 ^ 1'h1;
  assign T284 = {T293, T285};
  assign T285 = {T291, T286};
  assign T286 = {T289, T287};
  assign T287 = T275 & T288;
  assign T288 = T258 ^ 1'h1;
  assign T289 = T267 & T290;
  assign T290 = T258 ^ 1'h1;
  assign T291 = T259 & T292;
  assign T292 = T258 ^ 1'h1;
  assign T293 = {T299, T294};
  assign T294 = T298 & T295;
  assign T295 = T296 ^ 1'h1;
  assign T296 = T297[5'h16:5'h16];
  assign T297 = in_in1[5'h16:1'h0];
  assign T298 = T265 == 3'h7;
  assign T299 = T298 & T300;
  assign T300 = T297[5'h16:5'h16];
  assign T301 = in_rm[1'h0:1'h0];
  assign T338 = {63'h0, dcmp_out};
  assign dcmp_out = T302 != 3'h0;
  assign T302 = T304 & T339;
  assign T339 = {1'h0, T303};
  assign T303 = {dcmp_io_a_lt_b, dcmp_io_a_eq_b};
  assign T304 = ~ in_rm;
  assign T305 = T329 ? T308 : T340;
  assign T340 = {T341, T306};
  assign T306 = T307;
  assign T307 = T308[5'h1f:1'h0];
  assign T341 = T342 ? 32'hffffffff : 32'h0;
  assign T342 = T306[5'h1f:5'h1f];
  assign T308 = T58 ? T315 : T309;
  assign T309 = T310;
  assign T310 = T314 ? T313 : T311;
  assign T311 = T80 ? T312 : T69;
  assign T312 = ~ T69;
  assign T313 = T311 + 64'h1;
  assign T314 = T71 ^ T80;
  assign T315 = T327 ? 64'h8000000000000000 : T316;
  assign T316 = T325 ? 64'hffffffff80000000 : T317;
  assign T317 = T322 ? 64'h7fffffffffffffff : T343;
  assign T343 = {T344, T318};
  assign T318 = T319 ? 32'h7fffffff : 32'hffffffff;
  assign T319 = T321 & T320;
  assign T320 = T80 ^ 1'h1;
  assign T321 = T110 == 2'h1;
  assign T344 = T345 ? 32'hffffffff : 32'h0;
  assign T345 = T318[5'h1f:5'h1f];
  assign T322 = T324 & T323;
  assign T323 = T80 ^ 1'h1;
  assign T324 = T110 == 2'h3;
  assign T325 = T326 & T80;
  assign T326 = T110 == 2'h1;
  assign T327 = T328 & T80;
  assign T328 = T110 == 2'h3;
  assign T329 = in_typ[1'h1:1'h1];
  assign io_out_bits_store = unrec_out;
  assign io_out_bits_lt = dcmp_io_a_lt_b;
  assign io_out_valid = valid;
  recodedFloatNCompare dcmp(
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_a_eq_b( dcmp_io_a_eq_b ),
       .io_a_lt_b( dcmp_io_a_lt_b ),
       .io_a_eq_b_invalid( dcmp_io_a_eq_b_invalid ),
       .io_a_lt_b_invalid( dcmp_io_a_lt_b_invalid )
  );

  always @(posedge clk) begin
    if(T45) begin
      in_in2 <= T348;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(T45) begin
      in_in1 <= T25;
    end else if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      in_single <= io_in_bits_single;
    end
    valid <= io_in_valid;
  end
endmodule

module IntToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  reg [4:0] R0;
  wire[4:0] T1;
  reg [4:0] R2;
  wire[4:0] T3;
  wire[4:0] mux_exc;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[1:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[38:0] T12;
  wire[126:0] T13;
  wire[5:0] T14;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[5:0] T216;
  wire[5:0] T217;
  wire[5:0] T218;
  wire[5:0] T219;
  wire[5:0] T220;
  wire[5:0] T221;
  wire[5:0] T222;
  wire[5:0] T223;
  wire[5:0] T224;
  wire[5:0] T225;
  wire[5:0] T226;
  wire[5:0] T227;
  wire[5:0] T228;
  wire[5:0] T229;
  wire[5:0] T230;
  wire[5:0] T231;
  wire[5:0] T232;
  wire[5:0] T233;
  wire[5:0] T234;
  wire[5:0] T235;
  wire[5:0] T236;
  wire[5:0] T237;
  wire[5:0] T238;
  wire[4:0] T239;
  wire[4:0] T240;
  wire[4:0] T241;
  wire[4:0] T242;
  wire[4:0] T243;
  wire[4:0] T244;
  wire[4:0] T245;
  wire[4:0] T246;
  wire[4:0] T247;
  wire[4:0] T248;
  wire[4:0] T249;
  wire[4:0] T250;
  wire[4:0] T251;
  wire[4:0] T252;
  wire[4:0] T253;
  wire[4:0] T254;
  wire[3:0] T255;
  wire[3:0] T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[3:0] T262;
  wire[2:0] T263;
  wire[2:0] T264;
  wire[2:0] T265;
  wire[2:0] T266;
  wire[1:0] T267;
  wire[1:0] T268;
  wire T269;
  wire[63:0] T16;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[63:0] T17;
  wire[63:0] T332;
  wire[31:0] T18;
  wire[63:0] T19;
  wire[63:0] T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire[63:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  reg [1:0] R29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  reg  R38;
  wire T39;
  wire T40;
  wire[4:0] T41;
  reg [4:0] R42;
  wire[4:0] T43;
  wire[4:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire[2:0] T48;
  wire T49;
  wire[9:0] T50;
  wire[126:0] T51;
  wire[5:0] T52;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[5:0] T343;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[5:0] T349;
  wire[5:0] T350;
  wire[5:0] T351;
  wire[5:0] T352;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[5:0] T357;
  wire[5:0] T358;
  wire[5:0] T359;
  wire[5:0] T360;
  wire[5:0] T361;
  wire[5:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[4:0] T365;
  wire[4:0] T366;
  wire[4:0] T367;
  wire[4:0] T368;
  wire[4:0] T369;
  wire[4:0] T370;
  wire[4:0] T371;
  wire[4:0] T372;
  wire[4:0] T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire[4:0] T377;
  wire[4:0] T378;
  wire[4:0] T379;
  wire[4:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] T383;
  wire[3:0] T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[2:0] T389;
  wire[2:0] T390;
  wire[2:0] T391;
  wire[2:0] T392;
  wire[1:0] T393;
  wire[1:0] T394;
  wire T395;
  wire[63:0] T54;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire[63:0] T55;
  wire[63:0] T458;
  wire[31:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[1:0] T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T459;
  reg  R74;
  wire T460;
  reg [64:0] R75;
  wire[64:0] T76;
  reg [64:0] R77;
  wire[64:0] T78;
  wire[64:0] mux_data;
  wire[64:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[64:0] T82;
  wire[63:0] T83;
  wire[51:0] T84;
  wire[51:0] T85;
  wire[51:0] T86;
  wire[126:0] T87;
  wire[5:0] T88;
  wire[5:0] T461;
  wire[5:0] T462;
  wire[5:0] T463;
  wire[5:0] T464;
  wire[5:0] T465;
  wire[5:0] T466;
  wire[5:0] T467;
  wire[5:0] T468;
  wire[5:0] T469;
  wire[5:0] T470;
  wire[5:0] T471;
  wire[5:0] T472;
  wire[5:0] T473;
  wire[5:0] T474;
  wire[5:0] T475;
  wire[5:0] T476;
  wire[5:0] T477;
  wire[5:0] T478;
  wire[5:0] T479;
  wire[5:0] T480;
  wire[5:0] T481;
  wire[5:0] T482;
  wire[5:0] T483;
  wire[5:0] T484;
  wire[5:0] T485;
  wire[5:0] T486;
  wire[5:0] T487;
  wire[5:0] T488;
  wire[5:0] T489;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[5:0] T492;
  wire[4:0] T493;
  wire[4:0] T494;
  wire[4:0] T495;
  wire[4:0] T496;
  wire[4:0] T497;
  wire[4:0] T498;
  wire[4:0] T499;
  wire[4:0] T500;
  wire[4:0] T501;
  wire[4:0] T502;
  wire[4:0] T503;
  wire[4:0] T504;
  wire[4:0] T505;
  wire[4:0] T506;
  wire[4:0] T507;
  wire[4:0] T508;
  wire[3:0] T509;
  wire[3:0] T510;
  wire[3:0] T511;
  wire[3:0] T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[3:0] T516;
  wire[2:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire[2:0] T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire T523;
  wire[63:0] T90;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[63:0] T91;
  wire T92;
  wire[10:0] T93;
  wire[11:0] T94;
  wire[11:0] T586;
  wire[9:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[11:0] T101;
  wire[11:0] T587;
  wire[10:0] T102;
  wire[10:0] T103;
  wire[10:0] T588;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[11:0] T108;
  wire[11:0] T589;
  wire[11:0] T109;
  wire[11:0] T110;
  wire[5:0] T111;
  wire T112;
  wire[64:0] T113;
  wire[32:0] T114;
  wire[31:0] T115;
  wire[22:0] T116;
  wire[22:0] T117;
  wire[22:0] T118;
  wire[62:0] T119;
  wire[4:0] T120;
  wire[4:0] T590;
  wire[4:0] T591;
  wire[4:0] T592;
  wire[4:0] T593;
  wire[4:0] T594;
  wire[4:0] T595;
  wire[4:0] T596;
  wire[4:0] T597;
  wire[4:0] T598;
  wire[4:0] T599;
  wire[4:0] T600;
  wire[4:0] T601;
  wire[4:0] T602;
  wire[4:0] T603;
  wire[4:0] T604;
  wire[4:0] T605;
  wire[3:0] T606;
  wire[3:0] T607;
  wire[3:0] T608;
  wire[3:0] T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[3:0] T612;
  wire[3:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire[2:0] T616;
  wire[2:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire T620;
  wire[31:0] T122;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire[31:0] T123;
  wire T124;
  wire[7:0] T125;
  wire[8:0] T126;
  wire[8:0] T651;
  wire[6:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  wire[8:0] T133;
  wire[8:0] T652;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T653;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire[8:0] T140;
  wire[8:0] T654;
  wire[8:0] T141;
  wire[8:0] T142;
  wire[4:0] T143;
  wire T144;
  wire[64:0] T145;
  wire[32:0] T146;
  wire[31:0] T147;
  wire[22:0] T148;
  wire[24:0] T149;
  wire[24:0] T150;
  wire[23:0] T151;
  wire[24:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  reg [2:0] R159;
  wire[2:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire[1:0] T167;
  wire T168;
  wire[8:0] T169;
  wire[7:0] T170;
  wire[7:0] T171;
  wire[7:0] T655;
  wire T172;
  wire[7:0] T173;
  wire[6:0] T174;
  wire[5:0] T175;
  wire T176;
  wire[64:0] T177;
  wire[63:0] T178;
  wire[51:0] T179;
  wire[53:0] T180;
  wire[53:0] T181;
  wire[52:0] T182;
  wire[53:0] T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[1:0] T194;
  wire T195;
  wire[1:0] T196;
  wire T197;
  wire[11:0] T198;
  wire[10:0] T199;
  wire[10:0] T200;
  wire[10:0] T656;
  wire T201;
  wire[10:0] T202;
  wire[9:0] T203;
  wire[5:0] T204;
  wire T205;
  reg  R206;
  wire T657;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R2 = {1{$random}};
    R21 = {3{$random}};
    R29 = {1{$random}};
    R38 = {1{$random}};
    R42 = {1{$random}};
    R73 = {1{$random}};
    R74 = {1{$random}};
    R75 = {3{$random}};
    R77 = {3{$random}};
    R159 = {1{$random}};
    R206 = {1{$random}};
  end
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R74 ? R2 : R0;
  assign T3 = R73 ? mux_exc : R2;
  assign mux_exc = T4;
  assign T4 = T71 ? T44 : T5;
  assign T5 = T37 ? T6 : 5'h0;
  assign T6 = {3'h0, T7};
  assign T7 = {1'h0, T8};
  assign T8 = T9 != 2'h0;
  assign T9 = T10[1'h1:1'h0];
  assign T10 = {T36, T11};
  assign T11 = T12 != 39'h0;
  assign T12 = T13[6'h26:1'h0];
  assign T13 = T17 << T14;
  assign T14 = ~ T207;
  assign T207 = T331 ? 6'h3f : T208;
  assign T208 = T330 ? 6'h3e : T209;
  assign T209 = T329 ? 6'h3d : T210;
  assign T210 = T328 ? 6'h3c : T211;
  assign T211 = T327 ? 6'h3b : T212;
  assign T212 = T326 ? 6'h3a : T213;
  assign T213 = T325 ? 6'h39 : T214;
  assign T214 = T324 ? 6'h38 : T215;
  assign T215 = T323 ? 6'h37 : T216;
  assign T216 = T322 ? 6'h36 : T217;
  assign T217 = T321 ? 6'h35 : T218;
  assign T218 = T320 ? 6'h34 : T219;
  assign T219 = T319 ? 6'h33 : T220;
  assign T220 = T318 ? 6'h32 : T221;
  assign T221 = T317 ? 6'h31 : T222;
  assign T222 = T316 ? 6'h30 : T223;
  assign T223 = T315 ? 6'h2f : T224;
  assign T224 = T314 ? 6'h2e : T225;
  assign T225 = T313 ? 6'h2d : T226;
  assign T226 = T312 ? 6'h2c : T227;
  assign T227 = T311 ? 6'h2b : T228;
  assign T228 = T310 ? 6'h2a : T229;
  assign T229 = T309 ? 6'h29 : T230;
  assign T230 = T308 ? 6'h28 : T231;
  assign T231 = T307 ? 6'h27 : T232;
  assign T232 = T306 ? 6'h26 : T233;
  assign T233 = T305 ? 6'h25 : T234;
  assign T234 = T304 ? 6'h24 : T235;
  assign T235 = T303 ? 6'h23 : T236;
  assign T236 = T302 ? 6'h22 : T237;
  assign T237 = T301 ? 6'h21 : T238;
  assign T238 = T300 ? 6'h20 : T239;
  assign T239 = T299 ? 5'h1f : T240;
  assign T240 = T298 ? 5'h1e : T241;
  assign T241 = T297 ? 5'h1d : T242;
  assign T242 = T296 ? 5'h1c : T243;
  assign T243 = T295 ? 5'h1b : T244;
  assign T244 = T294 ? 5'h1a : T245;
  assign T245 = T293 ? 5'h19 : T246;
  assign T246 = T292 ? 5'h18 : T247;
  assign T247 = T291 ? 5'h17 : T248;
  assign T248 = T290 ? 5'h16 : T249;
  assign T249 = T289 ? 5'h15 : T250;
  assign T250 = T288 ? 5'h14 : T251;
  assign T251 = T287 ? 5'h13 : T252;
  assign T252 = T286 ? 5'h12 : T253;
  assign T253 = T285 ? 5'h11 : T254;
  assign T254 = T284 ? 5'h10 : T255;
  assign T255 = T283 ? 4'hf : T256;
  assign T256 = T282 ? 4'he : T257;
  assign T257 = T281 ? 4'hd : T258;
  assign T258 = T280 ? 4'hc : T259;
  assign T259 = T279 ? 4'hb : T260;
  assign T260 = T278 ? 4'ha : T261;
  assign T261 = T277 ? 4'h9 : T262;
  assign T262 = T276 ? 4'h8 : T263;
  assign T263 = T275 ? 3'h7 : T264;
  assign T264 = T274 ? 3'h6 : T265;
  assign T265 = T273 ? 3'h5 : T266;
  assign T266 = T272 ? 3'h4 : T267;
  assign T267 = T271 ? 2'h3 : T268;
  assign T268 = T270 ? 2'h2 : T269;
  assign T269 = T16[1'h1:1'h1];
  assign T16 = T17[6'h3f:1'h0];
  assign T270 = T16[2'h2:2'h2];
  assign T271 = T16[2'h3:2'h3];
  assign T272 = T16[3'h4:3'h4];
  assign T273 = T16[3'h5:3'h5];
  assign T274 = T16[3'h6:3'h6];
  assign T275 = T16[3'h7:3'h7];
  assign T276 = T16[4'h8:4'h8];
  assign T277 = T16[4'h9:4'h9];
  assign T278 = T16[4'ha:4'ha];
  assign T279 = T16[4'hb:4'hb];
  assign T280 = T16[4'hc:4'hc];
  assign T281 = T16[4'hd:4'hd];
  assign T282 = T16[4'he:4'he];
  assign T283 = T16[4'hf:4'hf];
  assign T284 = T16[5'h10:5'h10];
  assign T285 = T16[5'h11:5'h11];
  assign T286 = T16[5'h12:5'h12];
  assign T287 = T16[5'h13:5'h13];
  assign T288 = T16[5'h14:5'h14];
  assign T289 = T16[5'h15:5'h15];
  assign T290 = T16[5'h16:5'h16];
  assign T291 = T16[5'h17:5'h17];
  assign T292 = T16[5'h18:5'h18];
  assign T293 = T16[5'h19:5'h19];
  assign T294 = T16[5'h1a:5'h1a];
  assign T295 = T16[5'h1b:5'h1b];
  assign T296 = T16[5'h1c:5'h1c];
  assign T297 = T16[5'h1d:5'h1d];
  assign T298 = T16[5'h1e:5'h1e];
  assign T299 = T16[5'h1f:5'h1f];
  assign T300 = T16[6'h20:6'h20];
  assign T301 = T16[6'h21:6'h21];
  assign T302 = T16[6'h22:6'h22];
  assign T303 = T16[6'h23:6'h23];
  assign T304 = T16[6'h24:6'h24];
  assign T305 = T16[6'h25:6'h25];
  assign T306 = T16[6'h26:6'h26];
  assign T307 = T16[6'h27:6'h27];
  assign T308 = T16[6'h28:6'h28];
  assign T309 = T16[6'h29:6'h29];
  assign T310 = T16[6'h2a:6'h2a];
  assign T311 = T16[6'h2b:6'h2b];
  assign T312 = T16[6'h2c:6'h2c];
  assign T313 = T16[6'h2d:6'h2d];
  assign T314 = T16[6'h2e:6'h2e];
  assign T315 = T16[6'h2f:6'h2f];
  assign T316 = T16[6'h30:6'h30];
  assign T317 = T16[6'h31:6'h31];
  assign T318 = T16[6'h32:6'h32];
  assign T319 = T16[6'h33:6'h33];
  assign T320 = T16[6'h34:6'h34];
  assign T321 = T16[6'h35:6'h35];
  assign T322 = T16[6'h36:6'h36];
  assign T323 = T16[6'h37:6'h37];
  assign T324 = T16[6'h38:6'h38];
  assign T325 = T16[6'h39:6'h39];
  assign T326 = T16[6'h3a:6'h3a];
  assign T327 = T16[6'h3b:6'h3b];
  assign T328 = T16[6'h3c:6'h3c];
  assign T329 = T16[6'h3d:6'h3d];
  assign T330 = T16[6'h3e:6'h3e];
  assign T331 = T16[6'h3f:6'h3f];
  assign T17 = T33 ? T19 : T332;
  assign T332 = {32'h0, T18};
  assign T18 = T19[5'h1f:1'h0];
  assign T19 = T24 ? T23 : T20;
  assign T20 = R21[6'h3f:1'h0];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = 64'h0 - T20;
  assign T24 = T32 ? T31 : T25;
  assign T25 = T27 ? T26 : 1'h0;
  assign T26 = T20[6'h3f:6'h3f];
  assign T27 = T28 == 2'h3;
  assign T28 = R29 ^ 2'h1;
  assign T30 = io_in_valid ? io_in_bits_typ : R29;
  assign T31 = T20[5'h1f:5'h1f];
  assign T32 = T28 == 2'h1;
  assign T33 = T35 | T34;
  assign T34 = T28 == 2'h2;
  assign T35 = T28 == 2'h3;
  assign T36 = T13[6'h28:6'h27];
  assign T37 = T40 & R38;
  assign T39 = io_in_valid ? io_in_bits_single : R38;
  assign T40 = T41 == 5'h0;
  assign T41 = R42 & 5'h4;
  assign T43 = io_in_valid ? io_in_bits_cmd : R42;
  assign T44 = {3'h0, T45};
  assign T45 = {1'h0, T46};
  assign T46 = T47 != 2'h0;
  assign T47 = T48[1'h1:1'h0];
  assign T48 = {T70, T49};
  assign T49 = T50 != 10'h0;
  assign T50 = T51[4'h9:1'h0];
  assign T51 = T55 << T52;
  assign T52 = ~ T333;
  assign T333 = T457 ? 6'h3f : T334;
  assign T334 = T456 ? 6'h3e : T335;
  assign T335 = T455 ? 6'h3d : T336;
  assign T336 = T454 ? 6'h3c : T337;
  assign T337 = T453 ? 6'h3b : T338;
  assign T338 = T452 ? 6'h3a : T339;
  assign T339 = T451 ? 6'h39 : T340;
  assign T340 = T450 ? 6'h38 : T341;
  assign T341 = T449 ? 6'h37 : T342;
  assign T342 = T448 ? 6'h36 : T343;
  assign T343 = T447 ? 6'h35 : T344;
  assign T344 = T446 ? 6'h34 : T345;
  assign T345 = T445 ? 6'h33 : T346;
  assign T346 = T444 ? 6'h32 : T347;
  assign T347 = T443 ? 6'h31 : T348;
  assign T348 = T442 ? 6'h30 : T349;
  assign T349 = T441 ? 6'h2f : T350;
  assign T350 = T440 ? 6'h2e : T351;
  assign T351 = T439 ? 6'h2d : T352;
  assign T352 = T438 ? 6'h2c : T353;
  assign T353 = T437 ? 6'h2b : T354;
  assign T354 = T436 ? 6'h2a : T355;
  assign T355 = T435 ? 6'h29 : T356;
  assign T356 = T434 ? 6'h28 : T357;
  assign T357 = T433 ? 6'h27 : T358;
  assign T358 = T432 ? 6'h26 : T359;
  assign T359 = T431 ? 6'h25 : T360;
  assign T360 = T430 ? 6'h24 : T361;
  assign T361 = T429 ? 6'h23 : T362;
  assign T362 = T428 ? 6'h22 : T363;
  assign T363 = T427 ? 6'h21 : T364;
  assign T364 = T426 ? 6'h20 : T365;
  assign T365 = T425 ? 5'h1f : T366;
  assign T366 = T424 ? 5'h1e : T367;
  assign T367 = T423 ? 5'h1d : T368;
  assign T368 = T422 ? 5'h1c : T369;
  assign T369 = T421 ? 5'h1b : T370;
  assign T370 = T420 ? 5'h1a : T371;
  assign T371 = T419 ? 5'h19 : T372;
  assign T372 = T418 ? 5'h18 : T373;
  assign T373 = T417 ? 5'h17 : T374;
  assign T374 = T416 ? 5'h16 : T375;
  assign T375 = T415 ? 5'h15 : T376;
  assign T376 = T414 ? 5'h14 : T377;
  assign T377 = T413 ? 5'h13 : T378;
  assign T378 = T412 ? 5'h12 : T379;
  assign T379 = T411 ? 5'h11 : T380;
  assign T380 = T410 ? 5'h10 : T381;
  assign T381 = T409 ? 4'hf : T382;
  assign T382 = T408 ? 4'he : T383;
  assign T383 = T407 ? 4'hd : T384;
  assign T384 = T406 ? 4'hc : T385;
  assign T385 = T405 ? 4'hb : T386;
  assign T386 = T404 ? 4'ha : T387;
  assign T387 = T403 ? 4'h9 : T388;
  assign T388 = T402 ? 4'h8 : T389;
  assign T389 = T401 ? 3'h7 : T390;
  assign T390 = T400 ? 3'h6 : T391;
  assign T391 = T399 ? 3'h5 : T392;
  assign T392 = T398 ? 3'h4 : T393;
  assign T393 = T397 ? 2'h3 : T394;
  assign T394 = T396 ? 2'h2 : T395;
  assign T395 = T54[1'h1:1'h1];
  assign T54 = T55[6'h3f:1'h0];
  assign T396 = T54[2'h2:2'h2];
  assign T397 = T54[2'h3:2'h3];
  assign T398 = T54[3'h4:3'h4];
  assign T399 = T54[3'h5:3'h5];
  assign T400 = T54[3'h6:3'h6];
  assign T401 = T54[3'h7:3'h7];
  assign T402 = T54[4'h8:4'h8];
  assign T403 = T54[4'h9:4'h9];
  assign T404 = T54[4'ha:4'ha];
  assign T405 = T54[4'hb:4'hb];
  assign T406 = T54[4'hc:4'hc];
  assign T407 = T54[4'hd:4'hd];
  assign T408 = T54[4'he:4'he];
  assign T409 = T54[4'hf:4'hf];
  assign T410 = T54[5'h10:5'h10];
  assign T411 = T54[5'h11:5'h11];
  assign T412 = T54[5'h12:5'h12];
  assign T413 = T54[5'h13:5'h13];
  assign T414 = T54[5'h14:5'h14];
  assign T415 = T54[5'h15:5'h15];
  assign T416 = T54[5'h16:5'h16];
  assign T417 = T54[5'h17:5'h17];
  assign T418 = T54[5'h18:5'h18];
  assign T419 = T54[5'h19:5'h19];
  assign T420 = T54[5'h1a:5'h1a];
  assign T421 = T54[5'h1b:5'h1b];
  assign T422 = T54[5'h1c:5'h1c];
  assign T423 = T54[5'h1d:5'h1d];
  assign T424 = T54[5'h1e:5'h1e];
  assign T425 = T54[5'h1f:5'h1f];
  assign T426 = T54[6'h20:6'h20];
  assign T427 = T54[6'h21:6'h21];
  assign T428 = T54[6'h22:6'h22];
  assign T429 = T54[6'h23:6'h23];
  assign T430 = T54[6'h24:6'h24];
  assign T431 = T54[6'h25:6'h25];
  assign T432 = T54[6'h26:6'h26];
  assign T433 = T54[6'h27:6'h27];
  assign T434 = T54[6'h28:6'h28];
  assign T435 = T54[6'h29:6'h29];
  assign T436 = T54[6'h2a:6'h2a];
  assign T437 = T54[6'h2b:6'h2b];
  assign T438 = T54[6'h2c:6'h2c];
  assign T439 = T54[6'h2d:6'h2d];
  assign T440 = T54[6'h2e:6'h2e];
  assign T441 = T54[6'h2f:6'h2f];
  assign T442 = T54[6'h30:6'h30];
  assign T443 = T54[6'h31:6'h31];
  assign T444 = T54[6'h32:6'h32];
  assign T445 = T54[6'h33:6'h33];
  assign T446 = T54[6'h34:6'h34];
  assign T447 = T54[6'h35:6'h35];
  assign T448 = T54[6'h36:6'h36];
  assign T449 = T54[6'h37:6'h37];
  assign T450 = T54[6'h38:6'h38];
  assign T451 = T54[6'h39:6'h39];
  assign T452 = T54[6'h3a:6'h3a];
  assign T453 = T54[6'h3b:6'h3b];
  assign T454 = T54[6'h3c:6'h3c];
  assign T455 = T54[6'h3d:6'h3d];
  assign T456 = T54[6'h3e:6'h3e];
  assign T457 = T54[6'h3f:6'h3f];
  assign T55 = T67 ? T57 : T458;
  assign T458 = {32'h0, T56};
  assign T56 = T57[5'h1f:1'h0];
  assign T57 = T60 ? T59 : T58;
  assign T58 = R21[6'h3f:1'h0];
  assign T59 = 64'h0 - T58;
  assign T60 = T66 ? T65 : T61;
  assign T61 = T63 ? T62 : 1'h0;
  assign T62 = T58[6'h3f:6'h3f];
  assign T63 = T64 == 2'h3;
  assign T64 = R29 ^ 2'h1;
  assign T65 = T58[5'h1f:5'h1f];
  assign T66 = T64 == 2'h1;
  assign T67 = T69 | T68;
  assign T68 = T64 == 2'h2;
  assign T69 = T64 == 2'h3;
  assign T70 = T51[4'hb:4'ha];
  assign T71 = T40 & T72;
  assign T72 = R38 ^ 1'h1;
  assign T459 = reset ? 1'h0 : io_in_valid;
  assign T460 = reset ? 1'h0 : R73;
  assign io_out_bits_data = R75;
  assign T76 = R74 ? R77 : R75;
  assign T78 = R73 ? mux_data : R77;
  assign mux_data = T79;
  assign T79 = T71 ? T177 : T80;
  assign T80 = T37 ? T145 : T81;
  assign T81 = R38 ? T113 : T82;
  assign T82 = {T112, T83};
  assign T83 = {T94, T84};
  assign T84 = T92 ? T86 : T85;
  assign T85 = R21[6'h33:1'h0];
  assign T86 = T87[6'h3e:4'hb];
  assign T87 = T91 << T88;
  assign T88 = ~ T461;
  assign T461 = T585 ? 6'h3f : T462;
  assign T462 = T584 ? 6'h3e : T463;
  assign T463 = T583 ? 6'h3d : T464;
  assign T464 = T582 ? 6'h3c : T465;
  assign T465 = T581 ? 6'h3b : T466;
  assign T466 = T580 ? 6'h3a : T467;
  assign T467 = T579 ? 6'h39 : T468;
  assign T468 = T578 ? 6'h38 : T469;
  assign T469 = T577 ? 6'h37 : T470;
  assign T470 = T576 ? 6'h36 : T471;
  assign T471 = T575 ? 6'h35 : T472;
  assign T472 = T574 ? 6'h34 : T473;
  assign T473 = T573 ? 6'h33 : T474;
  assign T474 = T572 ? 6'h32 : T475;
  assign T475 = T571 ? 6'h31 : T476;
  assign T476 = T570 ? 6'h30 : T477;
  assign T477 = T569 ? 6'h2f : T478;
  assign T478 = T568 ? 6'h2e : T479;
  assign T479 = T567 ? 6'h2d : T480;
  assign T480 = T566 ? 6'h2c : T481;
  assign T481 = T565 ? 6'h2b : T482;
  assign T482 = T564 ? 6'h2a : T483;
  assign T483 = T563 ? 6'h29 : T484;
  assign T484 = T562 ? 6'h28 : T485;
  assign T485 = T561 ? 6'h27 : T486;
  assign T486 = T560 ? 6'h26 : T487;
  assign T487 = T559 ? 6'h25 : T488;
  assign T488 = T558 ? 6'h24 : T489;
  assign T489 = T557 ? 6'h23 : T490;
  assign T490 = T556 ? 6'h22 : T491;
  assign T491 = T555 ? 6'h21 : T492;
  assign T492 = T554 ? 6'h20 : T493;
  assign T493 = T553 ? 5'h1f : T494;
  assign T494 = T552 ? 5'h1e : T495;
  assign T495 = T551 ? 5'h1d : T496;
  assign T496 = T550 ? 5'h1c : T497;
  assign T497 = T549 ? 5'h1b : T498;
  assign T498 = T548 ? 5'h1a : T499;
  assign T499 = T547 ? 5'h19 : T500;
  assign T500 = T546 ? 5'h18 : T501;
  assign T501 = T545 ? 5'h17 : T502;
  assign T502 = T544 ? 5'h16 : T503;
  assign T503 = T543 ? 5'h15 : T504;
  assign T504 = T542 ? 5'h14 : T505;
  assign T505 = T541 ? 5'h13 : T506;
  assign T506 = T540 ? 5'h12 : T507;
  assign T507 = T539 ? 5'h11 : T508;
  assign T508 = T538 ? 5'h10 : T509;
  assign T509 = T537 ? 4'hf : T510;
  assign T510 = T536 ? 4'he : T511;
  assign T511 = T535 ? 4'hd : T512;
  assign T512 = T534 ? 4'hc : T513;
  assign T513 = T533 ? 4'hb : T514;
  assign T514 = T532 ? 4'ha : T515;
  assign T515 = T531 ? 4'h9 : T516;
  assign T516 = T530 ? 4'h8 : T517;
  assign T517 = T529 ? 3'h7 : T518;
  assign T518 = T528 ? 3'h6 : T519;
  assign T519 = T527 ? 3'h5 : T520;
  assign T520 = T526 ? 3'h4 : T521;
  assign T521 = T525 ? 2'h3 : T522;
  assign T522 = T524 ? 2'h2 : T523;
  assign T523 = T90[1'h1:1'h1];
  assign T90 = T91[6'h3f:1'h0];
  assign T524 = T90[2'h2:2'h2];
  assign T525 = T90[2'h3:2'h3];
  assign T526 = T90[3'h4:3'h4];
  assign T527 = T90[3'h5:3'h5];
  assign T528 = T90[3'h6:3'h6];
  assign T529 = T90[3'h7:3'h7];
  assign T530 = T90[4'h8:4'h8];
  assign T531 = T90[4'h9:4'h9];
  assign T532 = T90[4'ha:4'ha];
  assign T533 = T90[4'hb:4'hb];
  assign T534 = T90[4'hc:4'hc];
  assign T535 = T90[4'hd:4'hd];
  assign T536 = T90[4'he:4'he];
  assign T537 = T90[4'hf:4'hf];
  assign T538 = T90[5'h10:5'h10];
  assign T539 = T90[5'h11:5'h11];
  assign T540 = T90[5'h12:5'h12];
  assign T541 = T90[5'h13:5'h13];
  assign T542 = T90[5'h14:5'h14];
  assign T543 = T90[5'h15:5'h15];
  assign T544 = T90[5'h16:5'h16];
  assign T545 = T90[5'h17:5'h17];
  assign T546 = T90[5'h18:5'h18];
  assign T547 = T90[5'h19:5'h19];
  assign T548 = T90[5'h1a:5'h1a];
  assign T549 = T90[5'h1b:5'h1b];
  assign T550 = T90[5'h1c:5'h1c];
  assign T551 = T90[5'h1d:5'h1d];
  assign T552 = T90[5'h1e:5'h1e];
  assign T553 = T90[5'h1f:5'h1f];
  assign T554 = T90[6'h20:6'h20];
  assign T555 = T90[6'h21:6'h21];
  assign T556 = T90[6'h22:6'h22];
  assign T557 = T90[6'h23:6'h23];
  assign T558 = T90[6'h24:6'h24];
  assign T559 = T90[6'h25:6'h25];
  assign T560 = T90[6'h26:6'h26];
  assign T561 = T90[6'h27:6'h27];
  assign T562 = T90[6'h28:6'h28];
  assign T563 = T90[6'h29:6'h29];
  assign T564 = T90[6'h2a:6'h2a];
  assign T565 = T90[6'h2b:6'h2b];
  assign T566 = T90[6'h2c:6'h2c];
  assign T567 = T90[6'h2d:6'h2d];
  assign T568 = T90[6'h2e:6'h2e];
  assign T569 = T90[6'h2f:6'h2f];
  assign T570 = T90[6'h30:6'h30];
  assign T571 = T90[6'h31:6'h31];
  assign T572 = T90[6'h32:6'h32];
  assign T573 = T90[6'h33:6'h33];
  assign T574 = T90[6'h34:6'h34];
  assign T575 = T90[6'h35:6'h35];
  assign T576 = T90[6'h36:6'h36];
  assign T577 = T90[6'h37:6'h37];
  assign T578 = T90[6'h38:6'h38];
  assign T579 = T90[6'h39:6'h39];
  assign T580 = T90[6'h3a:6'h3a];
  assign T581 = T90[6'h3b:6'h3b];
  assign T582 = T90[6'h3c:6'h3c];
  assign T583 = T90[6'h3d:6'h3d];
  assign T584 = T90[6'h3e:6'h3e];
  assign T585 = T90[6'h3f:6'h3f];
  assign T91 = T85 << 4'hc;
  assign T92 = T93 == 11'h0;
  assign T93 = R21[6'h3e:6'h34];
  assign T94 = T101 | T586;
  assign T586 = {2'h0, T95};
  assign T95 = T96 << 4'h9;
  assign T96 = T99 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T85 == 52'h0;
  assign T99 = T100 == 2'h3;
  assign T100 = T101[4'hb:4'ha];
  assign T101 = T108 + T587;
  assign T587 = {1'h0, T102};
  assign T102 = T107 ? 11'h0 : T103;
  assign T103 = 11'h400 | T588;
  assign T588 = {9'h0, T104};
  assign T104 = T105 ? 2'h2 : 2'h1;
  assign T105 = T92 & T106;
  assign T106 = T98 ^ 1'h1;
  assign T107 = T92 & T98;
  assign T108 = T92 ? T109 : T589;
  assign T589 = {1'h0, T93};
  assign T109 = T98 ? 12'h0 : T110;
  assign T110 = {6'h3f, T111};
  assign T111 = ~ T88;
  assign T112 = R21[6'h3f:6'h3f];
  assign T113 = {32'hffffffff, T114};
  assign T114 = {T144, T115};
  assign T115 = {T126, T116};
  assign T116 = T124 ? T118 : T117;
  assign T117 = R21[5'h16:1'h0];
  assign T118 = T119[5'h1e:4'h8];
  assign T119 = T123 << T120;
  assign T120 = ~ T590;
  assign T590 = T650 ? 5'h1f : T591;
  assign T591 = T649 ? 5'h1e : T592;
  assign T592 = T648 ? 5'h1d : T593;
  assign T593 = T647 ? 5'h1c : T594;
  assign T594 = T646 ? 5'h1b : T595;
  assign T595 = T645 ? 5'h1a : T596;
  assign T596 = T644 ? 5'h19 : T597;
  assign T597 = T643 ? 5'h18 : T598;
  assign T598 = T642 ? 5'h17 : T599;
  assign T599 = T641 ? 5'h16 : T600;
  assign T600 = T640 ? 5'h15 : T601;
  assign T601 = T639 ? 5'h14 : T602;
  assign T602 = T638 ? 5'h13 : T603;
  assign T603 = T637 ? 5'h12 : T604;
  assign T604 = T636 ? 5'h11 : T605;
  assign T605 = T635 ? 5'h10 : T606;
  assign T606 = T634 ? 4'hf : T607;
  assign T607 = T633 ? 4'he : T608;
  assign T608 = T632 ? 4'hd : T609;
  assign T609 = T631 ? 4'hc : T610;
  assign T610 = T630 ? 4'hb : T611;
  assign T611 = T629 ? 4'ha : T612;
  assign T612 = T628 ? 4'h9 : T613;
  assign T613 = T627 ? 4'h8 : T614;
  assign T614 = T626 ? 3'h7 : T615;
  assign T615 = T625 ? 3'h6 : T616;
  assign T616 = T624 ? 3'h5 : T617;
  assign T617 = T623 ? 3'h4 : T618;
  assign T618 = T622 ? 2'h3 : T619;
  assign T619 = T621 ? 2'h2 : T620;
  assign T620 = T122[1'h1:1'h1];
  assign T122 = T123[5'h1f:1'h0];
  assign T621 = T122[2'h2:2'h2];
  assign T622 = T122[2'h3:2'h3];
  assign T623 = T122[3'h4:3'h4];
  assign T624 = T122[3'h5:3'h5];
  assign T625 = T122[3'h6:3'h6];
  assign T626 = T122[3'h7:3'h7];
  assign T627 = T122[4'h8:4'h8];
  assign T628 = T122[4'h9:4'h9];
  assign T629 = T122[4'ha:4'ha];
  assign T630 = T122[4'hb:4'hb];
  assign T631 = T122[4'hc:4'hc];
  assign T632 = T122[4'hd:4'hd];
  assign T633 = T122[4'he:4'he];
  assign T634 = T122[4'hf:4'hf];
  assign T635 = T122[5'h10:5'h10];
  assign T636 = T122[5'h11:5'h11];
  assign T637 = T122[5'h12:5'h12];
  assign T638 = T122[5'h13:5'h13];
  assign T639 = T122[5'h14:5'h14];
  assign T640 = T122[5'h15:5'h15];
  assign T641 = T122[5'h16:5'h16];
  assign T642 = T122[5'h17:5'h17];
  assign T643 = T122[5'h18:5'h18];
  assign T644 = T122[5'h19:5'h19];
  assign T645 = T122[5'h1a:5'h1a];
  assign T646 = T122[5'h1b:5'h1b];
  assign T647 = T122[5'h1c:5'h1c];
  assign T648 = T122[5'h1d:5'h1d];
  assign T649 = T122[5'h1e:5'h1e];
  assign T650 = T122[5'h1f:5'h1f];
  assign T123 = T117 << 4'h9;
  assign T124 = T125 == 8'h0;
  assign T125 = R21[5'h1e:5'h17];
  assign T126 = T133 | T651;
  assign T651 = {2'h0, T127};
  assign T127 = T128 << 3'h6;
  assign T128 = T131 & T129;
  assign T129 = T130 ^ 1'h1;
  assign T130 = T117 == 23'h0;
  assign T131 = T132 == 2'h3;
  assign T132 = T133[4'h8:3'h7];
  assign T133 = T140 + T652;
  assign T652 = {1'h0, T134};
  assign T134 = T139 ? 8'h0 : T135;
  assign T135 = 8'h80 | T653;
  assign T653 = {6'h0, T136};
  assign T136 = T137 ? 2'h2 : 2'h1;
  assign T137 = T124 & T138;
  assign T138 = T130 ^ 1'h1;
  assign T139 = T124 & T130;
  assign T140 = T124 ? T141 : T654;
  assign T654 = {1'h0, T125};
  assign T141 = T130 ? 9'h0 : T142;
  assign T142 = {4'hf, T143};
  assign T143 = ~ T120;
  assign T144 = R21[5'h1f:5'h1f];
  assign T145 = {32'hffffffff, T146};
  assign T146 = {T24, T147};
  assign T147 = {T169, T148};
  assign T148 = T149[5'h16:1'h0];
  assign T149 = T153 ? T152 : T150;
  assign T150 = {1'h0, T151};
  assign T151 = T13[6'h3f:6'h28];
  assign T152 = T150 + 25'h1;
  assign T153 = T168 ? T163 : T154;
  assign T154 = T162 ? T161 : T155;
  assign T155 = T158 ? T156 : 1'h0;
  assign T156 = T157 & T8;
  assign T157 = T24 ^ 1'h1;
  assign T158 = R159 == 3'h3;
  assign T160 = io_in_valid ? io_in_bits_rm : R159;
  assign T161 = T24 & T8;
  assign T162 = R159 == 3'h2;
  assign T163 = T166 | T164;
  assign T164 = T165 == 2'h3;
  assign T165 = T10[1'h1:1'h0];
  assign T166 = T167 == 2'h3;
  assign T167 = T10[2'h2:1'h1];
  assign T168 = R159 == 3'h0;
  assign T169 = {T176, T170};
  assign T170 = T171[3'h7:1'h0];
  assign T171 = T173 + T655;
  assign T655 = {7'h0, T172};
  assign T172 = T149[5'h18:5'h18];
  assign T173 = {1'h0, T174};
  assign T174 = {1'h0, T175};
  assign T175 = ~ T14;
  assign T176 = T13[6'h3f:6'h3f];
  assign T177 = {T60, T178};
  assign T178 = {T198, T179};
  assign T179 = T180[6'h33:1'h0];
  assign T180 = T184 ? T183 : T181;
  assign T181 = {1'h0, T182};
  assign T182 = T51[6'h3f:4'hb];
  assign T183 = T181 + 54'h1;
  assign T184 = T197 ? T192 : T185;
  assign T185 = T191 ? T190 : T186;
  assign T186 = T189 ? T187 : 1'h0;
  assign T187 = T188 & T46;
  assign T188 = T60 ^ 1'h1;
  assign T189 = R159 == 3'h3;
  assign T190 = T60 & T46;
  assign T191 = R159 == 3'h2;
  assign T192 = T195 | T193;
  assign T193 = T194 == 2'h3;
  assign T194 = T48[1'h1:1'h0];
  assign T195 = T196 == 2'h3;
  assign T196 = T48[2'h2:1'h1];
  assign T197 = R159 == 3'h0;
  assign T198 = {T205, T199};
  assign T199 = T200[4'ha:1'h0];
  assign T200 = T202 + T656;
  assign T656 = {10'h0, T201};
  assign T201 = T180[6'h35:6'h35];
  assign T202 = {1'h0, T203};
  assign T203 = {4'h0, T204};
  assign T204 = ~ T52;
  assign T205 = T51[6'h3f:6'h3f];
  assign io_out_valid = R206;
  assign T657 = reset ? 1'h0 : R74;

  always @(posedge clk) begin
    if(R74) begin
      R0 <= R2;
    end
    if(R73) begin
      R2 <= mux_exc;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R29 <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      R38 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R42 <= io_in_bits_cmd;
    end
    if(reset) begin
      R73 <= 1'h0;
    end else begin
      R73 <= io_in_valid;
    end
    if(reset) begin
      R74 <= 1'h0;
    end else begin
      R74 <= R73;
    end
    if(R74) begin
      R75 <= R77;
    end
    if(R73) begin
      R77 <= mux_data;
    end
    if(io_in_valid) begin
      R159 <= io_in_bits_rm;
    end
    if(reset) begin
      R206 <= 1'h0;
    end else begin
      R206 <= R74;
    end
  end
endmodule

module FPToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc,
    input  io_lt
);

  reg [4:0] R0;
  wire[4:0] T1;
  wire[4:0] mux_exc;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] minmax_exc;
  wire T5;
  wire issnan2;
  wire T6;
  wire T7;
  wire T8;
  reg [64:0] R9;
  wire[64:0] T10;
  wire T11;
  reg  R12;
  wire T13;
  wire isnan2;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire issnan1;
  wire T18;
  wire T19;
  wire T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire T23;
  wire isnan1;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire isSgnj;
  wire[4:0] T28;
  reg [4:0] R29;
  wire[4:0] T30;
  wire[4:0] T31;
  wire[2:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[2:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire[11:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[1:0] T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire[27:0] T56;
  wire[51:0] T57;
  wire T58;
  wire[23:0] T59;
  wire[48:0] T60;
  wire[4:0] T61;
  wire[11:0] T62;
  wire[11:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire[48:0] T67;
  wire[47:0] T68;
  wire[23:0] T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[24:0] T76;
  wire[24:0] T77;
  wire[24:0] T78;
  wire[24:0] T79;
  wire[55:0] T80;
  wire[4:0] T81;
  wire[24:0] T82;
  wire[22:0] T83;
  wire[24:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  reg [2:0] R92;
  wire[2:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[1:0] T98;
  wire T99;
  wire[1:0] T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire[4:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[22:0] T115;
  wire T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  reg  R120;
  wire T200;
  reg [64:0] R121;
  wire[64:0] T122;
  wire[64:0] mux_data;
  wire[64:0] T123;
  wire[64:0] T124;
  wire[64:0] T125;
  wire[64:0] fsgnj;
  wire[32:0] T126;
  wire[31:0] T127;
  wire sign_s;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire sign_d;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire isLHS;
  wire T150;
  wire T151;
  wire T152;
  wire isMax;
  wire[64:0] T153;
  wire[32:0] T154;
  wire[31:0] T155;
  wire[22:0] T156;
  wire[22:0] T157;
  wire[22:0] T158;
  wire[22:0] T159;
  wire[22:0] T160;
  wire[22:0] T201;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[22:0] T170;
  wire[22:0] T202;
  wire[8:0] T171;
  wire[8:0] T172;
  wire[8:0] T173;
  wire[8:0] T174;
  wire[8:0] T175;
  wire[8:0] T176;
  wire[8:0] T177;
  wire T178;
  wire[8:0] T203;
  wire[6:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire[64:0] T182;
  wire[63:0] T183;
  wire[51:0] T184;
  wire[51:0] T185;
  wire[51:0] T186;
  wire[51:0] T204;
  wire[11:0] T187;
  wire[11:0] T188;
  wire[11:0] T189;
  wire[11:0] T190;
  wire T191;
  wire[11:0] T192;
  wire[7:0] T196;
  wire T193;
  wire[11:0] T205;
  wire[10:0] T194;
  wire T195;
  wire[11:0] T206;
  wire T197;
  wire T198;
  reg  R199;
  wire T207;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R9 = {3{$random}};
    R12 = {1{$random}};
    R21 = {3{$random}};
    R29 = {1{$random}};
    R92 = {1{$random}};
    R120 = {1{$random}};
    R121 = {3{$random}};
    R199 = {1{$random}};
  end
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R120 ? mux_exc : R0;
  assign mux_exc = T2;
  assign T2 = T118 ? T111 : T3;
  assign T3 = T108 ? T31 : T4;
  assign T4 = isSgnj ? 5'h0 : minmax_exc;
  assign minmax_exc = {T5, 4'h0};
  assign T5 = issnan1 | issnan2;
  assign issnan2 = isnan2 & T6;
  assign T6 = ~ T7;
  assign T7 = R12 ? T11 : T8;
  assign T8 = R9[6'h33:6'h33];
  assign T10 = io_in_valid ? io_in_bits_in2 : R9;
  assign T11 = R9[5'h16:5'h16];
  assign T13 = io_in_valid ? io_in_bits_single : R12;
  assign isnan2 = R12 ? T16 : T14;
  assign T14 = T15 == 3'h7;
  assign T15 = R9[6'h3f:6'h3d];
  assign T16 = T17 == 3'h7;
  assign T17 = R9[5'h1f:5'h1d];
  assign issnan1 = isnan1 & T18;
  assign T18 = ~ T19;
  assign T19 = R12 ? T23 : T20;
  assign T20 = R21[6'h33:6'h33];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = R21[5'h16:5'h16];
  assign isnan1 = R12 ? T26 : T24;
  assign T24 = T25 == 3'h7;
  assign T25 = R21[6'h3f:6'h3d];
  assign T26 = T27 == 3'h7;
  assign T27 = R21[5'h1f:5'h1d];
  assign isSgnj = T28 == 5'h4;
  assign T28 = R29 & 5'h5;
  assign T30 = io_in_valid ? io_in_bits_cmd : R29;
  assign T31 = {T103, T32};
  assign T32 = {T73, T33};
  assign T33 = {T71, T34};
  assign T34 = T45 | T35;
  assign T35 = T43 & T36;
  assign T36 = T37 ^ 1'h1;
  assign T37 = T41 | T38;
  assign T38 = T39 == 2'h3;
  assign T39 = T40[2'h2:1'h1];
  assign T40 = R21[6'h3f:6'h3d];
  assign T41 = T42 ^ 1'h1;
  assign T42 = T40 != 3'h0;
  assign T43 = T44 < 12'h76a;
  assign T44 = R21[6'h3f:6'h34];
  assign T45 = T49 | T46;
  assign T46 = T48 & T47;
  assign T47 = T37 ^ 1'h1;
  assign T48 = 12'h87f < T44;
  assign T49 = T51 & T50;
  assign T50 = T37 ^ 1'h1;
  assign T51 = T52 != 2'h0;
  assign T52 = T53[1'h1:1'h0];
  assign T53 = {T70, T54};
  assign T54 = T58 | T55;
  assign T55 = T56 != 28'h0;
  assign T56 = T57[5'h1b:1'h0];
  assign T57 = R21[6'h33:1'h0];
  assign T58 = T59 != 24'h0;
  assign T59 = T60[5'h17:1'h0];
  assign T60 = T67 >> T61;
  assign T61 = T62[3'h4:1'h0];
  assign T62 = T64 ? T63 : 12'h0;
  assign T63 = 12'h782 - T44;
  assign T64 = T66 & T65;
  assign T65 = T44 <= 12'h781;
  assign T66 = 12'h76a <= T44;
  assign T67 = {1'h1, T68};
  assign T68 = {T69, 24'h0};
  assign T69 = T57[6'h33:5'h1c];
  assign T70 = T60[5'h19:5'h18];
  assign T71 = T35 | T72;
  assign T72 = T64 & T49;
  assign T73 = T46 | T74;
  assign T74 = T102 & T75;
  assign T75 = T76[5'h18:5'h18];
  assign T76 = T85 ? T84 : T77;
  assign T77 = T82 | T78;
  assign T78 = ~ T79;
  assign T79 = T80[5'h18:1'h0];
  assign T80 = 25'h1ffffff << T81;
  assign T81 = T61;
  assign T82 = {2'h1, T83};
  assign T83 = T57[6'h33:5'h1d];
  assign T84 = T77 + 25'h1;
  assign T85 = T101 ? T96 : T86;
  assign T86 = T95 ? T94 : T87;
  assign T87 = T91 ? T88 : 1'h0;
  assign T88 = T89 & T49;
  assign T89 = T90 ^ 1'h1;
  assign T90 = R21[7'h40:7'h40];
  assign T91 = R92 == 3'h3;
  assign T93 = io_in_valid ? io_in_bits_rm : R92;
  assign T94 = T90 & T49;
  assign T95 = R92 == 3'h2;
  assign T96 = T99 | T97;
  assign T97 = T98 == 2'h3;
  assign T98 = T53[2'h2:1'h1];
  assign T99 = T100 == 2'h3;
  assign T100 = T53[1'h1:1'h0];
  assign T101 = R92 == 3'h0;
  assign T102 = T44 == 12'h87f;
  assign T103 = {T104, 1'h0};
  assign T104 = T107 & T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = T57[6'h33:6'h33];
  assign T107 = T40 == 3'h7;
  assign T108 = T109 & R12;
  assign T109 = T110 == 5'h0;
  assign T110 = R29 & 5'h4;
  assign T111 = T112 << 3'h4;
  assign T112 = T116 & T113;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115[5'h16:5'h16];
  assign T115 = R21[5'h16:1'h0];
  assign T116 = T117 == 3'h7;
  assign T117 = R21[5'h1f:5'h1d];
  assign T118 = T109 & T119;
  assign T119 = R12 ^ 1'h1;
  assign T200 = reset ? 1'h0 : io_in_valid;
  assign io_out_bits_data = R121;
  assign T122 = R120 ? mux_data : R121;
  assign mux_data = T123;
  assign T123 = T118 ? T182 : T124;
  assign T124 = T108 ? T153 : T125;
  assign T125 = T149 ? fsgnj : R9;
  assign fsgnj = {T137, T126};
  assign T126 = {sign_s, T127};
  assign T127 = R21[5'h1f:1'h0];
  assign sign_s = T131 ^ T128;
  assign T128 = T130 & T129;
  assign T129 = R9[6'h20:6'h20];
  assign T130 = R12 & isSgnj;
  assign T131 = T134 ? T133 : T132;
  assign T132 = R92[1'h0:1'h0];
  assign T133 = R21[6'h20:6'h20];
  assign T134 = T136 | T135;
  assign T135 = T130 ^ 1'h1;
  assign T136 = R92[1'h1:1'h1];
  assign T137 = {sign_d, T138};
  assign T138 = R21[6'h3f:6'h21];
  assign sign_d = T143 ^ T139;
  assign T139 = T141 & T140;
  assign T140 = R9[7'h40:7'h40];
  assign T141 = T142 & isSgnj;
  assign T142 = R12 ^ 1'h1;
  assign T143 = T146 ? T145 : T144;
  assign T144 = R92[1'h0:1'h0];
  assign T145 = R21[7'h40:7'h40];
  assign T146 = T148 | T147;
  assign T147 = T141 ^ 1'h1;
  assign T148 = R92[1'h1:1'h1];
  assign T149 = isSgnj | isLHS;
  assign isLHS = isnan2 | T150;
  assign T150 = T152 & T151;
  assign T151 = isnan1 ^ 1'h1;
  assign T152 = isMax != io_lt;
  assign isMax = R92[1'h0:1'h0];
  assign T153 = {32'hffffffff, T154};
  assign T154 = {T90, T155};
  assign T155 = {T171, T156};
  assign T156 = T37 ? T170 : T157;
  assign T157 = T46 ? T160 : T158;
  assign T158 = T35 ? 23'h0 : T159;
  assign T159 = T76[5'h16:1'h0];
  assign T160 = 23'h0 - T201;
  assign T201 = {22'h0, T161};
  assign T161 = T162 ^ 1'h1;
  assign T162 = T164 | T163;
  assign T163 = R92 == 3'h0;
  assign T164 = T168 | T165;
  assign T165 = T167 & T166;
  assign T166 = T90 ^ 1'h1;
  assign T167 = R92 == 3'h3;
  assign T168 = T169 & T90;
  assign T169 = R92 == 3'h2;
  assign T170 = 23'h0 - T202;
  assign T202 = {22'h0, T107};
  assign T171 = T37 ? T181 : T172;
  assign T172 = T46 ? T180 : T173;
  assign T173 = T35 ? T203 : T174;
  assign T174 = T178 ? T177 : T175;
  assign T175 = T176 + 9'h100;
  assign T176 = T44[4'h8:1'h0];
  assign T177 = T175 + 9'h1;
  assign T178 = T76[5'h18:5'h18];
  assign T203 = {2'h0, T179};
  assign T179 = T164 ? 7'h6b : 7'h0;
  assign T180 = T162 ? 9'h180 : 9'h17f;
  assign T181 = T40 << 3'h6;
  assign T182 = {T198, T183};
  assign T183 = {T187, T184};
  assign T184 = T186 | T185;
  assign T185 = T115 << 5'h1d;
  assign T186 = 52'h0 - T204;
  assign T204 = {51'h0, T116};
  assign T187 = T197 ? T206 : T188;
  assign T188 = T195 ? T205 : T189;
  assign T189 = T193 ? T192 : T190;
  assign T190 = T191 ? 12'hc00 : 12'he00;
  assign T191 = T117 < 3'h7;
  assign T192 = {4'h8, T196};
  assign T196 = R21[5'h1e:5'h17];
  assign T193 = T117 < 3'h6;
  assign T205 = {1'h0, T194};
  assign T194 = {3'h7, T196};
  assign T195 = T117 < 3'h4;
  assign T206 = {4'h0, T196};
  assign T197 = T117 < 3'h1;
  assign T198 = R21[6'h20:6'h20];
  assign io_out_valid = R199;
  assign T207 = reset ? 1'h0 : R120;

  always @(posedge clk) begin
    if(R120) begin
      R0 <= mux_exc;
    end
    if(io_in_valid) begin
      R9 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      R12 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R29 <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      R92 <= io_in_bits_rm;
    end
    if(reset) begin
      R120 <= 1'h0;
    end else begin
      R120 <= io_in_valid;
    end
    if(R120) begin
      R121 <= mux_data;
    end
    if(reset) begin
      R199 <= 1'h0;
    end else begin
      R199 <= R120;
    end
  end
endmodule

module FPU(input clk, input reset,
    input  io_ctrl_valid,
    output io_ctrl_fcsr_rdy,
    output io_ctrl_nack_mem,
    output io_ctrl_illegal_rm,
    input  io_ctrl_killx,
    input  io_ctrl_killm,
    output[4:0] io_ctrl_dec_cmd,
    output io_ctrl_dec_ldst,
    output io_ctrl_dec_wen,
    output io_ctrl_dec_ren1,
    output io_ctrl_dec_ren2,
    output io_ctrl_dec_ren3,
    output io_ctrl_dec_swap23,
    output io_ctrl_dec_single,
    output io_ctrl_dec_fromint,
    output io_ctrl_dec_toint,
    output io_ctrl_dec_fastpipe,
    output io_ctrl_dec_fma,
    output io_ctrl_dec_round,
    output io_ctrl_sboard_set,
    output io_ctrl_sboard_clr,
    output[4:0] io_ctrl_sboard_clra,
    input [31:0] io_dpath_inst,
    input [63:0] io_dpath_fromint_data,
    input [2:0] io_dpath_fcsr_rm,
    output io_dpath_fcsr_flags_valid,
    output[4:0] io_dpath_fcsr_flags_bits,
    output[63:0] io_dpath_store_data,
    output[63:0] io_dpath_toint_data,
    input  io_dpath_dmem_resp_val,
    input [2:0] io_dpath_dmem_resp_type,
    input [4:0] io_dpath_dmem_resp_tag,
    input [63:0] io_dpath_dmem_resp_data
);

  wire[64:0] req_in3;
  wire[64:0] ex_rs3;
  reg [64:0] regfile [31:0];
  wire[64:0] T120;
  wire[64:0] T121;
  wire[96:0] wdata;
  wire[96:0] T122;
  wire[64:0] T123;
  wire T124;
  wire[1:0] T125;
  wire[1:0] wsrc;
  reg [6:0] winfo_0;
  wire[6:0] T5;
  wire[6:0] T6;
  reg [6:0] winfo_1;
  wire[6:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] memLatencyMask;
  wire[1:0] T11;
  wire T12;
  wire T13;
  reg  mem_ctrl_single;
  wire T14;
  reg  ex_ctrl_single;
  wire T15;
  reg  ex_reg_valid;
  wire T105;
  reg  mem_ctrl_fma;
  wire T16;
  reg  ex_ctrl_fma;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T106;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  reg  mem_ctrl_fromint;
  wire T22;
  reg  ex_ctrl_fromint;
  wire T23;
  wire[1:0] T107;
  reg  mem_ctrl_fastpipe;
  wire T24;
  reg  ex_ctrl_fastpipe;
  wire T25;
  wire T26;
  reg  write_port_busy;
  wire T27;
  wire T28;
  wire T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire[3:0] T35;
  wire[3:0] T108;
  wire[2:0] T36;
  wire T37;
  wire[3:0] T38;
  wire[3:0] T39;
  wire[3:0] T109;
  wire[2:0] T40;
  wire[3:0] T110;
  reg [1:0] wen;
  wire[1:0] T111;
  wire[1:0] T41;
  wire[1:0] T112;
  wire T42;
  wire[1:0] T43;
  wire[1:0] T113;
  wire T44;
  wire T45;
  wire T46;
  wire killm;
  wire T47;
  wire T48;
  wire[2:0] T49;
  wire[2:0] T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T114;
  wire[1:0] T55;
  wire T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T115;
  wire[1:0] T59;
  wire[2:0] T116;
  wire mem_wen;
  wire T60;
  wire T61;
  reg  mem_reg_valid;
  wire T117;
  wire T62;
  wire T63;
  wire T64;
  wire[6:0] mem_winfo;
  wire[4:0] T65;
  reg [31:0] mem_reg_inst;
  wire[31:0] T66;
  reg [31:0] ex_reg_inst;
  wire[31:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T118;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[96:0] T126;
  wire[96:0] T127;
  wire[96:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[4:0] T132;
  wire[4:0] waddr;
  wire[4:0] T93;
  wire[64:0] T133;
  wire[64:0] load_wb_data_recoded;
  wire[64:0] rec_d;
  wire[63:0] T134;
  wire[51:0] T135;
  wire[51:0] T136;
  reg [63:0] load_wb_data;
  wire[63:0] T137;
  wire[51:0] T138;
  wire[126:0] T139;
  wire[5:0] T140;
  wire[5:0] T141;
  wire[5:0] T142;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire[5:0] T146;
  wire[5:0] T147;
  wire[5:0] T148;
  wire[5:0] T149;
  wire[5:0] T150;
  wire[5:0] T151;
  wire[5:0] T152;
  wire[5:0] T153;
  wire[5:0] T154;
  wire[5:0] T155;
  wire[5:0] T156;
  wire[5:0] T157;
  wire[5:0] T158;
  wire[5:0] T159;
  wire[5:0] T160;
  wire[5:0] T161;
  wire[5:0] T162;
  wire[5:0] T163;
  wire[5:0] T164;
  wire[5:0] T165;
  wire[5:0] T166;
  wire[5:0] T167;
  wire[5:0] T168;
  wire[5:0] T169;
  wire[5:0] T170;
  wire[5:0] T171;
  wire[5:0] T172;
  wire[4:0] T173;
  wire[4:0] T174;
  wire[4:0] T175;
  wire[4:0] T176;
  wire[4:0] T177;
  wire[4:0] T178;
  wire[4:0] T179;
  wire[4:0] T180;
  wire[4:0] T181;
  wire[4:0] T182;
  wire[4:0] T183;
  wire[4:0] T184;
  wire[4:0] T185;
  wire[4:0] T186;
  wire[4:0] T187;
  wire[4:0] T188;
  wire[3:0] T189;
  wire[3:0] T190;
  wire[3:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[3:0] T195;
  wire[3:0] T196;
  wire[2:0] T197;
  wire[2:0] T198;
  wire[2:0] T199;
  wire[2:0] T200;
  wire[1:0] T201;
  wire[1:0] T202;
  wire T203;
  wire[63:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire[63:0] T267;
  wire T268;
  wire[10:0] T269;
  wire[11:0] T270;
  wire[11:0] T271;
  wire[9:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire[1:0] T277;
  wire[11:0] T278;
  wire[11:0] T279;
  wire[10:0] T280;
  wire[10:0] T281;
  wire[10:0] T282;
  wire[1:0] T283;
  wire T284;
  wire T285;
  wire T286;
  wire[11:0] T287;
  wire[11:0] T288;
  wire[11:0] T289;
  wire[11:0] T290;
  wire[5:0] T291;
  wire T292;
  wire[64:0] T293;
  wire[32:0] rec_s;
  wire[31:0] T294;
  wire[22:0] T295;
  wire[22:0] T296;
  wire[22:0] T297;
  wire[62:0] T298;
  wire[4:0] T299;
  wire[4:0] T300;
  wire[4:0] T301;
  wire[4:0] T302;
  wire[4:0] T303;
  wire[4:0] T304;
  wire[4:0] T305;
  wire[4:0] T306;
  wire[4:0] T307;
  wire[4:0] T308;
  wire[4:0] T309;
  wire[4:0] T310;
  wire[4:0] T311;
  wire[4:0] T312;
  wire[4:0] T313;
  wire[4:0] T314;
  wire[4:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[3:0] T318;
  wire[3:0] T319;
  wire[3:0] T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[2:0] T324;
  wire[2:0] T325;
  wire[2:0] T326;
  wire[2:0] T327;
  wire[1:0] T328;
  wire[1:0] T329;
  wire T330;
  wire[31:0] T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire[31:0] T362;
  wire T363;
  wire[7:0] T364;
  wire[8:0] T365;
  wire[8:0] T366;
  wire[6:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[1:0] T372;
  wire[8:0] T373;
  wire[8:0] T374;
  wire[7:0] T375;
  wire[7:0] T376;
  wire[7:0] T377;
  wire[1:0] T378;
  wire T379;
  wire T380;
  wire T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire[8:0] T384;
  wire[8:0] T385;
  wire[4:0] T386;
  wire T387;
  reg  load_wb_single;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  reg  load_wb;
  reg [4:0] load_wb_tag;
  wire[4:0] T392;
  reg [4:0] ex_ra3;
  wire[4:0] T393;
  wire[4:0] T394;
  wire[4:0] T395;
  wire T396;
  wire[4:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire[64:0] req_in2;
  wire[64:0] ex_rs2;
  reg [4:0] ex_ra2;
  wire[4:0] T402;
  wire[4:0] T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[64:0] req_in1;
  wire[64:0] ex_rs1;
  reg [4:0] ex_ra1;
  wire[4:0] T408;
  wire[4:0] T409;
  wire[4:0] T410;
  wire T411;
  wire[4:0] T412;
  wire T413;
  wire[1:0] req_typ;
  wire[1:0] T414;
  wire[2:0] req_rm;
  wire[2:0] ex_rm;
  wire[2:0] T99;
  wire T100;
  wire[2:0] T101;
  wire req_round;
  reg  ex_ctrl_round;
  wire T97;
  wire req_fma;
  wire req_fastpipe;
  wire req_toint;
  reg  ex_ctrl_toint;
  wire T87;
  wire req_fromint;
  wire req_single;
  wire req_swap23;
  reg  ex_ctrl_swap23;
  wire T415;
  wire req_ren3;
  reg  ex_ctrl_ren3;
  wire T416;
  wire req_ren2;
  reg  ex_ctrl_ren2;
  wire T417;
  wire req_ren1;
  reg  ex_ctrl_ren1;
  wire T418;
  wire req_wen;
  reg  ex_ctrl_wen;
  wire T419;
  wire req_ldst;
  reg  ex_ctrl_ldst;
  wire T420;
  wire[4:0] req_cmd;
  reg [4:0] ex_ctrl_cmd;
  wire[4:0] T421;
  wire T422;
  wire[64:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[4:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] wexc;
  wire[4:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[4:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire[4:0] T84;
  reg [4:0] wb_toint_exc;
  wire[4:0] T85;
  reg  mem_ctrl_toint;
  wire T86;
  wire wb_toint_valid;
  reg  wb_ctrl_toint;
  wire T88;
  reg  wb_reg_valid;
  wire T119;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T94;
  reg  R95;
  wire T96;
  wire T98;
  wire T102;
  wire fp_inflight;
  wire T103;
  wire T104;
  wire[4:0] fp_decoder_io_sigs_cmd;
  wire fp_decoder_io_sigs_ldst;
  wire fp_decoder_io_sigs_wen;
  wire fp_decoder_io_sigs_ren1;
  wire fp_decoder_io_sigs_ren2;
  wire fp_decoder_io_sigs_ren3;
  wire fp_decoder_io_sigs_swap23;
  wire fp_decoder_io_sigs_single;
  wire fp_decoder_io_sigs_fromint;
  wire fp_decoder_io_sigs_toint;
  wire fp_decoder_io_sigs_fastpipe;
  wire fp_decoder_io_sigs_fma;
  wire fp_decoder_io_sigs_round;
  wire[64:0] ifpu_io_out_bits_data;
  wire[4:0] ifpu_io_out_bits_exc;
  wire[64:0] fpmu_io_out_bits_data;
  wire[4:0] fpmu_io_out_bits_exc;
  wire[64:0] sfma_io_out_bits_data;
  wire[4:0] sfma_io_out_bits_exc;
  wire[64:0] dfma_io_out_bits_data;
  wire[4:0] dfma_io_out_bits_exc;
  wire fpiu_io_out_bits_lt;
  wire[63:0] fpiu_io_out_bits_store;
  wire[63:0] fpiu_io_out_bits_toint;
  wire[4:0] fpiu_io_out_bits_exc;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 32; initvar = initvar+1)
      regfile[initvar] = {3{$random}};
    winfo_0 = {1{$random}};
    winfo_1 = {1{$random}};
    mem_ctrl_single = {1{$random}};
    ex_ctrl_single = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_ctrl_fma = {1{$random}};
    ex_ctrl_fma = {1{$random}};
    mem_ctrl_fromint = {1{$random}};
    ex_ctrl_fromint = {1{$random}};
    mem_ctrl_fastpipe = {1{$random}};
    ex_ctrl_fastpipe = {1{$random}};
    write_port_busy = {1{$random}};
    wen = {1{$random}};
    mem_reg_valid = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    load_wb_data = {2{$random}};
    load_wb_single = {1{$random}};
    load_wb = {1{$random}};
    load_wb_tag = {1{$random}};
    ex_ra3 = {1{$random}};
    ex_ra2 = {1{$random}};
    ex_ra1 = {1{$random}};
    ex_ctrl_round = {1{$random}};
    ex_ctrl_toint = {1{$random}};
    ex_ctrl_swap23 = {1{$random}};
    ex_ctrl_ren3 = {1{$random}};
    ex_ctrl_ren2 = {1{$random}};
    ex_ctrl_ren1 = {1{$random}};
    ex_ctrl_wen = {1{$random}};
    ex_ctrl_ldst = {1{$random}};
    ex_ctrl_cmd = {1{$random}};
    wb_toint_exc = {1{$random}};
    mem_ctrl_toint = {1{$random}};
    wb_ctrl_toint = {1{$random}};
    wb_reg_valid = {1{$random}};
    R95 = {1{$random}};
  end
`endif

  assign req_in3 = ex_rs3;
  assign ex_rs3 = regfile[ex_ra3];
  assign T121 = wdata[7'h40:1'h0];
  assign wdata = T130 ? T126 : T122;
  assign T122 = {32'h0, T123};
  assign T123 = T124 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data;
  assign T124 = T125[1'h0:1'h0];
  assign T125 = wsrc;
  assign wsrc = winfo_0 >> 3'h5;
  assign T5 = T76 ? mem_winfo : T6;
  assign T6 = T64 ? winfo_1 : winfo_0;
  assign T7 = T8 ? mem_winfo : winfo_1;
  assign T8 = mem_wen & T9;
  assign T9 = T26 & T10;
  assign T10 = memLatencyMask[1'h1:1'h1];
  assign memLatencyMask = T18 | T11;
  assign T11 = T12 ? 2'h2 : 2'h0;
  assign T12 = mem_ctrl_fma & T13;
  assign T13 = mem_ctrl_single ^ 1'h1;
  assign T14 = ex_reg_valid ? ex_ctrl_single : mem_ctrl_single;
  assign T15 = io_ctrl_valid ? fp_decoder_io_sigs_single : ex_ctrl_single;
  assign T105 = reset ? 1'h0 : io_ctrl_valid;
  assign T16 = ex_reg_valid ? ex_ctrl_fma : mem_ctrl_fma;
  assign T17 = io_ctrl_valid ? fp_decoder_io_sigs_fma : ex_ctrl_fma;
  assign T18 = T20 | T106;
  assign T106 = {1'h0, T19};
  assign T19 = mem_ctrl_fma & mem_ctrl_single;
  assign T20 = T107 | T21;
  assign T21 = mem_ctrl_fromint ? 2'h2 : 2'h0;
  assign T22 = ex_reg_valid ? ex_ctrl_fromint : mem_ctrl_fromint;
  assign T23 = io_ctrl_valid ? fp_decoder_io_sigs_fromint : ex_ctrl_fromint;
  assign T107 = {1'h0, mem_ctrl_fastpipe};
  assign T24 = ex_reg_valid ? ex_ctrl_fastpipe : mem_ctrl_fastpipe;
  assign T25 = io_ctrl_valid ? fp_decoder_io_sigs_fastpipe : ex_ctrl_fastpipe;
  assign T26 = write_port_busy ^ 1'h1;
  assign T27 = ex_reg_valid ? T28 : write_port_busy;
  assign T28 = T47 | T29;
  assign T29 = T30 != 4'h0;
  assign T30 = T110 & T31;
  assign T31 = T35 | T32;
  assign T32 = T33 ? 4'h8 : 4'h0;
  assign T33 = ex_ctrl_fma & T34;
  assign T34 = ex_ctrl_single ^ 1'h1;
  assign T35 = T38 | T108;
  assign T108 = {1'h0, T36};
  assign T36 = T37 ? 3'h4 : 3'h0;
  assign T37 = ex_ctrl_fma & ex_ctrl_single;
  assign T38 = T109 | T39;
  assign T39 = ex_ctrl_fromint ? 4'h8 : 4'h0;
  assign T109 = {1'h0, T40};
  assign T40 = ex_ctrl_fastpipe ? 3'h4 : 3'h0;
  assign T110 = {2'h0, wen};
  assign T111 = reset ? 2'h0 : T41;
  assign T41 = T45 ? T43 : T112;
  assign T112 = {1'h0, T42};
  assign T42 = wen >> 1'h1;
  assign T43 = T113 | memLatencyMask;
  assign T113 = {1'h0, T44};
  assign T44 = wen >> 1'h1;
  assign T45 = mem_wen & T46;
  assign T46 = killm ^ 1'h1;
  assign killm = io_ctrl_killm | io_ctrl_nack_mem;
  assign T47 = mem_wen & T48;
  assign T48 = T49 != 3'h0;
  assign T49 = T116 & T50;
  assign T50 = T54 | T51;
  assign T51 = T52 ? 3'h4 : 3'h0;
  assign T52 = ex_ctrl_fma & T53;
  assign T53 = ex_ctrl_single ^ 1'h1;
  assign T54 = T57 | T114;
  assign T114 = {1'h0, T55};
  assign T55 = T56 ? 2'h2 : 2'h0;
  assign T56 = ex_ctrl_fma & ex_ctrl_single;
  assign T57 = T115 | T58;
  assign T58 = ex_ctrl_fromint ? 3'h4 : 3'h0;
  assign T115 = {1'h0, T59};
  assign T59 = ex_ctrl_fastpipe ? 2'h2 : 2'h0;
  assign T116 = {1'h0, memLatencyMask};
  assign mem_wen = mem_reg_valid & T60;
  assign T60 = T61 | mem_ctrl_fromint;
  assign T61 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T117 = reset ? 1'h0 : T62;
  assign T62 = ex_reg_valid & T63;
  assign T63 = io_ctrl_killx ^ 1'h1;
  assign T64 = wen[1'h1:1'h1];
  assign mem_winfo = {T68, T65};
  assign T65 = mem_reg_inst[4'hb:3'h7];
  assign T66 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T67 = io_ctrl_valid ? io_dpath_inst : ex_reg_inst;
  assign T68 = T72 | T69;
  assign T69 = T70 ? 2'h3 : 2'h0;
  assign T70 = mem_ctrl_fma & T71;
  assign T71 = mem_ctrl_single ^ 1'h1;
  assign T72 = T118 | T73;
  assign T73 = T74 ? 2'h2 : 2'h0;
  assign T74 = mem_ctrl_fma & mem_ctrl_single;
  assign T118 = {1'h0, T75};
  assign T75 = 1'h0 | mem_ctrl_fromint;
  assign T76 = mem_wen & T77;
  assign T77 = T79 & T78;
  assign T78 = memLatencyMask[1'h0:1'h0];
  assign T79 = write_port_busy ^ 1'h1;
  assign T126 = T129 ? T128 : T127;
  assign T127 = {32'hffffffff, sfma_io_out_bits_data};
  assign T128 = {32'h0, dfma_io_out_bits_data};
  assign T129 = T125[1'h0:1'h0];
  assign T130 = T125[1'h1:1'h1];
  assign T131 = wen[1'h0:1'h0];
  assign T132 = waddr[3'h4:1'h0];
  assign waddr = T93;
  assign T93 = winfo_0[3'h4:1'h0];
  assign load_wb_data_recoded = load_wb_single ? T293 : rec_d;
  assign rec_d = {T292, T134};
  assign T134 = {T270, T135};
  assign T135 = T268 ? T138 : T136;
  assign T136 = load_wb_data[6'h33:1'h0];
  assign T137 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_data : load_wb_data;
  assign T138 = T139[6'h3e:4'hb];
  assign T139 = T267 << T140;
  assign T140 = ~ T141;
  assign T141 = T266 ? 6'h3f : T142;
  assign T142 = T265 ? 6'h3e : T143;
  assign T143 = T264 ? 6'h3d : T144;
  assign T144 = T263 ? 6'h3c : T145;
  assign T145 = T262 ? 6'h3b : T146;
  assign T146 = T261 ? 6'h3a : T147;
  assign T147 = T260 ? 6'h39 : T148;
  assign T148 = T259 ? 6'h38 : T149;
  assign T149 = T258 ? 6'h37 : T150;
  assign T150 = T257 ? 6'h36 : T151;
  assign T151 = T256 ? 6'h35 : T152;
  assign T152 = T255 ? 6'h34 : T153;
  assign T153 = T254 ? 6'h33 : T154;
  assign T154 = T253 ? 6'h32 : T155;
  assign T155 = T252 ? 6'h31 : T156;
  assign T156 = T251 ? 6'h30 : T157;
  assign T157 = T250 ? 6'h2f : T158;
  assign T158 = T249 ? 6'h2e : T159;
  assign T159 = T248 ? 6'h2d : T160;
  assign T160 = T247 ? 6'h2c : T161;
  assign T161 = T246 ? 6'h2b : T162;
  assign T162 = T245 ? 6'h2a : T163;
  assign T163 = T244 ? 6'h29 : T164;
  assign T164 = T243 ? 6'h28 : T165;
  assign T165 = T242 ? 6'h27 : T166;
  assign T166 = T241 ? 6'h26 : T167;
  assign T167 = T240 ? 6'h25 : T168;
  assign T168 = T239 ? 6'h24 : T169;
  assign T169 = T238 ? 6'h23 : T170;
  assign T170 = T237 ? 6'h22 : T171;
  assign T171 = T236 ? 6'h21 : T172;
  assign T172 = T235 ? 6'h20 : T173;
  assign T173 = T234 ? 5'h1f : T174;
  assign T174 = T233 ? 5'h1e : T175;
  assign T175 = T232 ? 5'h1d : T176;
  assign T176 = T231 ? 5'h1c : T177;
  assign T177 = T230 ? 5'h1b : T178;
  assign T178 = T229 ? 5'h1a : T179;
  assign T179 = T228 ? 5'h19 : T180;
  assign T180 = T227 ? 5'h18 : T181;
  assign T181 = T226 ? 5'h17 : T182;
  assign T182 = T225 ? 5'h16 : T183;
  assign T183 = T224 ? 5'h15 : T184;
  assign T184 = T223 ? 5'h14 : T185;
  assign T185 = T222 ? 5'h13 : T186;
  assign T186 = T221 ? 5'h12 : T187;
  assign T187 = T220 ? 5'h11 : T188;
  assign T188 = T219 ? 5'h10 : T189;
  assign T189 = T218 ? 4'hf : T190;
  assign T190 = T217 ? 4'he : T191;
  assign T191 = T216 ? 4'hd : T192;
  assign T192 = T215 ? 4'hc : T193;
  assign T193 = T214 ? 4'hb : T194;
  assign T194 = T213 ? 4'ha : T195;
  assign T195 = T212 ? 4'h9 : T196;
  assign T196 = T211 ? 4'h8 : T197;
  assign T197 = T210 ? 3'h7 : T198;
  assign T198 = T209 ? 3'h6 : T199;
  assign T199 = T208 ? 3'h5 : T200;
  assign T200 = T207 ? 3'h4 : T201;
  assign T201 = T206 ? 2'h3 : T202;
  assign T202 = T205 ? 2'h2 : T203;
  assign T203 = T204[1'h1:1'h1];
  assign T204 = T267[6'h3f:1'h0];
  assign T205 = T204[2'h2:2'h2];
  assign T206 = T204[2'h3:2'h3];
  assign T207 = T204[3'h4:3'h4];
  assign T208 = T204[3'h5:3'h5];
  assign T209 = T204[3'h6:3'h6];
  assign T210 = T204[3'h7:3'h7];
  assign T211 = T204[4'h8:4'h8];
  assign T212 = T204[4'h9:4'h9];
  assign T213 = T204[4'ha:4'ha];
  assign T214 = T204[4'hb:4'hb];
  assign T215 = T204[4'hc:4'hc];
  assign T216 = T204[4'hd:4'hd];
  assign T217 = T204[4'he:4'he];
  assign T218 = T204[4'hf:4'hf];
  assign T219 = T204[5'h10:5'h10];
  assign T220 = T204[5'h11:5'h11];
  assign T221 = T204[5'h12:5'h12];
  assign T222 = T204[5'h13:5'h13];
  assign T223 = T204[5'h14:5'h14];
  assign T224 = T204[5'h15:5'h15];
  assign T225 = T204[5'h16:5'h16];
  assign T226 = T204[5'h17:5'h17];
  assign T227 = T204[5'h18:5'h18];
  assign T228 = T204[5'h19:5'h19];
  assign T229 = T204[5'h1a:5'h1a];
  assign T230 = T204[5'h1b:5'h1b];
  assign T231 = T204[5'h1c:5'h1c];
  assign T232 = T204[5'h1d:5'h1d];
  assign T233 = T204[5'h1e:5'h1e];
  assign T234 = T204[5'h1f:5'h1f];
  assign T235 = T204[6'h20:6'h20];
  assign T236 = T204[6'h21:6'h21];
  assign T237 = T204[6'h22:6'h22];
  assign T238 = T204[6'h23:6'h23];
  assign T239 = T204[6'h24:6'h24];
  assign T240 = T204[6'h25:6'h25];
  assign T241 = T204[6'h26:6'h26];
  assign T242 = T204[6'h27:6'h27];
  assign T243 = T204[6'h28:6'h28];
  assign T244 = T204[6'h29:6'h29];
  assign T245 = T204[6'h2a:6'h2a];
  assign T246 = T204[6'h2b:6'h2b];
  assign T247 = T204[6'h2c:6'h2c];
  assign T248 = T204[6'h2d:6'h2d];
  assign T249 = T204[6'h2e:6'h2e];
  assign T250 = T204[6'h2f:6'h2f];
  assign T251 = T204[6'h30:6'h30];
  assign T252 = T204[6'h31:6'h31];
  assign T253 = T204[6'h32:6'h32];
  assign T254 = T204[6'h33:6'h33];
  assign T255 = T204[6'h34:6'h34];
  assign T256 = T204[6'h35:6'h35];
  assign T257 = T204[6'h36:6'h36];
  assign T258 = T204[6'h37:6'h37];
  assign T259 = T204[6'h38:6'h38];
  assign T260 = T204[6'h39:6'h39];
  assign T261 = T204[6'h3a:6'h3a];
  assign T262 = T204[6'h3b:6'h3b];
  assign T263 = T204[6'h3c:6'h3c];
  assign T264 = T204[6'h3d:6'h3d];
  assign T265 = T204[6'h3e:6'h3e];
  assign T266 = T204[6'h3f:6'h3f];
  assign T267 = T136 << 4'hc;
  assign T268 = T269 == 11'h0;
  assign T269 = load_wb_data[6'h3e:6'h34];
  assign T270 = T278 | T271;
  assign T271 = {2'h0, T272};
  assign T272 = T273 << 4'h9;
  assign T273 = T276 & T274;
  assign T274 = T275 ^ 1'h1;
  assign T275 = T136 == 52'h0;
  assign T276 = T277 == 2'h3;
  assign T277 = T278[4'hb:4'ha];
  assign T278 = T287 + T279;
  assign T279 = {1'h0, T280};
  assign T280 = T286 ? 11'h0 : T281;
  assign T281 = 11'h400 | T282;
  assign T282 = {9'h0, T283};
  assign T283 = T284 ? 2'h2 : 2'h1;
  assign T284 = T268 & T285;
  assign T285 = T275 ^ 1'h1;
  assign T286 = T268 & T275;
  assign T287 = T268 ? T289 : T288;
  assign T288 = {1'h0, T269};
  assign T289 = T275 ? 12'h0 : T290;
  assign T290 = {6'h3f, T291};
  assign T291 = ~ T140;
  assign T292 = load_wb_data[6'h3f:6'h3f];
  assign T293 = {32'hffffffff, rec_s};
  assign rec_s = {T387, T294};
  assign T294 = {T365, T295};
  assign T295 = T363 ? T297 : T296;
  assign T296 = load_wb_data[5'h16:1'h0];
  assign T297 = T298[5'h1e:4'h8];
  assign T298 = T362 << T299;
  assign T299 = ~ T300;
  assign T300 = T361 ? 5'h1f : T301;
  assign T301 = T360 ? 5'h1e : T302;
  assign T302 = T359 ? 5'h1d : T303;
  assign T303 = T358 ? 5'h1c : T304;
  assign T304 = T357 ? 5'h1b : T305;
  assign T305 = T356 ? 5'h1a : T306;
  assign T306 = T355 ? 5'h19 : T307;
  assign T307 = T354 ? 5'h18 : T308;
  assign T308 = T353 ? 5'h17 : T309;
  assign T309 = T352 ? 5'h16 : T310;
  assign T310 = T351 ? 5'h15 : T311;
  assign T311 = T350 ? 5'h14 : T312;
  assign T312 = T349 ? 5'h13 : T313;
  assign T313 = T348 ? 5'h12 : T314;
  assign T314 = T347 ? 5'h11 : T315;
  assign T315 = T346 ? 5'h10 : T316;
  assign T316 = T345 ? 4'hf : T317;
  assign T317 = T344 ? 4'he : T318;
  assign T318 = T343 ? 4'hd : T319;
  assign T319 = T342 ? 4'hc : T320;
  assign T320 = T341 ? 4'hb : T321;
  assign T321 = T340 ? 4'ha : T322;
  assign T322 = T339 ? 4'h9 : T323;
  assign T323 = T338 ? 4'h8 : T324;
  assign T324 = T337 ? 3'h7 : T325;
  assign T325 = T336 ? 3'h6 : T326;
  assign T326 = T335 ? 3'h5 : T327;
  assign T327 = T334 ? 3'h4 : T328;
  assign T328 = T333 ? 2'h3 : T329;
  assign T329 = T332 ? 2'h2 : T330;
  assign T330 = T331[1'h1:1'h1];
  assign T331 = T362[5'h1f:1'h0];
  assign T332 = T331[2'h2:2'h2];
  assign T333 = T331[2'h3:2'h3];
  assign T334 = T331[3'h4:3'h4];
  assign T335 = T331[3'h5:3'h5];
  assign T336 = T331[3'h6:3'h6];
  assign T337 = T331[3'h7:3'h7];
  assign T338 = T331[4'h8:4'h8];
  assign T339 = T331[4'h9:4'h9];
  assign T340 = T331[4'ha:4'ha];
  assign T341 = T331[4'hb:4'hb];
  assign T342 = T331[4'hc:4'hc];
  assign T343 = T331[4'hd:4'hd];
  assign T344 = T331[4'he:4'he];
  assign T345 = T331[4'hf:4'hf];
  assign T346 = T331[5'h10:5'h10];
  assign T347 = T331[5'h11:5'h11];
  assign T348 = T331[5'h12:5'h12];
  assign T349 = T331[5'h13:5'h13];
  assign T350 = T331[5'h14:5'h14];
  assign T351 = T331[5'h15:5'h15];
  assign T352 = T331[5'h16:5'h16];
  assign T353 = T331[5'h17:5'h17];
  assign T354 = T331[5'h18:5'h18];
  assign T355 = T331[5'h19:5'h19];
  assign T356 = T331[5'h1a:5'h1a];
  assign T357 = T331[5'h1b:5'h1b];
  assign T358 = T331[5'h1c:5'h1c];
  assign T359 = T331[5'h1d:5'h1d];
  assign T360 = T331[5'h1e:5'h1e];
  assign T361 = T331[5'h1f:5'h1f];
  assign T362 = T296 << 4'h9;
  assign T363 = T364 == 8'h0;
  assign T364 = load_wb_data[5'h1e:5'h17];
  assign T365 = T373 | T366;
  assign T366 = {2'h0, T367};
  assign T367 = T368 << 3'h6;
  assign T368 = T371 & T369;
  assign T369 = T370 ^ 1'h1;
  assign T370 = T296 == 23'h0;
  assign T371 = T372 == 2'h3;
  assign T372 = T373[4'h8:3'h7];
  assign T373 = T382 + T374;
  assign T374 = {1'h0, T375};
  assign T375 = T381 ? 8'h0 : T376;
  assign T376 = 8'h80 | T377;
  assign T377 = {6'h0, T378};
  assign T378 = T379 ? 2'h2 : 2'h1;
  assign T379 = T363 & T380;
  assign T380 = T370 ^ 1'h1;
  assign T381 = T363 & T370;
  assign T382 = T363 ? T384 : T383;
  assign T383 = {1'h0, T364};
  assign T384 = T370 ? 9'h0 : T385;
  assign T385 = {4'hf, T386};
  assign T386 = ~ T299;
  assign T387 = load_wb_data[5'h1f:5'h1f];
  assign T388 = io_dpath_dmem_resp_val ? T389 : load_wb_single;
  assign T389 = T391 | T390;
  assign T390 = io_dpath_dmem_resp_type == 3'h6;
  assign T391 = io_dpath_dmem_resp_type == 3'h2;
  assign T392 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_tag : load_wb_tag;
  assign T393 = T398 ? T397 : T394;
  assign T394 = T396 ? T395 : ex_ra3;
  assign T395 = io_dpath_inst[5'h1f:5'h1b];
  assign T396 = io_ctrl_valid & fp_decoder_io_sigs_ren3;
  assign T397 = io_dpath_inst[5'h18:5'h14];
  assign T398 = T401 & T399;
  assign T399 = T400 & fp_decoder_io_sigs_swap23;
  assign T400 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign T401 = io_ctrl_valid & fp_decoder_io_sigs_ren2;
  assign req_in2 = ex_rs2;
  assign ex_rs2 = regfile[ex_ra2];
  assign T402 = T404 ? T403 : ex_ra2;
  assign T403 = io_dpath_inst[5'h18:5'h14];
  assign T404 = T401 & T405;
  assign T405 = T407 & T406;
  assign T406 = fp_decoder_io_sigs_swap23 ^ 1'h1;
  assign T407 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign req_in1 = ex_rs1;
  assign ex_rs1 = regfile[ex_ra1];
  assign T408 = T413 ? T412 : T409;
  assign T409 = T411 ? T410 : ex_ra1;
  assign T410 = io_dpath_inst[5'h13:4'hf];
  assign T411 = io_ctrl_valid & fp_decoder_io_sigs_ren1;
  assign T412 = io_dpath_inst[5'h18:5'h14];
  assign T413 = T401 & fp_decoder_io_sigs_ldst;
  assign req_typ = T414;
  assign T414 = ex_reg_inst[5'h15:5'h14];
  assign req_rm = ex_rm;
  assign ex_rm = T100 ? io_dpath_fcsr_rm : T99;
  assign T99 = ex_reg_inst[4'he:4'hc];
  assign T100 = T101 == 3'h7;
  assign T101 = ex_reg_inst[4'he:4'hc];
  assign req_round = ex_ctrl_round;
  assign T97 = io_ctrl_valid ? fp_decoder_io_sigs_round : ex_ctrl_round;
  assign req_fma = ex_ctrl_fma;
  assign req_fastpipe = ex_ctrl_fastpipe;
  assign req_toint = ex_ctrl_toint;
  assign T87 = io_ctrl_valid ? fp_decoder_io_sigs_toint : ex_ctrl_toint;
  assign req_fromint = ex_ctrl_fromint;
  assign req_single = ex_ctrl_single;
  assign req_swap23 = ex_ctrl_swap23;
  assign T415 = io_ctrl_valid ? fp_decoder_io_sigs_swap23 : ex_ctrl_swap23;
  assign req_ren3 = ex_ctrl_ren3;
  assign T416 = io_ctrl_valid ? fp_decoder_io_sigs_ren3 : ex_ctrl_ren3;
  assign req_ren2 = ex_ctrl_ren2;
  assign T417 = io_ctrl_valid ? fp_decoder_io_sigs_ren2 : ex_ctrl_ren2;
  assign req_ren1 = ex_ctrl_ren1;
  assign T418 = io_ctrl_valid ? fp_decoder_io_sigs_ren1 : ex_ctrl_ren1;
  assign req_wen = ex_ctrl_wen;
  assign T419 = io_ctrl_valid ? fp_decoder_io_sigs_wen : ex_ctrl_wen;
  assign req_ldst = ex_ctrl_ldst;
  assign T420 = io_ctrl_valid ? fp_decoder_io_sigs_ldst : ex_ctrl_ldst;
  assign req_cmd = ex_ctrl_cmd;
  assign T421 = io_ctrl_valid ? fp_decoder_io_sigs_cmd : ex_ctrl_cmd;
  assign T422 = ex_reg_valid & ex_ctrl_fastpipe;
  assign T423 = {1'h0, io_dpath_fromint_data};
  assign T424 = ex_reg_valid & ex_ctrl_fromint;
  assign T425 = ex_reg_valid & T426;
  assign T426 = ex_ctrl_toint | T427;
  assign T427 = T428 == 5'h5;
  assign T428 = ex_ctrl_cmd & 5'hd;
  assign T429 = T431 & T430;
  assign T430 = ex_ctrl_single ^ 1'h1;
  assign T431 = ex_reg_valid & ex_ctrl_fma;
  assign T432 = T433 & ex_ctrl_single;
  assign T433 = ex_reg_valid & ex_ctrl_fma;
  assign io_dpath_toint_data = fpiu_io_out_bits_toint;
  assign io_dpath_store_data = fpiu_io_out_bits_store;
  assign io_dpath_fcsr_flags_bits = T0;
  assign T0 = T84 | T1;
  assign T1 = T83 ? wexc : 5'h0;
  assign wexc = T82 ? T80 : T2;
  assign T2 = T3 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = wsrc;
  assign T80 = T81 ? dfma_io_out_bits_exc : sfma_io_out_bits_exc;
  assign T81 = T4[1'h0:1'h0];
  assign T82 = T4[1'h1:1'h1];
  assign T83 = wen[1'h0:1'h0];
  assign T84 = wb_toint_valid ? wb_toint_exc : 5'h0;
  assign T85 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign T86 = ex_reg_valid ? ex_ctrl_toint : mem_ctrl_toint;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign T88 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign T119 = reset ? 1'h0 : T89;
  assign T89 = mem_reg_valid & T90;
  assign T90 = killm ^ 1'h1;
  assign io_dpath_fcsr_flags_valid = T91;
  assign T91 = wb_toint_valid | T92;
  assign T92 = wen[1'h0:1'h0];
  assign io_ctrl_sboard_clra = waddr;
  assign io_ctrl_sboard_clr = 1'h0;
  assign io_ctrl_sboard_set = T94;
  assign T94 = wb_reg_valid & R95;
  assign io_ctrl_dec_round = fp_decoder_io_sigs_round;
  assign io_ctrl_dec_fma = fp_decoder_io_sigs_fma;
  assign io_ctrl_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_ctrl_dec_toint = fp_decoder_io_sigs_toint;
  assign io_ctrl_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_ctrl_dec_single = fp_decoder_io_sigs_single;
  assign io_ctrl_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_ctrl_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_ctrl_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_ctrl_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_ctrl_dec_wen = fp_decoder_io_sigs_wen;
  assign io_ctrl_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_ctrl_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_ctrl_illegal_rm = T96;
  assign T96 = T98 & ex_ctrl_round;
  assign T98 = ex_rm[2'h2:2'h2];
  assign io_ctrl_nack_mem = write_port_busy;
  assign io_ctrl_fcsr_rdy = T102;
  assign T102 = fp_inflight ^ 1'h1;
  assign fp_inflight = T104 | T103;
  assign T103 = wen != 2'h0;
  assign T104 = wb_reg_valid & wb_ctrl_toint;
  FPUDecoder fp_decoder(
       .io_inst( io_dpath_inst ),
       .io_sigs_cmd( fp_decoder_io_sigs_cmd ),
       .io_sigs_ldst( fp_decoder_io_sigs_ldst ),
       .io_sigs_wen( fp_decoder_io_sigs_wen ),
       .io_sigs_ren1( fp_decoder_io_sigs_ren1 ),
       .io_sigs_ren2( fp_decoder_io_sigs_ren2 ),
       .io_sigs_ren3( fp_decoder_io_sigs_ren3 ),
       .io_sigs_swap23( fp_decoder_io_sigs_swap23 ),
       .io_sigs_single( fp_decoder_io_sigs_single ),
       .io_sigs_fromint( fp_decoder_io_sigs_fromint ),
       .io_sigs_toint( fp_decoder_io_sigs_toint ),
       .io_sigs_fastpipe( fp_decoder_io_sigs_fastpipe ),
       .io_sigs_fma( fp_decoder_io_sigs_fma ),
       .io_sigs_round( fp_decoder_io_sigs_round )
  );
  FPUFMAPipe_0 sfma(.clk(clk), .reset(reset),
       .io_in_valid( T432 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( sfma_io_out_bits_data ),
       .io_out_bits_exc( sfma_io_out_bits_exc )
  );
  FPUFMAPipe_1 dfma(.clk(clk), .reset(reset),
       .io_in_valid( T429 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( dfma_io_out_bits_data ),
       .io_out_bits_exc( dfma_io_out_bits_exc )
  );
  FPToInt fpiu(.clk(clk),
       .io_in_valid( T425 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_lt( fpiu_io_out_bits_lt ),
       .io_out_bits_store( fpiu_io_out_bits_store ),
       .io_out_bits_toint( fpiu_io_out_bits_toint ),
       .io_out_bits_exc( fpiu_io_out_bits_exc )
  );
  IntToFP ifpu(.clk(clk), .reset(reset),
       .io_in_valid( T424 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( T423 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( ifpu_io_out_bits_data ),
       .io_out_bits_exc( ifpu_io_out_bits_exc )
  );
  FPToFP fpmu(.clk(clk), .reset(reset),
       .io_in_valid( T422 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( fpmu_io_out_bits_data ),
       .io_out_bits_exc( fpmu_io_out_bits_exc ),
       .io_lt( fpiu_io_out_bits_lt )
  );

  always @(posedge clk) begin
    if (T131)
      regfile[T132] <= T121;
    if(T76) begin
      winfo_0 <= mem_winfo;
    end else if(T64) begin
      winfo_0 <= winfo_1;
    end
    if(T8) begin
      winfo_1 <= mem_winfo;
    end
    if(ex_reg_valid) begin
      mem_ctrl_single <= ex_ctrl_single;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_single <= fp_decoder_io_sigs_single;
    end
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_ctrl_valid;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fma <= ex_ctrl_fma;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fromint <= ex_ctrl_fromint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_ctrl_fastpipe;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if(ex_reg_valid) begin
      write_port_busy <= T28;
    end
    if(reset) begin
      wen <= 2'h0;
    end else if(T45) begin
      wen <= T43;
    end else begin
      wen <= T112;
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T62;
    end
    if(ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(io_ctrl_valid) begin
      ex_reg_inst <= io_dpath_inst;
    end
    if (load_wb)
      regfile[load_wb_tag] <= load_wb_data_recoded;
    if(io_dpath_dmem_resp_val) begin
      load_wb_data <= io_dpath_dmem_resp_data;
    end
    if(io_dpath_dmem_resp_val) begin
      load_wb_single <= T389;
    end
    load_wb <= io_dpath_dmem_resp_val;
    if(io_dpath_dmem_resp_val) begin
      load_wb_tag <= io_dpath_dmem_resp_tag;
    end
    if(T398) begin
      ex_ra3 <= T397;
    end else if(T396) begin
      ex_ra3 <= T395;
    end
    if(T404) begin
      ex_ra2 <= T403;
    end
    if(T413) begin
      ex_ra1 <= T412;
    end else if(T411) begin
      ex_ra1 <= T410;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_round <= fp_decoder_io_sigs_round;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren1 <= fp_decoder_io_sigs_ren1;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_wen <= fp_decoder_io_sigs_wen;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ldst <= fp_decoder_io_sigs_ldst;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_cmd <= fp_decoder_io_sigs_cmd;
    end
    if(mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if(ex_reg_valid) begin
      mem_ctrl_toint <= ex_ctrl_toint;
    end
    if(mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T89;
    end
    R95 <= 1'h0;
  end
endmodule

module Core(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[43:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_mispredict,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready
);

  wire[2:0] ctrl_io_dpath_sel_pc;
  wire ctrl_io_dpath_killd;
  wire ctrl_io_dpath_ren_1;
  wire ctrl_io_dpath_ren_0;
  wire[2:0] ctrl_io_dpath_sel_alu2;
  wire[1:0] ctrl_io_dpath_sel_alu1;
  wire[2:0] ctrl_io_dpath_sel_imm;
  wire ctrl_io_dpath_fn_dw;
  wire[3:0] ctrl_io_dpath_fn_alu;
  wire ctrl_io_dpath_div_mul_val;
  wire ctrl_io_dpath_div_mul_kill;
  wire[2:0] ctrl_io_dpath_csr;
  wire ctrl_io_dpath_sret;
  wire ctrl_io_dpath_mem_load;
  wire ctrl_io_dpath_wb_load;
  wire ctrl_io_dpath_ex_fp_val;
  wire ctrl_io_dpath_mem_fp_val;
  wire ctrl_io_dpath_ex_wen;
  wire ctrl_io_dpath_ex_valid;
  wire ctrl_io_dpath_mem_jalr;
  wire ctrl_io_dpath_mem_branch;
  wire ctrl_io_dpath_mem_wen;
  wire ctrl_io_dpath_wb_wen;
  wire[2:0] ctrl_io_dpath_ex_mem_type;
  wire ctrl_io_dpath_ex_rs2_val;
  wire ctrl_io_dpath_ex_rocc_val;
  wire ctrl_io_dpath_mem_rocc_val;
  wire ctrl_io_dpath_bypass_1;
  wire ctrl_io_dpath_bypass_0;
  wire[1:0] ctrl_io_dpath_bypass_src_1;
  wire[1:0] ctrl_io_dpath_bypass_src_0;
  wire ctrl_io_dpath_ll_ready;
  wire ctrl_io_dpath_retire;
  wire ctrl_io_dpath_exception;
  wire[63:0] ctrl_io_dpath_cause;
  wire ctrl_io_dpath_badvaddr_wen;
  wire ctrl_io_imem_req_valid;
  wire ctrl_io_imem_resp_ready;
  wire ctrl_io_imem_btb_update_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  wire[42:0] ctrl_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire ctrl_io_imem_btb_update_bits_taken;
  wire ctrl_io_imem_btb_update_bits_isJump;
  wire ctrl_io_imem_btb_update_bits_isCall;
  wire ctrl_io_imem_btb_update_bits_isReturn;
  wire ctrl_io_imem_btb_update_bits_mispredict;
  wire ctrl_io_imem_invalidate;
  wire ctrl_io_dmem_req_valid;
  wire ctrl_io_dmem_req_bits_kill;
  wire[2:0] ctrl_io_dmem_req_bits_typ;
  wire ctrl_io_dmem_req_bits_phys;
  wire[4:0] ctrl_io_dmem_req_bits_cmd;
  wire ctrl_io_fpu_valid;
  wire ctrl_io_fpu_killx;
  wire ctrl_io_fpu_killm;
  wire ctrl_io_rocc_cmd_valid;
  wire ctrl_io_rocc_s;
  wire ctrl_io_rocc_exception;
  wire dpath_io_host_pcr_req_ready;
  wire dpath_io_host_pcr_rep_valid;
  wire[63:0] dpath_io_host_pcr_rep_bits;
  wire dpath_io_host_ipi_req_valid;
  wire dpath_io_host_ipi_req_bits;
  wire dpath_io_host_ipi_rep_ready;
  wire dpath_io_host_debug_stats_pcr;
  wire[31:0] dpath_io_ctrl_inst;
  wire dpath_io_ctrl_mem_br_taken;
  wire dpath_io_ctrl_mem_misprediction;
  wire dpath_io_ctrl_div_mul_rdy;
  wire dpath_io_ctrl_ll_wen;
  wire[4:0] dpath_io_ctrl_ll_waddr;
  wire[4:0] dpath_io_ctrl_ex_waddr;
  wire dpath_io_ctrl_mem_rs1_ra;
  wire[4:0] dpath_io_ctrl_mem_waddr;
  wire[4:0] dpath_io_ctrl_wb_waddr;
  wire[7:0] dpath_io_ctrl_status_ip;
  wire[7:0] dpath_io_ctrl_status_im;
  wire[6:0] dpath_io_ctrl_status_zero;
  wire dpath_io_ctrl_status_er;
  wire dpath_io_ctrl_status_vm;
  wire dpath_io_ctrl_status_s64;
  wire dpath_io_ctrl_status_u64;
  wire dpath_io_ctrl_status_ef;
  wire dpath_io_ctrl_status_pei;
  wire dpath_io_ctrl_status_ei;
  wire dpath_io_ctrl_status_ps;
  wire dpath_io_ctrl_status_s;
  wire dpath_io_ctrl_fp_sboard_clr;
  wire[4:0] dpath_io_ctrl_fp_sboard_clra;
  wire dpath_io_ctrl_csr_replay;
  wire[43:0] dpath_io_dmem_req_bits_addr;
  wire[63:0] dpath_io_dmem_req_bits_data;
  wire[7:0] dpath_io_dmem_req_bits_tag;
  wire[31:0] dpath_io_ptw_ptbr;
  wire dpath_io_ptw_invalidate;
  wire dpath_io_ptw_sret;
  wire[7:0] dpath_io_ptw_status_ip;
  wire[7:0] dpath_io_ptw_status_im;
  wire[6:0] dpath_io_ptw_status_zero;
  wire dpath_io_ptw_status_er;
  wire dpath_io_ptw_status_vm;
  wire dpath_io_ptw_status_s64;
  wire dpath_io_ptw_status_u64;
  wire dpath_io_ptw_status_ef;
  wire dpath_io_ptw_status_pei;
  wire dpath_io_ptw_status_ei;
  wire dpath_io_ptw_status_ps;
  wire dpath_io_ptw_status_s;
  wire[43:0] dpath_io_imem_req_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_target;
  wire[42:0] dpath_io_imem_btb_update_bits_returnAddr;
  wire[31:0] dpath_io_fpu_inst;
  wire[63:0] dpath_io_fpu_fromint_data;
  wire[2:0] dpath_io_fpu_fcsr_rm;
  wire dpath_io_fpu_dmem_resp_val;
  wire[2:0] dpath_io_fpu_dmem_resp_type;
  wire[4:0] dpath_io_fpu_dmem_resp_tag;
  wire[63:0] dpath_io_fpu_dmem_resp_data;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_funct;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs1;
  wire dpath_io_rocc_cmd_bits_inst_xd;
  wire dpath_io_rocc_cmd_bits_inst_xs1;
  wire dpath_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rd;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] dpath_io_rocc_cmd_bits_rs1;
  wire[63:0] dpath_io_rocc_cmd_bits_rs2;
  wire dpath_io_temac_rx_axis_fifo_tready;
  wire[7:0] dpath_io_temac_tx_axis_fifo_tdata;
  wire dpath_io_temac_tx_axis_fifo_tvalid;
  wire dpath_io_temac_tx_axis_fifo_tlast;
  wire[11:0] dpath_io_temac_s_axi_awaddr;
  wire dpath_io_temac_s_axi_awvalid;
  wire[31:0] dpath_io_temac_s_axi_wdata;
  wire dpath_io_temac_s_axi_wvalid;
  wire dpath_io_temac_s_axi_bready;
  wire[11:0] dpath_io_temac_s_axi_araddr;
  wire dpath_io_temac_s_axi_arvalid;
  wire dpath_io_temac_s_axi_rready;
  wire FPU_io_ctrl_fcsr_rdy;
  wire FPU_io_ctrl_nack_mem;
  wire FPU_io_ctrl_illegal_rm;
  wire[4:0] FPU_io_ctrl_dec_cmd;
  wire FPU_io_ctrl_dec_ldst;
  wire FPU_io_ctrl_dec_wen;
  wire FPU_io_ctrl_dec_ren1;
  wire FPU_io_ctrl_dec_ren2;
  wire FPU_io_ctrl_dec_ren3;
  wire FPU_io_ctrl_dec_swap23;
  wire FPU_io_ctrl_dec_single;
  wire FPU_io_ctrl_dec_fromint;
  wire FPU_io_ctrl_dec_toint;
  wire FPU_io_ctrl_dec_fastpipe;
  wire FPU_io_ctrl_dec_fma;
  wire FPU_io_ctrl_dec_round;
  wire FPU_io_ctrl_sboard_set;
  wire FPU_io_ctrl_sboard_clr;
  wire[4:0] FPU_io_ctrl_sboard_clra;
  wire FPU_io_dpath_fcsr_flags_valid;
  wire[4:0] FPU_io_dpath_fcsr_flags_bits;
  wire[63:0] FPU_io_dpath_store_data;
  wire[63:0] FPU_io_dpath_toint_data;


  assign io_temac_s_axi_rready = dpath_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = dpath_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = dpath_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = dpath_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = dpath_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = dpath_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = dpath_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = dpath_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = dpath_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = dpath_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = dpath_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = dpath_io_temac_rx_axis_fifo_tready;
  assign io_rocc_exception = ctrl_io_rocc_exception;
  assign io_rocc_s = ctrl_io_rocc_s;
  assign io_rocc_cmd_bits_rs2 = dpath_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = dpath_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = dpath_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = dpath_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = dpath_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = dpath_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = dpath_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = dpath_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = dpath_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = dpath_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = ctrl_io_rocc_cmd_valid;
  assign io_ptw_status_s = dpath_io_ptw_status_s;
  assign io_ptw_status_ps = dpath_io_ptw_status_ps;
  assign io_ptw_status_ei = dpath_io_ptw_status_ei;
  assign io_ptw_status_pei = dpath_io_ptw_status_pei;
  assign io_ptw_status_ef = dpath_io_ptw_status_ef;
  assign io_ptw_status_u64 = dpath_io_ptw_status_u64;
  assign io_ptw_status_s64 = dpath_io_ptw_status_s64;
  assign io_ptw_status_vm = dpath_io_ptw_status_vm;
  assign io_ptw_status_er = dpath_io_ptw_status_er;
  assign io_ptw_status_zero = dpath_io_ptw_status_zero;
  assign io_ptw_status_im = dpath_io_ptw_status_im;
  assign io_ptw_status_ip = dpath_io_ptw_status_ip;
  assign io_ptw_sret = dpath_io_ptw_sret;
  assign io_ptw_invalidate = dpath_io_ptw_invalidate;
  assign io_ptw_ptbr = dpath_io_ptw_ptbr;
  assign io_dmem_req_bits_cmd = ctrl_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_tag = dpath_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_phys = ctrl_io_dmem_req_bits_phys;
  assign io_dmem_req_bits_typ = ctrl_io_dmem_req_bits_typ;
  assign io_dmem_req_bits_kill = ctrl_io_dmem_req_bits_kill;
  assign io_dmem_req_valid = ctrl_io_dmem_req_valid;
  assign io_imem_invalidate = ctrl_io_imem_invalidate;
  assign io_imem_btb_update_bits_mispredict = ctrl_io_imem_btb_update_bits_mispredict;
  assign io_imem_btb_update_bits_isReturn = ctrl_io_imem_btb_update_bits_isReturn;
  assign io_imem_btb_update_bits_isCall = ctrl_io_imem_btb_update_bits_isCall;
  assign io_imem_btb_update_bits_isJump = ctrl_io_imem_btb_update_bits_isJump;
  assign io_imem_btb_update_bits_taken = ctrl_io_imem_btb_update_bits_taken;
  assign io_imem_btb_update_bits_returnAddr = dpath_io_imem_btb_update_bits_returnAddr;
  assign io_imem_btb_update_bits_target = dpath_io_imem_btb_update_bits_target;
  assign io_imem_btb_update_bits_pc = dpath_io_imem_btb_update_bits_pc;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = ctrl_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = ctrl_io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_btb_update_bits_prediction_valid = ctrl_io_imem_btb_update_bits_prediction_valid;
  assign io_imem_btb_update_valid = ctrl_io_imem_btb_update_valid;
  assign io_imem_resp_ready = ctrl_io_imem_resp_ready;
  assign io_imem_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign io_imem_req_valid = ctrl_io_imem_req_valid;
  assign io_host_debug_stats_pcr = dpath_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = dpath_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = dpath_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = dpath_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = dpath_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = dpath_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = dpath_io_host_pcr_req_ready;
  Control ctrl(.clk(clk), .reset(reset),
       .io_dpath_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_dpath_killd( ctrl_io_dpath_killd ),
       .io_dpath_ren_1( ctrl_io_dpath_ren_1 ),
       .io_dpath_ren_0( ctrl_io_dpath_ren_0 ),
       .io_dpath_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_dpath_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_dpath_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_dpath_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_dpath_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_dpath_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_dpath_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_dpath_div_val(  )
       //.io_dpath_div_kill(  )
       .io_dpath_csr( ctrl_io_dpath_csr ),
       .io_dpath_sret( ctrl_io_dpath_sret ),
       .io_dpath_mem_load( ctrl_io_dpath_mem_load ),
       .io_dpath_wb_load( ctrl_io_dpath_wb_load ),
       .io_dpath_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_dpath_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_dpath_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_dpath_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_dpath_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_dpath_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_dpath_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_dpath_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_dpath_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_dpath_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_dpath_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_dpath_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_dpath_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_dpath_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_dpath_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_dpath_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_dpath_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_dpath_retire( ctrl_io_dpath_retire ),
       .io_dpath_exception( ctrl_io_dpath_exception ),
       .io_dpath_cause( ctrl_io_dpath_cause ),
       .io_dpath_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_dpath_inst( dpath_io_ctrl_inst ),
       //.io_dpath_jalr_eq(  )
       .io_dpath_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_dpath_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_dpath_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_dpath_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_dpath_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_dpath_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_dpath_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_dpath_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_dpath_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_dpath_status_ip( dpath_io_ctrl_status_ip ),
       .io_dpath_status_im( dpath_io_ctrl_status_im ),
       .io_dpath_status_zero( dpath_io_ctrl_status_zero ),
       .io_dpath_status_er( dpath_io_ctrl_status_er ),
       .io_dpath_status_vm( dpath_io_ctrl_status_vm ),
       .io_dpath_status_s64( dpath_io_ctrl_status_s64 ),
       .io_dpath_status_u64( dpath_io_ctrl_status_u64 ),
       .io_dpath_status_ef( dpath_io_ctrl_status_ef ),
       .io_dpath_status_pei( dpath_io_ctrl_status_pei ),
       .io_dpath_status_ei( dpath_io_ctrl_status_ei ),
       .io_dpath_status_ps( dpath_io_ctrl_status_ps ),
       .io_dpath_status_s( dpath_io_ctrl_status_s ),
       .io_dpath_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_dpath_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_dpath_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_imem_req_valid( ctrl_io_imem_req_valid ),
       //.io_imem_req_bits_pc(  )
       .io_imem_resp_ready( ctrl_io_imem_resp_ready ),
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( io_imem_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( ctrl_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( ctrl_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( ctrl_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( ctrl_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( ctrl_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( ctrl_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( ctrl_io_imem_btb_update_bits_prediction_bits_bht_value ),
       //.io_imem_btb_update_bits_pc(  )
       //.io_imem_btb_update_bits_target(  )
       //.io_imem_btb_update_bits_returnAddr(  )
       .io_imem_btb_update_bits_taken( ctrl_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( ctrl_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( ctrl_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( ctrl_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_mispredict( ctrl_io_imem_btb_update_bits_mispredict ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( ctrl_io_imem_invalidate ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       .io_dmem_req_valid( ctrl_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( ctrl_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( ctrl_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( ctrl_io_dmem_req_bits_phys ),
       //.io_dmem_req_bits_addr(  )
       //.io_dmem_req_bits_data(  )
       //.io_dmem_req_bits_tag(  )
       .io_dmem_req_bits_cmd( ctrl_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_fpu_valid( ctrl_io_fpu_valid ),
       .io_fpu_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_fpu_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_fpu_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_fpu_killx( ctrl_io_fpu_killx ),
       .io_fpu_killm( ctrl_io_fpu_killm ),
       .io_fpu_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_fpu_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_fpu_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_fpu_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_fpu_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_fpu_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_fpu_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_fpu_dec_single( FPU_io_ctrl_dec_single ),
       .io_fpu_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_fpu_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_fpu_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_fpu_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_fpu_dec_round( FPU_io_ctrl_dec_round ),
       .io_fpu_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_fpu_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_fpu_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( ctrl_io_rocc_cmd_valid ),
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( ctrl_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( ctrl_io_rocc_exception )
  );
  Datapath dpath(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( dpath_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( dpath_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( dpath_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( dpath_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( dpath_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( dpath_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( dpath_io_host_debug_stats_pcr ),
       .io_ctrl_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_ctrl_killd( ctrl_io_dpath_killd ),
       .io_ctrl_ren_1( ctrl_io_dpath_ren_1 ),
       .io_ctrl_ren_0( ctrl_io_dpath_ren_0 ),
       .io_ctrl_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_ctrl_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_ctrl_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_ctrl_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_ctrl_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_ctrl_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_ctrl_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_ctrl_div_val(  )
       //.io_ctrl_div_kill(  )
       .io_ctrl_csr( ctrl_io_dpath_csr ),
       .io_ctrl_sret( ctrl_io_dpath_sret ),
       .io_ctrl_mem_load( ctrl_io_dpath_mem_load ),
       .io_ctrl_wb_load( ctrl_io_dpath_wb_load ),
       .io_ctrl_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_ctrl_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_ctrl_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_ctrl_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_ctrl_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_ctrl_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_ctrl_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_ctrl_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_ctrl_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_ctrl_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_ctrl_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_ctrl_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_ctrl_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_ctrl_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_ctrl_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_ctrl_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_ctrl_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_ctrl_retire( ctrl_io_dpath_retire ),
       .io_ctrl_exception( ctrl_io_dpath_exception ),
       .io_ctrl_cause( ctrl_io_dpath_cause ),
       .io_ctrl_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_ctrl_inst( dpath_io_ctrl_inst ),
       //.io_ctrl_jalr_eq(  )
       .io_ctrl_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_ctrl_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_ctrl_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_ctrl_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_ctrl_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_ctrl_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_ctrl_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_ctrl_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_ctrl_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_ctrl_status_ip( dpath_io_ctrl_status_ip ),
       .io_ctrl_status_im( dpath_io_ctrl_status_im ),
       .io_ctrl_status_zero( dpath_io_ctrl_status_zero ),
       .io_ctrl_status_er( dpath_io_ctrl_status_er ),
       .io_ctrl_status_vm( dpath_io_ctrl_status_vm ),
       .io_ctrl_status_s64( dpath_io_ctrl_status_s64 ),
       .io_ctrl_status_u64( dpath_io_ctrl_status_u64 ),
       .io_ctrl_status_ef( dpath_io_ctrl_status_ef ),
       .io_ctrl_status_pei( dpath_io_ctrl_status_pei ),
       .io_ctrl_status_ei( dpath_io_ctrl_status_ei ),
       .io_ctrl_status_ps( dpath_io_ctrl_status_ps ),
       .io_ctrl_status_s( dpath_io_ctrl_status_s ),
       .io_ctrl_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_ctrl_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_ctrl_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       //.io_dmem_req_valid(  )
       //.io_dmem_req_bits_kill(  )
       //.io_dmem_req_bits_typ(  )
       //.io_dmem_req_bits_phys(  )
       .io_dmem_req_bits_addr( dpath_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( dpath_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( dpath_io_dmem_req_bits_tag ),
       //.io_dmem_req_bits_cmd(  )
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_ptw_ptbr( dpath_io_ptw_ptbr ),
       .io_ptw_invalidate( dpath_io_ptw_invalidate ),
       .io_ptw_sret( dpath_io_ptw_sret ),
       .io_ptw_status_ip( dpath_io_ptw_status_ip ),
       .io_ptw_status_im( dpath_io_ptw_status_im ),
       .io_ptw_status_zero( dpath_io_ptw_status_zero ),
       .io_ptw_status_er( dpath_io_ptw_status_er ),
       .io_ptw_status_vm( dpath_io_ptw_status_vm ),
       .io_ptw_status_s64( dpath_io_ptw_status_s64 ),
       .io_ptw_status_u64( dpath_io_ptw_status_u64 ),
       .io_ptw_status_ef( dpath_io_ptw_status_ef ),
       .io_ptw_status_pei( dpath_io_ptw_status_pei ),
       .io_ptw_status_ei( dpath_io_ptw_status_ei ),
       .io_ptw_status_ps( dpath_io_ptw_status_ps ),
       .io_ptw_status_s( dpath_io_ptw_status_s ),
       //.io_imem_req_valid(  )
       .io_imem_req_bits_pc( dpath_io_imem_req_bits_pc ),
       //.io_imem_resp_ready(  )
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( io_imem_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       //.io_imem_btb_update_valid(  )
       //.io_imem_btb_update_bits_prediction_valid(  )
       //.io_imem_btb_update_bits_prediction_bits_taken(  )
       //.io_imem_btb_update_bits_prediction_bits_target(  )
       //.io_imem_btb_update_bits_prediction_bits_entry(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_history(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_value(  )
       .io_imem_btb_update_bits_pc( dpath_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( dpath_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( dpath_io_imem_btb_update_bits_returnAddr ),
       //.io_imem_btb_update_bits_taken(  )
       //.io_imem_btb_update_bits_isJump(  )
       //.io_imem_btb_update_bits_isCall(  )
       //.io_imem_btb_update_bits_isReturn(  )
       //.io_imem_btb_update_bits_mispredict(  )
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       //.io_imem_invalidate(  )
       .io_fpu_inst( dpath_io_fpu_inst ),
       .io_fpu_fromint_data( dpath_io_fpu_fromint_data ),
       .io_fpu_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_fpu_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_fpu_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_fpu_store_data( FPU_io_dpath_store_data ),
       .io_fpu_toint_data( FPU_io_dpath_toint_data ),
       .io_fpu_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_fpu_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_fpu_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_fpu_dmem_resp_data( dpath_io_fpu_dmem_resp_data ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       .io_rocc_cmd_bits_inst_funct( dpath_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( dpath_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( dpath_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( dpath_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( dpath_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( dpath_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( dpath_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( dpath_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( dpath_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( dpath_io_rocc_cmd_bits_rs2 ),
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( dpath_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( dpath_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( dpath_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( dpath_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( dpath_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( dpath_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( dpath_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( dpath_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( dpath_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( dpath_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( dpath_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( dpath_io_temac_s_axi_rready )
  );
  FPU FPU(.clk(clk), .reset(reset),
       .io_ctrl_valid( ctrl_io_fpu_valid ),
       .io_ctrl_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_ctrl_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_ctrl_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_ctrl_killx( ctrl_io_fpu_killx ),
       .io_ctrl_killm( ctrl_io_fpu_killm ),
       .io_ctrl_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_ctrl_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_ctrl_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_ctrl_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_ctrl_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_ctrl_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_ctrl_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_ctrl_dec_single( FPU_io_ctrl_dec_single ),
       .io_ctrl_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_ctrl_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_ctrl_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_ctrl_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_ctrl_dec_round( FPU_io_ctrl_dec_round ),
       .io_ctrl_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_ctrl_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_ctrl_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_dpath_inst( dpath_io_fpu_inst ),
       .io_dpath_fromint_data( dpath_io_fpu_fromint_data ),
       .io_dpath_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_dpath_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_dpath_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_dpath_store_data( FPU_io_dpath_store_data ),
       .io_dpath_toint_data( FPU_io_dpath_toint_data ),
       .io_dpath_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_dpath_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_dpath_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_dpath_dmem_resp_data( dpath_io_fpu_dmem_resp_data )
  );
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input  io_requestor_1_req_bits_kill,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_phys,
    input [43:0] io_requestor_1_req_bits_addr,
    input [63:0] io_requestor_1_req_bits_data,
    input [7:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output[2:0] io_requestor_1_resp_bits_typ,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[7:0] io_requestor_1_resp_bits_tag,
    output[3:0] io_requestor_1_resp_bits_cmd,
    output[43:0] io_requestor_1_resp_bits_addr,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[7:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    //input  io_requestor_1_ptw_req_ready
    //output io_requestor_1_ptw_req_valid
    //output[29:0] io_requestor_1_ptw_req_bits
    //input  io_requestor_1_ptw_resp_valid
    //input  io_requestor_1_ptw_resp_bits_error
    //input [18:0] io_requestor_1_ptw_resp_bits_ppn
    //input [5:0] io_requestor_1_ptw_resp_bits_perm
    //input [7:0] io_requestor_1_ptw_status_ip
    //input [7:0] io_requestor_1_ptw_status_im
    //input [6:0] io_requestor_1_ptw_status_zero
    //input  io_requestor_1_ptw_status_er
    //input  io_requestor_1_ptw_status_vm
    //input  io_requestor_1_ptw_status_s64
    //input  io_requestor_1_ptw_status_u64
    //input  io_requestor_1_ptw_status_ef
    //input  io_requestor_1_ptw_status_pei
    //input  io_requestor_1_ptw_status_ei
    //input  io_requestor_1_ptw_status_ps
    //input  io_requestor_1_ptw_status_s
    //input  io_requestor_1_ptw_invalidate
    //input  io_requestor_1_ptw_sret
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input  io_requestor_0_req_bits_kill,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_phys,
    input [43:0] io_requestor_0_req_bits_addr,
    input [63:0] io_requestor_0_req_bits_data,
    input [7:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output[2:0] io_requestor_0_resp_bits_typ,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[7:0] io_requestor_0_resp_bits_tag,
    output[3:0] io_requestor_0_resp_bits_cmd,
    output[43:0] io_requestor_0_resp_bits_addr,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[7:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_ptw_req_ready
    //output io_requestor_0_ptw_req_valid
    //output[29:0] io_requestor_0_ptw_req_bits
    //input  io_requestor_0_ptw_resp_valid
    //input  io_requestor_0_ptw_resp_bits_error
    //input [18:0] io_requestor_0_ptw_resp_bits_ppn
    //input [5:0] io_requestor_0_ptw_resp_bits_perm
    //input [7:0] io_requestor_0_ptw_status_ip
    //input [7:0] io_requestor_0_ptw_status_im
    //input [6:0] io_requestor_0_ptw_status_zero
    //input  io_requestor_0_ptw_status_er
    //input  io_requestor_0_ptw_status_vm
    //input  io_requestor_0_ptw_status_s64
    //input  io_requestor_0_ptw_status_u64
    //input  io_requestor_0_ptw_status_ef
    //input  io_requestor_0_ptw_status_pei
    //input  io_requestor_0_ptw_status_ei
    //input  io_requestor_0_ptw_status_ps
    //input  io_requestor_0_ptw_status_s
    //input  io_requestor_0_ptw_invalidate
    //input  io_requestor_0_ptw_sret
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    output[63:0] io_mem_req_bits_data,
    output[7:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered
);

  wire[4:0] T0;
  wire[7:0] T32;
  wire[8:0] T1;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[63:0] T4;
  reg  r_valid_0;
  wire[43:0] T5;
  wire T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire[7:0] T33;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[7:0] T34;
  wire[6:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[7:0] T35;
  wire[6:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[7:0] T36;
  wire[6:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
`endif

  assign io_mem_req_bits_cmd = T0;
  assign T0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T32;
  assign T32 = T1[3'h7:1'h0];
  assign T1 = io_requestor_0_req_valid ? T3 : T2;
  assign T2 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T3 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_data = T4;
  assign T4 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_addr = T5;
  assign T5 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_bits_phys = T6;
  assign T6 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_typ = T7;
  assign T7 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_kill = T8;
  assign T8 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_valid = T9;
  assign T9 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T33;
  assign T33 = {1'h0, T10};
  assign T10 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T11;
  assign T11 = io_mem_replay_next_valid & T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T34;
  assign T34 = {1'h0, T14};
  assign T14 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_replay = T15;
  assign T15 = io_mem_resp_bits_replay & T16;
  assign T16 = T17 == 1'h0;
  assign T17 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T18;
  assign T18 = io_mem_resp_bits_nack & T16;
  assign io_requestor_0_resp_valid = T19;
  assign T19 = io_mem_resp_valid & T16;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T35;
  assign T35 = {1'h0, T20};
  assign T20 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T21;
  assign T21 = io_mem_replay_next_valid & T22;
  assign T22 = T23 == 1'h1;
  assign T23 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T36;
  assign T36 = {1'h0, T24};
  assign T24 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_replay = T25;
  assign T25 = io_mem_resp_bits_replay & T26;
  assign T26 = T27 == 1'h1;
  assign T27 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T28;
  assign T28 = io_mem_resp_bits_nack & T26;
  assign io_requestor_1_resp_valid = T29;
  assign T29 = io_mem_resp_valid & T26;
  assign io_requestor_1_req_ready = T30;
  assign T30 = io_requestor_0_req_ready & T31;
  assign T31 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T36;
  wire T6;
  wire T7;
  wire[3:0] T8;
  wire T9;
  wire[2:0] T10;
  wire[5:0] T11;
  wire[2:0] T12;
  wire[511:0] T13;
  wire[1:0] T14;
  wire[25:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T36 = reset ? 1'h0 : T6;
  assign T6 = T7 ? T0 : R5;
  assign T7 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_atomic_opcode = T8;
  assign T8 = T9 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T9 = T0;
  assign io_out_bits_payload_subword_addr = T10;
  assign T10 = T9 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign io_out_bits_payload_write_mask = T11;
  assign T11 = T9 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign io_out_bits_payload_a_type = T12;
  assign T12 = T9 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign io_out_bits_payload_data = T13;
  assign T13 = T9 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign io_out_bits_payload_client_xact_id = T14;
  assign T14 = T9 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr = T15;
  assign T15 = T9 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign io_out_bits_header_dst = T16;
  assign T16 = T9 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T17;
  assign T17 = T9 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T18;
  assign T18 = T9 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T27 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T25 | T23;
  assign T23 = io_in_1_valid & T24;
  assign T24 = R5 < 1'h1;
  assign T25 = io_in_0_valid & T26;
  assign T26 = R5 < 1'h0;
  assign T27 = R5 < 1'h0;
  assign io_in_1_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T33 | T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T32 | io_in_0_valid;
  assign T32 = T25 | T23;
  assign T33 = T35 & T34;
  assign T34 = R5 < 1'h1;
  assign T35 = T25 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T7) begin
      R5 <= T0;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T30;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T30 = reset ? 1'h0 : T6;
  assign T6 = T7 ? T0 : R5;
  assign T7 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_master_xact_id = T8;
  assign T8 = T9 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T9 = T0;
  assign io_out_bits_header_dst = T10;
  assign T10 = T9 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T11;
  assign T11 = T9 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T12;
  assign T12 = T9 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T13;
  assign T13 = T14 & io_out_ready;
  assign T14 = T21 | T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = T19 | T17;
  assign T17 = io_in_1_valid & T18;
  assign T18 = R5 < 1'h1;
  assign T19 = io_in_0_valid & T20;
  assign T20 = R5 < 1'h0;
  assign T21 = R5 < 1'h0;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T27 | T24;
  assign T24 = T25 ^ 1'h1;
  assign T25 = T26 | io_in_0_valid;
  assign T26 = T19 | T17;
  assign T27 = T29 & T28;
  assign T28 = R5 < 1'h1;
  assign T29 = T19 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T7) begin
      R5 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatAppendsArbiterId(input clk, input reset,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [1:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[1:0] io_in_1_grant_bits_payload_client_xact_id,
    output[2:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [2:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [1:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[1:0] io_in_0_grant_bits_payload_client_xact_id,
    output[2:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [2:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [2:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[2:0] io_out_finish_bits_payload_master_xact_id
);

  wire[1:0] T14;
  wire[2:0] T15;
  wire[1:0] T16;
  wire[2:0] T17;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[1:0] T12;
  wire T8;
  wire T9;
  wire[1:0] T13;
  wire T10;
  wire T11;
  wire RRArbiter_0_io_in_1_ready;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_0_io_out_valid;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire[2:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[5:0] RRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_0_io_out_bits_payload_subword_addr;
  wire[3:0] RRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire RRArbiter_1_io_in_1_ready;
  wire RRArbiter_1_io_in_0_ready;
  wire RRArbiter_1_io_out_valid;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[2:0] RRArbiter_1_io_out_bits_payload_master_xact_id;


  assign T14 = T15[1'h1:1'h0];
  assign T15 = {io_in_0_acquire_bits_payload_client_xact_id, 1'h0};
  assign T16 = T17[1'h1:1'h0];
  assign T17 = {io_in_1_acquire_bits_payload_client_xact_id, 1'h1};
  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T5 ? io_in_1_grant_ready : T1;
  assign T1 = T2 ? io_in_0_grant_ready : 1'h0;
  assign T2 = T3 == 1'h0;
  assign T3 = T4;
  assign T4 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign T5 = T6 == 1'h1;
  assign T6 = T7;
  assign T7 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = T12;
  assign T12 = {1'h0, T8};
  assign T8 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T9;
  assign T9 = T2 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = T13;
  assign T13 = {1'h0, T10};
  assign T10 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T11;
  assign T11 = T5 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  RRArbiter_1 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T16 ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T14 ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_2 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketTile(input clk, input reset,
    input  io_tilelink_acquire_ready,
    output io_tilelink_acquire_valid,
    output[1:0] io_tilelink_acquire_bits_header_src,
    output[1:0] io_tilelink_acquire_bits_header_dst,
    output[25:0] io_tilelink_acquire_bits_payload_addr,
    output[1:0] io_tilelink_acquire_bits_payload_client_xact_id,
    output[511:0] io_tilelink_acquire_bits_payload_data,
    output[2:0] io_tilelink_acquire_bits_payload_a_type,
    output[5:0] io_tilelink_acquire_bits_payload_write_mask,
    output[2:0] io_tilelink_acquire_bits_payload_subword_addr,
    output[3:0] io_tilelink_acquire_bits_payload_atomic_opcode,
    output io_tilelink_grant_ready,
    input  io_tilelink_grant_valid,
    input [1:0] io_tilelink_grant_bits_header_src,
    input [1:0] io_tilelink_grant_bits_header_dst,
    input [511:0] io_tilelink_grant_bits_payload_data,
    input [1:0] io_tilelink_grant_bits_payload_client_xact_id,
    input [2:0] io_tilelink_grant_bits_payload_master_xact_id,
    input [3:0] io_tilelink_grant_bits_payload_g_type,
    input  io_tilelink_finish_ready,
    output io_tilelink_finish_valid,
    output[1:0] io_tilelink_finish_bits_header_src,
    output[1:0] io_tilelink_finish_bits_header_dst,
    output[2:0] io_tilelink_finish_bits_payload_master_xact_id,
    output io_tilelink_probe_ready,
    input  io_tilelink_probe_valid,
    input [1:0] io_tilelink_probe_bits_header_src,
    input [1:0] io_tilelink_probe_bits_header_dst,
    input [25:0] io_tilelink_probe_bits_payload_addr,
    input [2:0] io_tilelink_probe_bits_payload_master_xact_id,
    input [1:0] io_tilelink_probe_bits_payload_p_type,
    input  io_tilelink_release_ready,
    output io_tilelink_release_valid,
    output[1:0] io_tilelink_release_bits_header_src,
    output[1:0] io_tilelink_release_bits_header_dst,
    output[25:0] io_tilelink_release_bits_payload_addr,
    output[1:0] io_tilelink_release_bits_payload_client_xact_id,
    output[2:0] io_tilelink_release_bits_payload_master_xact_id,
    output[511:0] io_tilelink_release_bits_payload_data,
    output[2:0] io_tilelink_release_bits_payload_r_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready
);

  wire[1:0] T1;
  wire[2:0] T0;
  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_subword;
  wire[7:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[7:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_subword;
  wire[7:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[7:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire dcArb_io_mem_req_bits_kill;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_phys;
  wire[43:0] dcArb_io_mem_req_bits_addr;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire[7:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[18:0] ptw_io_requestor_1_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_1_resp_bits_perm;
  wire[7:0] ptw_io_requestor_1_status_ip;
  wire[7:0] ptw_io_requestor_1_status_im;
  wire[6:0] ptw_io_requestor_1_status_zero;
  wire ptw_io_requestor_1_status_er;
  wire ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_s64;
  wire ptw_io_requestor_1_status_u64;
  wire ptw_io_requestor_1_status_ef;
  wire ptw_io_requestor_1_status_pei;
  wire ptw_io_requestor_1_status_ei;
  wire ptw_io_requestor_1_status_ps;
  wire ptw_io_requestor_1_status_s;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_1_sret;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[18:0] ptw_io_requestor_0_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_0_resp_bits_perm;
  wire[7:0] ptw_io_requestor_0_status_ip;
  wire[7:0] ptw_io_requestor_0_status_im;
  wire[6:0] ptw_io_requestor_0_status_zero;
  wire ptw_io_requestor_0_status_er;
  wire ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_s64;
  wire ptw_io_requestor_0_status_u64;
  wire ptw_io_requestor_0_status_ef;
  wire ptw_io_requestor_0_status_pei;
  wire ptw_io_requestor_0_status_ei;
  wire ptw_io_requestor_0_status_ps;
  wire ptw_io_requestor_0_status_s;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_requestor_0_sret;
  wire ptw_io_mem_req_valid;
  wire ptw_io_mem_req_bits_kill;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_phys;
  wire[43:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire memArb_io_in_1_acquire_ready;
  wire memArb_io_in_1_grant_valid;
  wire[1:0] memArb_io_in_1_grant_bits_header_src;
  wire[1:0] memArb_io_in_1_grant_bits_header_dst;
  wire[511:0] memArb_io_in_1_grant_bits_payload_data;
  wire[1:0] memArb_io_in_1_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_1_grant_bits_payload_master_xact_id;
  wire[3:0] memArb_io_in_1_grant_bits_payload_g_type;
  wire memArb_io_in_1_finish_ready;
  wire memArb_io_in_0_acquire_ready;
  wire memArb_io_in_0_grant_valid;
  wire[1:0] memArb_io_in_0_grant_bits_header_src;
  wire[1:0] memArb_io_in_0_grant_bits_header_dst;
  wire[511:0] memArb_io_in_0_grant_bits_payload_data;
  wire[1:0] memArb_io_in_0_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_0_grant_bits_payload_master_xact_id;
  wire[3:0] memArb_io_in_0_grant_bits_payload_g_type;
  wire memArb_io_in_0_finish_ready;
  wire memArb_io_out_acquire_valid;
  wire[1:0] memArb_io_out_acquire_bits_header_src;
  wire[1:0] memArb_io_out_acquire_bits_header_dst;
  wire[25:0] memArb_io_out_acquire_bits_payload_addr;
  wire[1:0] memArb_io_out_acquire_bits_payload_client_xact_id;
  wire[511:0] memArb_io_out_acquire_bits_payload_data;
  wire[2:0] memArb_io_out_acquire_bits_payload_a_type;
  wire[5:0] memArb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] memArb_io_out_acquire_bits_payload_subword_addr;
  wire[3:0] memArb_io_out_acquire_bits_payload_atomic_opcode;
  wire memArb_io_out_grant_ready;
  wire memArb_io_out_finish_valid;
  wire[1:0] memArb_io_out_finish_bits_header_src;
  wire[1:0] memArb_io_out_finish_bits_header_dst;
  wire[2:0] memArb_io_out_finish_bits_payload_master_xact_id;
  wire icache_io_cpu_resp_valid;
  wire[43:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data;
  wire icache_io_cpu_resp_bits_xcpt_ma;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire[42:0] icache_io_cpu_btb_resp_bits_target;
  wire[5:0] icache_io_cpu_btb_resp_bits_entry;
  wire[6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire icache_io_cpu_ptw_req_valid;
  wire[29:0] icache_io_cpu_ptw_req_bits;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[7:0] dcache_io_cpu_resp_bits_tag;
  wire[3:0] dcache_io_cpu_resp_bits_cmd;
  wire[43:0] dcache_io_cpu_resp_bits_addr;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[7:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ptw_req_valid;
  wire[29:0] dcache_io_cpu_ptw_req_bits;
  wire dcache_io_cpu_ordered;
  wire dcache_io_mem_acquire_valid;
  wire[1:0] dcache_io_mem_acquire_bits_header_src;
  wire[1:0] dcache_io_mem_acquire_bits_header_dst;
  wire[25:0] dcache_io_mem_acquire_bits_payload_addr;
  wire[1:0] dcache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] dcache_io_mem_acquire_bits_payload_data;
  wire[2:0] dcache_io_mem_acquire_bits_payload_a_type;
  wire[5:0] dcache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] dcache_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] dcache_io_mem_acquire_bits_payload_atomic_opcode;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_finish_valid;
  wire[1:0] dcache_io_mem_finish_bits_header_src;
  wire[1:0] dcache_io_mem_finish_bits_header_dst;
  wire[2:0] dcache_io_mem_finish_bits_payload_master_xact_id;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_header_src;
  wire[1:0] dcache_io_mem_release_bits_header_dst;
  wire[25:0] dcache_io_mem_release_bits_payload_addr;
  wire[1:0] dcache_io_mem_release_bits_payload_client_xact_id;
  wire[2:0] dcache_io_mem_release_bits_payload_master_xact_id;
  wire[511:0] dcache_io_mem_release_bits_payload_data;
  wire[2:0] dcache_io_mem_release_bits_payload_r_type;
  wire core_io_host_pcr_req_ready;
  wire core_io_host_pcr_rep_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_pcr;
  wire core_io_imem_req_valid;
  wire[43:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire[42:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[42:0] core_io_imem_btb_update_bits_pc;
  wire[42:0] core_io_imem_btb_update_bits_target;
  wire[42:0] core_io_imem_btb_update_bits_returnAddr;
  wire core_io_imem_btb_update_bits_taken;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isCall;
  wire core_io_imem_btb_update_bits_isReturn;
  wire core_io_imem_btb_update_bits_mispredict;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire core_io_dmem_req_bits_kill;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_phys;
  wire[43:0] core_io_dmem_req_bits_addr;
  wire[63:0] core_io_dmem_req_bits_data;
  wire[7:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_sret;
  wire[7:0] core_io_ptw_status_ip;
  wire[7:0] core_io_ptw_status_im;
  wire[6:0] core_io_ptw_status_zero;
  wire core_io_ptw_status_er;
  wire core_io_ptw_status_vm;
  wire core_io_ptw_status_s64;
  wire core_io_ptw_status_u64;
  wire core_io_ptw_status_ef;
  wire core_io_ptw_status_pei;
  wire core_io_ptw_status_ei;
  wire core_io_ptw_status_ps;
  wire core_io_ptw_status_s;
  wire core_io_temac_rx_axis_fifo_tready;
  wire[7:0] core_io_temac_tx_axis_fifo_tdata;
  wire core_io_temac_tx_axis_fifo_tvalid;
  wire core_io_temac_tx_axis_fifo_tlast;
  wire[11:0] core_io_temac_s_axi_awaddr;
  wire core_io_temac_s_axi_awvalid;
  wire[31:0] core_io_temac_s_axi_wdata;
  wire core_io_temac_s_axi_wvalid;
  wire core_io_temac_s_axi_bready;
  wire[11:0] core_io_temac_s_axi_araddr;
  wire core_io_temac_s_axi_arvalid;
  wire core_io_temac_s_axi_rready;


  assign io_temac_s_axi_rready = core_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = core_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = core_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = core_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = core_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = core_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = core_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = core_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = core_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = core_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = core_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = core_io_temac_rx_axis_fifo_tready;
  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_tilelink_release_bits_payload_r_type = dcache_io_mem_release_bits_payload_r_type;
  assign io_tilelink_release_bits_payload_data = dcache_io_mem_release_bits_payload_data;
  assign io_tilelink_release_bits_payload_master_xact_id = dcache_io_mem_release_bits_payload_master_xact_id;
  assign io_tilelink_release_bits_payload_client_xact_id = T1;
  assign T1 = T0[1'h1:1'h0];
  assign T0 = {dcache_io_mem_release_bits_payload_client_xact_id, 1'h0};
  assign io_tilelink_release_bits_payload_addr = dcache_io_mem_release_bits_payload_addr;
  assign io_tilelink_release_bits_header_dst = dcache_io_mem_release_bits_header_dst;
  assign io_tilelink_release_bits_header_src = dcache_io_mem_release_bits_header_src;
  assign io_tilelink_release_valid = dcache_io_mem_release_valid;
  assign io_tilelink_probe_ready = dcache_io_mem_probe_ready;
  assign io_tilelink_finish_bits_payload_master_xact_id = memArb_io_out_finish_bits_payload_master_xact_id;
  assign io_tilelink_finish_bits_header_dst = memArb_io_out_finish_bits_header_dst;
  assign io_tilelink_finish_bits_header_src = memArb_io_out_finish_bits_header_src;
  assign io_tilelink_finish_valid = memArb_io_out_finish_valid;
  assign io_tilelink_grant_ready = memArb_io_out_grant_ready;
  assign io_tilelink_acquire_bits_payload_atomic_opcode = memArb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_tilelink_acquire_bits_payload_subword_addr = memArb_io_out_acquire_bits_payload_subword_addr;
  assign io_tilelink_acquire_bits_payload_write_mask = memArb_io_out_acquire_bits_payload_write_mask;
  assign io_tilelink_acquire_bits_payload_a_type = memArb_io_out_acquire_bits_payload_a_type;
  assign io_tilelink_acquire_bits_payload_data = memArb_io_out_acquire_bits_payload_data;
  assign io_tilelink_acquire_bits_payload_client_xact_id = memArb_io_out_acquire_bits_payload_client_xact_id;
  assign io_tilelink_acquire_bits_payload_addr = memArb_io_out_acquire_bits_payload_addr;
  assign io_tilelink_acquire_bits_header_dst = memArb_io_out_acquire_bits_header_dst;
  assign io_tilelink_acquire_bits_header_src = memArb_io_out_acquire_bits_header_src;
  assign io_tilelink_acquire_valid = memArb_io_out_acquire_valid;
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_cpu_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_cpu_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_mispredict( core_io_imem_btb_update_bits_mispredict ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_cpu_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_0_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_0_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_0_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_0_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_0_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_0_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_0_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_0_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_0_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_0_sret ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_mem_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_1_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_1_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_cpu_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_1_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_1_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_1_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_1_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_1_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_1_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_1_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_1_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_1_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_1_sret ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_mem_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_mem_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_mem_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_0_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_0_finish_ready ),
       .io_mem_finish_valid( dcache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_tilelink_probe_valid ),
       .io_mem_probe_bits_header_src( io_tilelink_probe_bits_header_src ),
       .io_mem_probe_bits_header_dst( io_tilelink_probe_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( io_tilelink_probe_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( io_tilelink_probe_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( io_tilelink_probe_bits_payload_p_type ),
       .io_mem_release_ready( io_tilelink_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_mem_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_mem_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( dcache_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_requestor_1_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_requestor_1_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_requestor_1_status_ip( ptw_io_requestor_1_status_ip ),
       .io_requestor_1_status_im( ptw_io_requestor_1_status_im ),
       .io_requestor_1_status_zero( ptw_io_requestor_1_status_zero ),
       .io_requestor_1_status_er( ptw_io_requestor_1_status_er ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_requestor_1_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_requestor_1_status_ef( ptw_io_requestor_1_status_ef ),
       .io_requestor_1_status_pei( ptw_io_requestor_1_status_pei ),
       .io_requestor_1_status_ei( ptw_io_requestor_1_status_ei ),
       .io_requestor_1_status_ps( ptw_io_requestor_1_status_ps ),
       .io_requestor_1_status_s( ptw_io_requestor_1_status_s ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_1_sret( ptw_io_requestor_1_sret ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_requestor_0_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_requestor_0_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_requestor_0_status_ip( ptw_io_requestor_0_status_ip ),
       .io_requestor_0_status_im( ptw_io_requestor_0_status_im ),
       .io_requestor_0_status_zero( ptw_io_requestor_0_status_zero ),
       .io_requestor_0_status_er( ptw_io_requestor_0_status_er ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_requestor_0_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_requestor_0_status_ef( ptw_io_requestor_0_status_ef ),
       .io_requestor_0_status_pei( ptw_io_requestor_0_status_pei ),
       .io_requestor_0_status_ei( ptw_io_requestor_0_status_ei ),
       .io_requestor_0_status_ps( ptw_io_requestor_0_status_ps ),
       .io_requestor_0_status_s( ptw_io_requestor_0_status_s ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_requestor_0_sret( ptw_io_requestor_0_sret ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_data(  )
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       //.io_mem_ptw_req_valid(  )
       //.io_mem_ptw_req_bits(  )
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_sret( core_io_ptw_sret ),
       .io_dpath_status_ip( core_io_ptw_status_ip ),
       .io_dpath_status_im( core_io_ptw_status_im ),
       .io_dpath_status_zero( core_io_ptw_status_zero ),
       .io_dpath_status_er( core_io_ptw_status_er ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_s64( core_io_ptw_status_s64 ),
       .io_dpath_status_u64( core_io_ptw_status_u64 ),
       .io_dpath_status_ef( core_io_ptw_status_ef ),
       .io_dpath_status_pei( core_io_ptw_status_pei ),
       .io_dpath_status_ei( core_io_ptw_status_ei ),
       .io_dpath_status_ps( core_io_ptw_status_ps ),
       .io_dpath_status_s( core_io_ptw_status_s )
  );
  Core core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_imem_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_mispredict( core_io_imem_btb_update_bits_mispredict ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_imem_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       //.io_dmem_ptw_req_valid(  )
       //.io_dmem_ptw_req_bits(  )
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_sret( core_io_ptw_sret ),
       .io_ptw_status_ip( core_io_ptw_status_ip ),
       .io_ptw_status_im( core_io_ptw_status_im ),
       .io_ptw_status_zero( core_io_ptw_status_zero ),
       .io_ptw_status_er( core_io_ptw_status_er ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_s64( core_io_ptw_status_s64 ),
       .io_ptw_status_u64( core_io_ptw_status_u64 ),
       .io_ptw_status_ef( core_io_ptw_status_ef ),
       .io_ptw_status_pei( core_io_ptw_status_pei ),
       .io_ptw_status_ei( core_io_ptw_status_ei ),
       .io_ptw_status_ps( core_io_ptw_status_ps ),
       .io_ptw_status_s( core_io_ptw_status_s ),
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_write_mask(  )
       //.io_rocc_imem_acquire_bits_payload_subword_addr(  )
       //.io_rocc_imem_acquire_bits_payload_atomic_opcode(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       //.io_rocc_imem_finish_valid(  )
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( core_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( core_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( core_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( core_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( core_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( core_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( core_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( core_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( core_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( core_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( core_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( core_io_temac_s_axi_rready )
  );
  `ifndef SYNTHESIS
    assign core.io_dmem_ptw_req_valid = {1{$random}};
    assign core.io_dmem_ptw_req_bits = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_ptw_req_ready = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_valid = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_error = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_ppn = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_perm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ip = {1{$random}};
    assign core.io_rocc_mem_ptw_status_im = {1{$random}};
    assign core.io_rocc_mem_ptw_status_zero = {1{$random}};
    assign core.io_rocc_mem_ptw_status_er = {1{$random}};
    assign core.io_rocc_mem_ptw_status_vm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_u64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ef = {1{$random}};
    assign core.io_rocc_mem_ptw_status_pei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ps = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s = {1{$random}};
    assign core.io_rocc_mem_ptw_invalidate = {1{$random}};
    assign core.io_rocc_mem_ptw_sret = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_data = {16{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_write_mask = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_subword_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_atomic_opcode = {1{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_imem_finish_valid = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_finish_bits_payload_master_xact_id = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits = {1{$random}};
  `endif
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_requestor_1_ptw_req_ready(  )
       //.io_requestor_1_ptw_req_valid(  )
       //.io_requestor_1_ptw_req_bits(  )
       //.io_requestor_1_ptw_resp_valid(  )
       //.io_requestor_1_ptw_resp_bits_error(  )
       //.io_requestor_1_ptw_resp_bits_ppn(  )
       //.io_requestor_1_ptw_resp_bits_perm(  )
       //.io_requestor_1_ptw_status_ip(  )
       //.io_requestor_1_ptw_status_im(  )
       //.io_requestor_1_ptw_status_zero(  )
       //.io_requestor_1_ptw_status_er(  )
       //.io_requestor_1_ptw_status_vm(  )
       //.io_requestor_1_ptw_status_s64(  )
       //.io_requestor_1_ptw_status_u64(  )
       //.io_requestor_1_ptw_status_ef(  )
       //.io_requestor_1_ptw_status_pei(  )
       //.io_requestor_1_ptw_status_ei(  )
       //.io_requestor_1_ptw_status_ps(  )
       //.io_requestor_1_ptw_status_s(  )
       //.io_requestor_1_ptw_invalidate(  )
       //.io_requestor_1_ptw_sret(  )
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_data(  )
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_ptw_req_ready(  )
       //.io_requestor_0_ptw_req_valid(  )
       //.io_requestor_0_ptw_req_bits(  )
       //.io_requestor_0_ptw_resp_valid(  )
       //.io_requestor_0_ptw_resp_bits_error(  )
       //.io_requestor_0_ptw_resp_bits_ppn(  )
       //.io_requestor_0_ptw_resp_bits_perm(  )
       //.io_requestor_0_ptw_status_ip(  )
       //.io_requestor_0_ptw_status_im(  )
       //.io_requestor_0_ptw_status_zero(  )
       //.io_requestor_0_ptw_status_er(  )
       //.io_requestor_0_ptw_status_vm(  )
       //.io_requestor_0_ptw_status_s64(  )
       //.io_requestor_0_ptw_status_u64(  )
       //.io_requestor_0_ptw_status_ef(  )
       //.io_requestor_0_ptw_status_pei(  )
       //.io_requestor_0_ptw_status_ei(  )
       //.io_requestor_0_ptw_status_ps(  )
       //.io_requestor_0_ptw_status_s(  )
       //.io_requestor_0_ptw_invalidate(  )
       //.io_requestor_0_ptw_sret(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_mem_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
  `ifndef SYNTHESIS
    assign dcArb.io_requestor_0_req_bits_data = {2{$random}};
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
  `endif
  UncachedTileLinkIOArbiterThatAppendsArbiterId memArb(.clk(clk), .reset(reset),
       .io_in_1_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_in_1_acquire_bits_header_src(  )
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( icache_io_mem_grant_ready ),
       .io_in_1_grant_valid( memArb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( memArb_io_in_1_finish_ready ),
       .io_in_1_finish_valid( icache_io_mem_finish_valid ),
       .io_in_1_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_in_1_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_in_1_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_in_0_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_in_0_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( dcache_io_mem_grant_ready ),
       .io_in_0_grant_valid( memArb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( memArb_io_in_0_finish_ready ),
       .io_in_0_finish_valid( dcache_io_mem_finish_valid ),
       .io_in_0_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_in_0_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_in_0_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_acquire_ready( io_tilelink_acquire_ready ),
       .io_out_acquire_valid( memArb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( memArb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( memArb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( memArb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( memArb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( memArb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( memArb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( memArb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( memArb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( memArb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( memArb_io_out_grant_ready ),
       .io_out_grant_valid( io_tilelink_grant_valid ),
       .io_out_grant_bits_header_src( io_tilelink_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_tilelink_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_tilelink_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_tilelink_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_tilelink_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_tilelink_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_tilelink_finish_ready ),
       .io_out_finish_valid( memArb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( memArb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( memArb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( memArb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign memArb.io_in_1_acquire_bits_header_src = {1{$random}};
    assign memArb.io_in_1_acquire_bits_header_dst = {1{$random}};
  `endif
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [1:0] io_enq_bits_client_xact_id,
    input [511:0] io_enq_bits_data,
    input [2:0] io_enq_bits_a_type,
    input [5:0] io_enq_bits_write_mask,
    input [2:0] io_enq_bits_subword_addr,
    input [3:0] io_enq_bits_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[1:0] io_deq_bits_client_xact_id,
    output[511:0] io_deq_bits_data,
    output[2:0] io_deq_bits_a_type,
    output[5:0] io_deq_bits_write_mask,
    output[2:0] io_deq_bits_subword_addr,
    output[3:0] io_deq_bits_atomic_opcode,
    output io_count
);

  wire T21;
  wire[1:0] T0;
  reg  full;
  wire T22;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[3:0] T3;
  wire[555:0] T4;
  reg [555:0] ram [0:0];
  wire[555:0] T5;
  wire[555:0] T6;
  wire[555:0] T7;
  wire[15:0] T8;
  wire[6:0] T9;
  wire[8:0] T10;
  wire[539:0] T11;
  wire[513:0] T12;
  wire[2:0] T13;
  wire[5:0] T14;
  wire[2:0] T15;
  wire[511:0] T16;
  wire[1:0] T17;
  wire[25:0] T18;
  wire T19;
  wire empty;
  wire T20;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {18{$random}};
  end
`endif

  assign io_count = T21;
  assign T21 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T22 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_atomic_opcode = T3;
  assign T3 = T4[2'h3:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_subword_addr, io_enq_bits_atomic_opcode};
  assign T10 = {io_enq_bits_a_type, io_enq_bits_write_mask};
  assign T11 = {io_enq_bits_addr, T12};
  assign T12 = {io_enq_bits_client_xact_id, io_enq_bits_data};
  assign io_deq_bits_subword_addr = T13;
  assign T13 = T4[3'h6:3'h4];
  assign io_deq_bits_write_mask = T14;
  assign T14 = T4[4'hc:3'h7];
  assign io_deq_bits_a_type = T15;
  assign T15 = T4[4'hf:4'hd];
  assign io_deq_bits_data = T16;
  assign T16 = T4[10'h20f:5'h10];
  assign io_deq_bits_client_xact_id = T17;
  assign T17 = T4[10'h211:10'h210];
  assign io_deq_bits_addr = T18;
  assign T18 = T4[10'h22b:10'h212];
  assign io_deq_valid = T19;
  assign T19 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[4:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    //output[1:0] io_mem_finish_bits_header_src
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [2:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    //output[1:0] io_mem_release_bits_header_src
    //output[1:0] io_mem_release_bits_header_dst
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[2:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire T350;
  reg [3:0] cmd;
  wire[3:0] T20;
  wire[3:0] next_cmd;
  wire[63:0] rx_shifter_in;
  wire[47:0] T30;
  reg [63:0] rx_shifter;
  wire[63:0] T31;
  wire T59;
  wire T21;
  wire T22;
  reg [14:0] rx_count;
  wire[14:0] T337;
  wire[14:0] T23;
  wire[14:0] T24;
  wire[14:0] T25;
  wire T26;
  wire T27;
  wire[12:0] T338;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T28;
  wire[11:0] T29;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire nack;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire bad_mem_packet;
  wire T44;
  wire[2:0] T45;
  reg [39:0] addr;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire T96;
  wire T97;
  reg [3:0] state;
  wire[3:0] T336;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  wire[3:0] rx_cmd;
  wire T60;
  wire[12:0] rx_word_count;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire rx_done;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire T69;
  wire[12:0] T340;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire rx_word_done;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  reg  mem_acked;
  wire T341;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire[3:0] T88;
  wire T89;
  wire T90;
  reg [8:0] pos;
  wire[8:0] T91;
  wire[8:0] T92;
  wire[8:0] T93;
  wire[8:0] T94;
  wire T95;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T112;
  wire T113;
  wire T114;
  wire[4:0] pcr_addr;
  wire T115;
  wire T116;
  wire[1:0] pcr_coreid;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T339;
  wire[14:0] T55;
  wire[14:0] T56;
  wire[14:0] T57;
  wire T58;
  wire T102;
  wire tx_done;
  wire T103;
  wire T104;
  wire T105;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T106;
  wire T107;
  wire T108;
  wire[12:0] T342;
  wire T109;
  wire T110;
  wire[1:0] tx_subword_count;
  wire T111;
  wire[2:0] T351;
  wire[2:0] T352;
  wire[2:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[2:0] T357;
  wire[2:0] T358;
  wire[2:0] T359;
  wire[511:0] T360;
  wire[511:0] T361;
  wire[511:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[25:0] T366;
  wire[25:0] T367;
  wire[25:0] T368;
  wire[36:0] init_addr;
  wire[39:0] T369;
  wire[25:0] T370;
  wire[25:0] T371;
  wire T372;
  wire T373;
  wire T374;
  wire[63:0] pcr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  wire[63:0] T121;
  wire[63:0] T122;
  wire T123;
  wire T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire T128;
  wire[63:0] T129;
  wire[63:0] T130;
  wire T131;
  wire T132;
  wire[63:0] T133;
  wire[63:0] T134;
  wire T135;
  wire T136;
  wire[63:0] T137;
  wire[63:0] T138;
  wire T139;
  wire T140;
  wire[63:0] T141;
  wire[63:0] T142;
  wire T143;
  wire T144;
  wire[63:0] T145;
  wire[63:0] T146;
  wire T147;
  wire T148;
  wire[63:0] T149;
  wire T150;
  wire[2:0] T151;
  wire[2:0] T152;
  wire[5:0] T153;
  wire[5:0] scr_addr;
  wire T154;
  wire T155;
  reg [2:0] mem_gxid;
  wire[2:0] T156;
  reg [1:0] mem_gsrc;
  wire[1:0] T157;
  wire T158;
  reg  mem_needs_ack;
  wire T159;
  wire T160;
  wire T161;
  wire[511:0] mem_req_data;
  wire[447:0] T162;
  wire[383:0] T163;
  wire[319:0] T164;
  wire[255:0] T165;
  wire[191:0] T166;
  wire[127:0] T167;
  wire[63:0] T168;
  wire[63:0] T169;
  wire[63:0] T170;
  wire[63:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[63:0] T174;
  wire[63:0] T175;
  reg  R176;
  wire T343;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  reg  R186;
  wire T344;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[15:0] T345;
  wire[63:0] T191;
  wire[5:0] T192;
  wire[1:0] T193;
  wire[63:0] tx_data;
  wire[63:0] T194;
  wire[63:0] T195;
  reg [63:0] pcrReadData;
  wire[63:0] T196;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T346;
  wire[63:0] T199;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  wire[63:0] T203;
  wire[63:0] T204;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T205;
  wire[5:0] T206;
  wire[63:0] T207;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T208;
  wire T209;
  wire[63:0] T210;
  wire[63:0] T211;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T212;
  wire[63:0] T213;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T214;
  wire T215;
  wire T216;
  wire[63:0] T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T220;
  wire[63:0] T221;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T222;
  wire T223;
  wire[63:0] T224;
  wire[63:0] T225;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T226;
  wire[63:0] T227;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[63:0] T232;
  wire[63:0] T233;
  wire[63:0] T234;
  wire[63:0] T235;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T236;
  wire[63:0] T237;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T238;
  wire T239;
  wire[63:0] T240;
  wire[63:0] T241;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T242;
  wire[63:0] T243;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T244;
  wire T245;
  wire T246;
  wire[63:0] T247;
  wire[63:0] T248;
  wire[63:0] T249;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T250;
  wire[63:0] T251;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T252;
  wire T253;
  wire[63:0] T254;
  wire[63:0] T255;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T256;
  wire[63:0] T257;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire[63:0] T263;
  wire[63:0] T264;
  wire[63:0] T265;
  wire[63:0] T266;
  wire[63:0] T267;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T268;
  wire[63:0] T269;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T270;
  wire T271;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T274;
  wire[63:0] T275;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T276;
  wire T277;
  wire T278;
  wire[63:0] T279;
  wire[63:0] T280;
  wire[63:0] T281;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T282;
  wire[63:0] T283;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T284;
  wire T285;
  wire[63:0] T286;
  wire[63:0] T287;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T288;
  wire[63:0] T289;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[63:0] T294;
  wire[63:0] T295;
  wire[63:0] T296;
  wire[63:0] T297;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T298;
  wire[63:0] T299;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T300;
  wire T301;
  wire[63:0] T302;
  wire[63:0] T303;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T304;
  wire[63:0] T305;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T306;
  wire T307;
  wire T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T312;
  wire[63:0] T313;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T314;
  wire T315;
  wire[63:0] T316;
  wire[63:0] T317;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T318;
  wire[63:0] T319;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[63:0] tx_header;
  wire[15:0] T329;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T330;
  reg [7:0] seqno;
  wire[7:0] T331;
  wire[7:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire acq_q_io_enq_ready;
  wire acq_q_io_deq_valid;
  wire[25:0] acq_q_io_deq_bits_addr;
  wire[1:0] acq_q_io_deq_bits_client_xact_id;
  wire[2:0] acq_q_io_deq_bits_a_type;
  wire[5:0] acq_q_io_deq_bits_write_mask;
  wire[2:0] acq_q_io_deq_bits_subword_addr;
  wire[3:0] acq_q_io_deq_bits_atomic_opcode;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cmd = {1{$random}};
    rx_shifter = {2{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    addr = {2{$random}};
    state = {1{$random}};
    mem_acked = {1{$random}};
    pos = {1{$random}};
    tx_count = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    mem_gxid = {1{$random}};
    mem_gsrc = {1{$random}};
    mem_needs_ack = {1{$random}};
    R176 = {1{$random}};
    R186 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
`endif

  assign T347 = T350 ? T349 : T348;
  assign T348 = 4'h0;
  assign T349 = 4'h0;
  assign T350 = cmd == 4'h1;
  assign T20 = T21 ? next_cmd : cmd;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign rx_shifter_in = {io_host_in_bits, T30};
  assign T30 = rx_shifter[6'h3f:5'h10];
  assign T31 = T59 ? rx_shifter_in : rx_shifter;
  assign T59 = io_host_in_valid & io_host_in_ready;
  assign T21 = T59 & T22;
  assign T22 = rx_count == 15'h3;
  assign T337 = reset ? 15'h0 : T23;
  assign T23 = T26 ? 15'h0 : T24;
  assign T24 = T59 ? T25 : rx_count;
  assign T25 = rx_count + 15'h1;
  assign T26 = T102 & T27;
  assign T27 = tx_word_count == T338;
  assign T338 = {1'h0, tx_size};
  assign tx_size = T32 ? size : 12'h0;
  assign T28 = T21 ? T29 : size;
  assign T29 = rx_shifter_in[4'hf:3'h4];
  assign T32 = T38 & T33;
  assign T33 = T35 | T34;
  assign T34 = cmd == 4'h3;
  assign T35 = T37 | T36;
  assign T36 = cmd == 4'h2;
  assign T37 = cmd == 4'h0;
  assign T38 = nack ^ 1'h1;
  assign nack = T52 ? bad_mem_packet : T39;
  assign T39 = T41 ? T40 : 1'h1;
  assign T40 = size != 12'h1;
  assign T41 = T43 | T42;
  assign T42 = cmd == 4'h3;
  assign T43 = cmd == 4'h2;
  assign bad_mem_packet = T50 | T44;
  assign T44 = T45 != 3'h0;
  assign T45 = addr[2'h2:1'h0];
  assign T46 = T96 ? T49 : T47;
  assign T47 = T21 ? T48 : addr;
  assign T48 = rx_shifter_in[6'h3f:5'h18];
  assign T49 = addr + 40'h8;
  assign T96 = T97 & io_mem_finish_ready;
  assign T97 = state == 4'h7;
  assign T336 = reset ? 4'h0 : T4;
  assign T4 = T118 ? 4'h8 : T5;
  assign T5 = io_cpu_0_pcr_rep_valid ? 4'h8 : T6;
  assign T6 = T113 ? 4'h8 : T7;
  assign T7 = T112 ? 4'h2 : T8;
  assign T8 = T102 ? T98 : T9;
  assign T9 = T96 ? T88 : T10;
  assign T10 = T87 ? 4'h7 : T11;
  assign T11 = T81 ? 4'h7 : T12;
  assign T12 = T79 ? 4'h5 : T13;
  assign T13 = T77 ? 4'h6 : T14;
  assign T14 = T64 ? T15 : state;
  assign T15 = T63 ? 4'h3 : T16;
  assign T16 = T62 ? 4'h4 : T17;
  assign T17 = T18 ? 4'h1 : 4'h8;
  assign T18 = T61 | T19;
  assign T19 = rx_cmd == 4'h3;
  assign rx_cmd = T60 ? next_cmd : cmd;
  assign T60 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T61 = rx_cmd == 4'h2;
  assign T62 = rx_cmd == 4'h1;
  assign T63 = rx_cmd == 4'h0;
  assign T64 = T76 & rx_done;
  assign rx_done = rx_word_done & T65;
  assign T65 = T73 ? T70 : T66;
  assign T66 = T69 | T67;
  assign T67 = T68 == 3'h0;
  assign T68 = rx_word_count[2'h2:1'h0];
  assign T69 = rx_word_count == T340;
  assign T340 = {1'h0, size};
  assign T70 = T72 & T71;
  assign T71 = next_cmd != 4'h3;
  assign T72 = next_cmd != 4'h1;
  assign T73 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T74;
  assign T74 = T75 == 2'h3;
  assign T75 = rx_count[1'h1:1'h0];
  assign T76 = state == 4'h0;
  assign T77 = T78 & acq_q_io_enq_ready;
  assign T78 = state == 4'h4;
  assign T79 = T80 & acq_q_io_enq_ready;
  assign T80 = state == 4'h3;
  assign T81 = T86 & mem_acked;
  assign T341 = reset ? 1'h0 : T82;
  assign T82 = T85 ? 1'h0 : T83;
  assign T83 = T81 ? 1'h0 : T84;
  assign T84 = io_mem_grant_valid ? 1'h1 : mem_acked;
  assign T85 = state == 4'h5;
  assign T86 = state == 4'h6;
  assign T87 = T85 & io_mem_grant_valid;
  assign T88 = T89 ? 4'h8 : 4'h0;
  assign T89 = T95 | T90;
  assign T90 = pos == 9'h1;
  assign T91 = T96 ? T94 : T92;
  assign T92 = T21 ? T93 : pos;
  assign T93 = rx_shifter_in[4'hf:3'h7];
  assign T94 = pos - 9'h1;
  assign T95 = cmd == 4'h0;
  assign T98 = T99 ? 4'h3 : 4'h0;
  assign T99 = T101 & T100;
  assign T100 = pos != 9'h0;
  assign T101 = cmd == 4'h0;
  assign T112 = io_cpu_0_pcr_req_valid & io_cpu_0_pcr_req_ready;
  assign T113 = T115 & T114;
  assign T114 = pcr_addr == 5'h1d;
  assign pcr_addr = addr[3'h4:1'h0];
  assign T115 = T117 & T116;
  assign T116 = pcr_coreid == 2'h0;
  assign pcr_coreid = addr[5'h15:5'h14];
  assign T117 = state == 4'h1;
  assign T118 = T120 & T119;
  assign T119 = pcr_coreid == 2'h3;
  assign T120 = state == 4'h1;
  assign T50 = T51 != 3'h0;
  assign T51 = size[2'h2:1'h0];
  assign T52 = T54 | T53;
  assign T53 = cmd == 4'h1;
  assign T54 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T339 = reset ? 15'h0 : T55;
  assign T55 = T26 ? 15'h0 : T56;
  assign T56 = T58 ? T57 : tx_count;
  assign T57 = tx_count + 15'h1;
  assign T58 = io_host_out_valid & io_host_out_ready;
  assign T102 = T111 & tx_done;
  assign tx_done = T109 & T103;
  assign T103 = T108 | T104;
  assign T104 = T107 & T105;
  assign T105 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T106 - 3'h1;
  assign T106 = tx_word_count[2'h2:1'h0];
  assign T107 = 13'h0 < tx_word_count;
  assign T108 = tx_word_count == T342;
  assign T342 = {1'h0, tx_size};
  assign T109 = io_host_out_ready & T110;
  assign T110 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T111 = state == 4'h8;
  assign T351 = T350 ? T353 : T352;
  assign T352 = 3'h0;
  assign T353 = 3'h0;
  assign T354 = T350 ? T356 : T355;
  assign T355 = 6'h0;
  assign T356 = 6'h0;
  assign T357 = T350 ? T359 : T358;
  assign T358 = 3'h2;
  assign T359 = 3'h3;
  assign T360 = T350 ? T362 : T361;
  assign T361 = 512'h0;
  assign T362 = 512'h0;
  assign T363 = T350 ? T365 : T364;
  assign T364 = 2'h0;
  assign T365 = 2'h0;
  assign T366 = T350 ? T370 : T367;
  assign T367 = T368;
  assign T368 = init_addr[5'h19:1'h0];
  assign init_addr = T369 >> 2'h3;
  assign T369 = addr;
  assign T370 = T371;
  assign T371 = init_addr[5'h19:1'h0];
  assign T372 = T374 | T373;
  assign T373 = state == 4'h4;
  assign T374 = state == 4'h3;
  assign io_scr_wdata = pcr_wdata;
  assign pcr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_payload_data[9'h1ff:9'h1c0];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 4'h5;
  assign T122 = io_mem_grant_bits_payload_data[9'h1bf:9'h180];
  assign T123 = T124 & io_mem_grant_valid;
  assign T124 = state == 4'h5;
  assign T126 = io_mem_grant_bits_payload_data[9'h17f:9'h140];
  assign T127 = T128 & io_mem_grant_valid;
  assign T128 = state == 4'h5;
  assign T130 = io_mem_grant_bits_payload_data[9'h13f:9'h100];
  assign T131 = T132 & io_mem_grant_valid;
  assign T132 = state == 4'h5;
  assign T134 = io_mem_grant_bits_payload_data[8'hff:8'hc0];
  assign T135 = T136 & io_mem_grant_valid;
  assign T136 = state == 4'h5;
  assign T138 = io_mem_grant_bits_payload_data[8'hbf:8'h80];
  assign T139 = T140 & io_mem_grant_valid;
  assign T140 = state == 4'h5;
  assign T142 = io_mem_grant_bits_payload_data[7'h7f:7'h40];
  assign T143 = T144 & io_mem_grant_valid;
  assign T144 = state == 4'h5;
  assign T146 = io_mem_grant_bits_payload_data[6'h3f:1'h0];
  assign T147 = T148 & io_mem_grant_valid;
  assign T148 = state == 4'h5;
  assign T150 = rx_word_done & io_host_in_ready;
  assign T151 = T152 - 3'h1;
  assign T152 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T153;
  assign T153 = scr_addr;
  assign scr_addr = addr[3'h5:1'h0];
  assign io_scr_wen = T154;
  assign T154 = T118 ? T155 : 1'h0;
  assign T155 = cmd == 4'h3;
  assign io_mem_release_valid = 1'h0;
  assign io_mem_probe_ready = 1'h0;
  assign io_mem_finish_bits_payload_master_xact_id = mem_gxid;
  assign T156 = io_mem_grant_valid ? io_mem_grant_bits_payload_master_xact_id : mem_gxid;
  assign io_mem_finish_bits_header_dst = mem_gsrc;
  assign T157 = io_mem_grant_valid ? io_mem_grant_bits_header_src : mem_gsrc;
  assign io_mem_finish_valid = T158;
  assign T158 = T161 & mem_needs_ack;
  assign T159 = io_mem_grant_valid ? T160 : mem_needs_ack;
  assign T160 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T161 = state == 4'h7;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_payload_atomic_opcode = acq_q_io_deq_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = acq_q_io_deq_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = acq_q_io_deq_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = acq_q_io_deq_bits_a_type;
  assign io_mem_acquire_bits_payload_data = mem_req_data;
  assign mem_req_data = {T175, T162};
  assign T162 = {T174, T163};
  assign T163 = {T173, T164};
  assign T164 = {T172, T165};
  assign T165 = {T171, T166};
  assign T166 = {T170, T167};
  assign T167 = {T169, T168};
  assign T168 = packet_ram[3'h0];
  assign T169 = packet_ram[3'h1];
  assign T170 = packet_ram[3'h2];
  assign T171 = packet_ram[3'h3];
  assign T172 = packet_ram[3'h4];
  assign T173 = packet_ram[3'h5];
  assign T174 = packet_ram[3'h6];
  assign T175 = packet_ram[3'h7];
  assign io_mem_acquire_bits_payload_client_xact_id = acq_q_io_deq_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = acq_q_io_deq_bits_addr;
  assign io_mem_acquire_bits_header_dst = 2'h0;
  assign io_mem_acquire_bits_header_src = 2'h2;
  assign io_mem_acquire_valid = acq_q_io_deq_valid;
  assign io_cpu_0_ipi_rep_valid = R176;
  assign T343 = reset ? 1'h0 : T177;
  assign T177 = T179 ? 1'h1 : T178;
  assign T178 = io_cpu_0_ipi_rep_ready ? 1'h0 : R176;
  assign T179 = io_cpu_0_ipi_req_valid & T180;
  assign T180 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = pcr_wdata;
  assign io_cpu_0_pcr_req_bits_addr = pcr_addr;
  assign io_cpu_0_pcr_req_bits_rw = T181;
  assign T181 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T182;
  assign T182 = T184 & T183;
  assign T183 = pcr_addr != 5'h1d;
  assign T184 = T185 & T116;
  assign T185 = state == 4'h1;
  assign io_cpu_0_reset = R186;
  assign T344 = reset ? 1'h1 : T187;
  assign T187 = T189 ? T188 : R186;
  assign T188 = pcr_wdata[1'h0:1'h0];
  assign T189 = T113 & T190;
  assign T190 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T345;
  assign T345 = T191[4'hf:1'h0];
  assign T191 = tx_data >> T192;
  assign T192 = {T193, 4'h0};
  assign T193 = tx_count[1'h1:1'h0];
  assign tx_data = T333 ? tx_header : T194;
  assign T194 = T326 ? pcrReadData : T195;
  assign T195 = packet_ram[packet_ram_raddr];
  assign T196 = T118 ? T199 : T197;
  assign T197 = io_cpu_0_pcr_rep_valid ? io_cpu_0_pcr_rep_bits : T198;
  assign T198 = T113 ? T346 : pcrReadData;
  assign T346 = {63'h0, R186};
  assign T199 = T325 ? T263 : T200;
  assign T200 = T262 ? T232 : T201;
  assign T201 = T231 ? T217 : T202;
  assign T202 = T216 ? T210 : T203;
  assign T203 = T209 ? T207 : T204;
  assign T204 = T205 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T205 = T206[1'h0:1'h0];
  assign T206 = scr_addr;
  assign T207 = T208 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T208 = T206[1'h0:1'h0];
  assign T209 = T206[1'h1:1'h1];
  assign T210 = T215 ? T213 : T211;
  assign T211 = T212 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T212 = T206[1'h0:1'h0];
  assign T213 = T214 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T214 = T206[1'h0:1'h0];
  assign T215 = T206[1'h1:1'h1];
  assign T216 = T206[2'h2:2'h2];
  assign T217 = T230 ? T224 : T218;
  assign T218 = T223 ? T221 : T219;
  assign T219 = T220 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T220 = T206[1'h0:1'h0];
  assign T221 = T222 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T222 = T206[1'h0:1'h0];
  assign T223 = T206[1'h1:1'h1];
  assign T224 = T229 ? T227 : T225;
  assign T225 = T226 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T226 = T206[1'h0:1'h0];
  assign T227 = T228 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T228 = T206[1'h0:1'h0];
  assign T229 = T206[1'h1:1'h1];
  assign T230 = T206[2'h2:2'h2];
  assign T231 = T206[2'h3:2'h3];
  assign T232 = T261 ? T247 : T233;
  assign T233 = T246 ? T240 : T234;
  assign T234 = T239 ? T237 : T235;
  assign T235 = T236 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T236 = T206[1'h0:1'h0];
  assign T237 = T238 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T238 = T206[1'h0:1'h0];
  assign T239 = T206[1'h1:1'h1];
  assign T240 = T245 ? T243 : T241;
  assign T241 = T242 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T242 = T206[1'h0:1'h0];
  assign T243 = T244 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T244 = T206[1'h0:1'h0];
  assign T245 = T206[1'h1:1'h1];
  assign T246 = T206[2'h2:2'h2];
  assign T247 = T260 ? T254 : T248;
  assign T248 = T253 ? T251 : T249;
  assign T249 = T250 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T250 = T206[1'h0:1'h0];
  assign T251 = T252 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T252 = T206[1'h0:1'h0];
  assign T253 = T206[1'h1:1'h1];
  assign T254 = T259 ? T257 : T255;
  assign T255 = T256 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T256 = T206[1'h0:1'h0];
  assign T257 = T258 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T258 = T206[1'h0:1'h0];
  assign T259 = T206[1'h1:1'h1];
  assign T260 = T206[2'h2:2'h2];
  assign T261 = T206[2'h3:2'h3];
  assign T262 = T206[3'h4:3'h4];
  assign T263 = T324 ? T294 : T264;
  assign T264 = T293 ? T279 : T265;
  assign T265 = T278 ? T272 : T266;
  assign T266 = T271 ? T269 : T267;
  assign T267 = T268 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T268 = T206[1'h0:1'h0];
  assign T269 = T270 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T270 = T206[1'h0:1'h0];
  assign T271 = T206[1'h1:1'h1];
  assign T272 = T277 ? T275 : T273;
  assign T273 = T274 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T274 = T206[1'h0:1'h0];
  assign T275 = T276 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T276 = T206[1'h0:1'h0];
  assign T277 = T206[1'h1:1'h1];
  assign T278 = T206[2'h2:2'h2];
  assign T279 = T292 ? T286 : T280;
  assign T280 = T285 ? T283 : T281;
  assign T281 = T282 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T282 = T206[1'h0:1'h0];
  assign T283 = T284 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T284 = T206[1'h0:1'h0];
  assign T285 = T206[1'h1:1'h1];
  assign T286 = T291 ? T289 : T287;
  assign T287 = T288 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T288 = T206[1'h0:1'h0];
  assign T289 = T290 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T290 = T206[1'h0:1'h0];
  assign T291 = T206[1'h1:1'h1];
  assign T292 = T206[2'h2:2'h2];
  assign T293 = T206[2'h3:2'h3];
  assign T294 = T323 ? T309 : T295;
  assign T295 = T308 ? T302 : T296;
  assign T296 = T301 ? T299 : T297;
  assign T297 = T298 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T298 = T206[1'h0:1'h0];
  assign T299 = T300 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T300 = T206[1'h0:1'h0];
  assign T301 = T206[1'h1:1'h1];
  assign T302 = T307 ? T305 : T303;
  assign T303 = T304 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T304 = T206[1'h0:1'h0];
  assign T305 = T306 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T306 = T206[1'h0:1'h0];
  assign T307 = T206[1'h1:1'h1];
  assign T308 = T206[2'h2:2'h2];
  assign T309 = T322 ? T316 : T310;
  assign T310 = T315 ? T313 : T311;
  assign T311 = T312 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T312 = T206[1'h0:1'h0];
  assign T313 = T314 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T314 = T206[1'h0:1'h0];
  assign T315 = T206[1'h1:1'h1];
  assign T316 = T321 ? T319 : T317;
  assign T317 = T318 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T318 = T206[1'h0:1'h0];
  assign T319 = T320 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T320 = T206[1'h0:1'h0];
  assign T321 = T206[1'h1:1'h1];
  assign T322 = T206[2'h2:2'h2];
  assign T323 = T206[2'h3:2'h3];
  assign T324 = T206[3'h4:3'h4];
  assign T325 = T206[3'h5:3'h5];
  assign T326 = T328 | T327;
  assign T327 = cmd == 4'h3;
  assign T328 = cmd == 4'h2;
  assign tx_header = {T330, T329};
  assign T329 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T330 = {addr, seqno};
  assign T331 = T21 ? T332 : seqno;
  assign T332 = rx_shifter_in[5'h17:5'h10];
  assign T333 = tx_word_count == 13'h0;
  assign io_host_out_valid = T334;
  assign T334 = state == 4'h8;
  assign io_host_in_ready = T335;
  assign T335 = state == 4'h0;
  Queue_8 acq_q(.clk(clk), .reset(reset),
       .io_enq_ready( acq_q_io_enq_ready ),
       .io_enq_valid( T372 ),
       .io_enq_bits_addr( T366 ),
       .io_enq_bits_client_xact_id( T363 ),
       .io_enq_bits_data( T360 ),
       .io_enq_bits_a_type( T357 ),
       .io_enq_bits_write_mask( T354 ),
       .io_enq_bits_subword_addr( T351 ),
       .io_enq_bits_atomic_opcode( T347 ),
       .io_deq_ready( io_mem_acquire_ready ),
       .io_deq_valid( acq_q_io_deq_valid ),
       .io_deq_bits_addr( acq_q_io_deq_bits_addr ),
       .io_deq_bits_client_xact_id( acq_q_io_deq_bits_client_xact_id ),
       //.io_deq_bits_data(  )
       .io_deq_bits_a_type( acq_q_io_deq_bits_a_type ),
       .io_deq_bits_write_mask( acq_q_io_deq_bits_write_mask ),
       .io_deq_bits_subword_addr( acq_q_io_deq_bits_subword_addr ),
       .io_deq_bits_atomic_opcode( acq_q_io_deq_bits_atomic_opcode )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T21) begin
      cmd <= next_cmd;
    end
    if(T59) begin
      rx_shifter <= rx_shifter_in;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T26) begin
      rx_count <= 15'h0;
    end else if(T59) begin
      rx_count <= T25;
    end
    if(T21) begin
      size <= T29;
    end
    if(T96) begin
      addr <= T49;
    end else if(T21) begin
      addr <= T48;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T118) begin
      state <= 4'h8;
    end else if(io_cpu_0_pcr_rep_valid) begin
      state <= 4'h8;
    end else if(T113) begin
      state <= 4'h8;
    end else if(T112) begin
      state <= 4'h2;
    end else if(T102) begin
      state <= T98;
    end else if(T96) begin
      state <= T88;
    end else if(T87) begin
      state <= 4'h7;
    end else if(T81) begin
      state <= 4'h7;
    end else if(T79) begin
      state <= 4'h5;
    end else if(T77) begin
      state <= 4'h6;
    end else if(T64) begin
      state <= T15;
    end
    if(reset) begin
      mem_acked <= 1'h0;
    end else if(T85) begin
      mem_acked <= 1'h0;
    end else if(T81) begin
      mem_acked <= 1'h0;
    end else if(io_mem_grant_valid) begin
      mem_acked <= 1'h1;
    end
    if(T96) begin
      pos <= T94;
    end else if(T21) begin
      pos <= T93;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T26) begin
      tx_count <= 15'h0;
    end else if(T58) begin
      tx_count <= T57;
    end
    if (T2)
      packet_ram[3'h7] <= T1;
    if (T123)
      packet_ram[3'h6] <= T122;
    if (T127)
      packet_ram[3'h5] <= T126;
    if (T131)
      packet_ram[3'h4] <= T130;
    if (T135)
      packet_ram[3'h3] <= T134;
    if (T139)
      packet_ram[3'h2] <= T138;
    if (T143)
      packet_ram[3'h1] <= T142;
    if (T147)
      packet_ram[3'h0] <= T146;
    if (T150)
      packet_ram[T151] <= rx_shifter_in;
    if(io_mem_grant_valid) begin
      mem_gxid <= io_mem_grant_bits_payload_master_xact_id;
    end
    if(io_mem_grant_valid) begin
      mem_gsrc <= io_mem_grant_bits_header_src;
    end
    if(io_mem_grant_valid) begin
      mem_needs_ack <= T160;
    end
    if(reset) begin
      R176 <= 1'h0;
    end else if(T179) begin
      R176 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R176 <= 1'h0;
    end
    if(reset) begin
      R186 <= 1'h1;
    end else if(T189) begin
      R186 <= T188;
    end
    if(T118) begin
      pcrReadData <= T199;
    end else if(io_cpu_0_pcr_rep_valid) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T113) begin
      pcrReadData <= T346;
    end
    if(T21) begin
      seqno <= T332;
    end
  end
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T83;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[5:0] T19;
  wire[5:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire T25;
  wire T26;
  wire[511:0] T27;
  wire[511:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[25:0] T35;
  wire[25:0] T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T83 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_atomic_opcode = T10;
  assign T10 = T14 ? io_in_2_bits_payload_atomic_opcode : T11;
  assign T11 = T12 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_subword_addr = T15;
  assign T15 = T18 ? io_in_2_bits_payload_subword_addr : T16;
  assign T16 = T17 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_write_mask = T19;
  assign T19 = T22 ? io_in_2_bits_payload_write_mask : T20;
  assign T20 = T21 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T23;
  assign T23 = T26 ? io_in_2_bits_payload_a_type : T24;
  assign T24 = T25 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T27;
  assign T27 = T30 ? io_in_2_bits_payload_data : T28;
  assign T28 = T29 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T31;
  assign T31 = T34 ? io_in_2_bits_payload_client_xact_id : T32;
  assign T32 = T33 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T35;
  assign T35 = T38 ? io_in_2_bits_payload_addr : T36;
  assign T36 = T37 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T39;
  assign T39 = T42 ? io_in_2_bits_header_dst : T40;
  assign T40 = T41 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T41 = T13[1'h0:1'h0];
  assign T42 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T43;
  assign T43 = T46 ? io_in_2_bits_header_src : T44;
  assign T44 = T45 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T45 = T13[1'h0:1'h0];
  assign T46 = T13[1'h1:1'h1];
  assign io_out_valid = T47;
  assign T47 = T50 ? io_in_2_valid : T48;
  assign T48 = T49 ? io_in_1_valid : io_in_0_valid;
  assign T49 = T13[1'h0:1'h0];
  assign T50 = T13[1'h1:1'h1];
  assign io_in_0_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T62 | T53;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T57 | T55;
  assign T55 = io_in_2_valid & T56;
  assign T56 = last_grant < 2'h2;
  assign T57 = T60 | T58;
  assign T58 = io_in_1_valid & T59;
  assign T59 = last_grant < 2'h1;
  assign T60 = io_in_0_valid & T61;
  assign T61 = last_grant < 2'h0;
  assign T62 = last_grant < 2'h0;
  assign io_in_1_ready = T63;
  assign T63 = T64 & io_out_ready;
  assign T64 = T69 | T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_0_valid;
  assign T67 = T68 | T55;
  assign T68 = T60 | T58;
  assign T69 = T71 & T70;
  assign T70 = last_grant < 2'h1;
  assign T71 = T60 ^ 1'h1;
  assign io_in_2_ready = T72;
  assign T72 = T73 & io_out_ready;
  assign T73 = T79 | T74;
  assign T74 = T75 ^ 1'h1;
  assign T75 = T76 | io_in_1_valid;
  assign T76 = T77 | io_in_0_valid;
  assign T77 = T78 | T55;
  assign T78 = T60 | T58;
  assign T79 = T81 & T80;
  assign T80 = last_grant < 2'h2;
  assign T81 = T82 ^ 1'h1;
  assign T82 = T60 | T58;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_a_type,
    output[5:0] io_out_2_bits_payload_write_mask,
    output[2:0] io_out_2_bits_payload_subword_addr,
    output[3:0] io_out_2_bits_payload_atomic_opcode,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_a_type,
    output[5:0] io_out_1_bits_payload_write_mask,
    output[2:0] io_out_1_bits_payload_subword_addr,
    output[3:0] io_out_1_bits_payload_atomic_opcode,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_a_type,
    output[5:0] io_out_0_bits_payload_write_mask,
    output[2:0] io_out_0_bits_payload_subword_addr,
    output[3:0] io_out_0_bits_payload_atomic_opcode
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_0_io_in_2_ready;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire LockingRRArbiter_0_io_out_valid;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_a_type;
  wire[5:0] LockingRRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_a_type;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_a_type;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_atomic_opcode = LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_0_bits_payload_subword_addr = LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_0_bits_payload_write_mask = LockingRRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_atomic_opcode = LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  assign io_out_1_bits_payload_subword_addr = LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  assign io_out_1_bits_payload_write_mask = LockingRRArbiter_1_io_out_bits_payload_write_mask;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_1_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_atomic_opcode = LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;
  assign io_out_2_bits_payload_subword_addr = LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  assign io_out_2_bits_payload_write_mask = LockingRRArbiter_2_io_out_bits_payload_write_mask;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_2_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_1_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_0_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_2_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_1_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_0_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_2_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_1_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_0_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_0 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_1_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_1_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_1_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_1_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_2_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_2_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_2_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T75;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[511:0] T15;
  wire[511:0] T16;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[25:0] T27;
  wire[25:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T75 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_r_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_r_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T15;
  assign T15 = T18 ? io_in_2_bits_payload_data : T16;
  assign T16 = T17 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T19;
  assign T19 = T22 ? io_in_2_bits_payload_master_xact_id : T20;
  assign T20 = T21 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T23;
  assign T23 = T26 ? io_in_2_bits_payload_client_xact_id : T24;
  assign T24 = T25 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T27;
  assign T27 = T30 ? io_in_2_bits_payload_addr : T28;
  assign T28 = T29 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T31;
  assign T31 = T34 ? io_in_2_bits_header_dst : T32;
  assign T32 = T33 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T35;
  assign T35 = T38 ? io_in_2_bits_header_src : T36;
  assign T36 = T37 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_out_valid = T39;
  assign T39 = T42 ? io_in_2_valid : T40;
  assign T40 = T41 ? io_in_1_valid : io_in_0_valid;
  assign T41 = T13[1'h0:1'h0];
  assign T42 = T13[1'h1:1'h1];
  assign io_in_0_ready = T43;
  assign T43 = T44 & io_out_ready;
  assign T44 = T54 | T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T49 | T47;
  assign T47 = io_in_2_valid & T48;
  assign T48 = last_grant < 2'h2;
  assign T49 = T52 | T50;
  assign T50 = io_in_1_valid & T51;
  assign T51 = last_grant < 2'h1;
  assign T52 = io_in_0_valid & T53;
  assign T53 = last_grant < 2'h0;
  assign T54 = last_grant < 2'h0;
  assign io_in_1_ready = T55;
  assign T55 = T56 & io_out_ready;
  assign T56 = T61 | T57;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T59 | io_in_0_valid;
  assign T59 = T60 | T47;
  assign T60 = T52 | T50;
  assign T61 = T63 & T62;
  assign T62 = last_grant < 2'h1;
  assign T63 = T52 ^ 1'h1;
  assign io_in_2_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T71 | T66;
  assign T66 = T67 ^ 1'h1;
  assign T67 = T68 | io_in_1_valid;
  assign T68 = T69 | io_in_0_valid;
  assign T69 = T70 | T47;
  assign T70 = T52 | T50;
  assign T71 = T73 & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T52 | T50;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_r_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_r_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_r_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[1:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_3_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_master_xact_id;
  wire[511:0] LockingRRArbiter_3_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_r_type;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[1:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_4_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_master_xact_id;
  wire[511:0] LockingRRArbiter_4_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_r_type;
  wire LockingRRArbiter_5_io_in_2_ready;
  wire LockingRRArbiter_5_io_in_1_ready;
  wire LockingRRArbiter_5_io_in_0_ready;
  wire LockingRRArbiter_5_io_out_valid;
  wire[1:0] LockingRRArbiter_5_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_5_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_5_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_5_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_5_io_out_bits_payload_master_xact_id;
  wire[511:0] LockingRRArbiter_5_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_5_io_out_bits_payload_r_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_3_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_3_io_out_bits_payload_data;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_3_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_3_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_4_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_4_io_out_bits_payload_data;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_4_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_4_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_4_io_out_valid;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_5_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_5_io_out_bits_payload_data;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_5_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_5_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_5_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_5_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_5_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_5_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_5_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_4_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_3_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_5_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_4_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_3_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_5_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_4_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_3_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_1 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_3_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_3_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_3_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_3_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_3_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_4_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_4_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_4_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_4_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_4_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_5(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_5_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_5_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_5_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_5_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_5_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_5_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_5_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_5_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_5_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_5_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_5_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T67;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[25:0] T19;
  wire[25:0] T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T67 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_p_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_p_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T15;
  assign T15 = T18 ? io_in_2_bits_payload_master_xact_id : T16;
  assign T16 = T17 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T19;
  assign T19 = T22 ? io_in_2_bits_payload_addr : T20;
  assign T20 = T21 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T23;
  assign T23 = T26 ? io_in_2_bits_header_dst : T24;
  assign T24 = T25 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T27;
  assign T27 = T30 ? io_in_2_bits_header_src : T28;
  assign T28 = T29 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_valid = T31;
  assign T31 = T34 ? io_in_2_valid : T32;
  assign T32 = T33 ? io_in_1_valid : io_in_0_valid;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_in_0_ready = T35;
  assign T35 = T36 & io_out_ready;
  assign T36 = T46 | T37;
  assign T37 = T38 ^ 1'h1;
  assign T38 = T41 | T39;
  assign T39 = io_in_2_valid & T40;
  assign T40 = last_grant < 2'h2;
  assign T41 = T44 | T42;
  assign T42 = io_in_1_valid & T43;
  assign T43 = last_grant < 2'h1;
  assign T44 = io_in_0_valid & T45;
  assign T45 = last_grant < 2'h0;
  assign T46 = last_grant < 2'h0;
  assign io_in_1_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T53 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_0_valid;
  assign T51 = T52 | T39;
  assign T52 = T44 | T42;
  assign T53 = T55 & T54;
  assign T54 = last_grant < 2'h1;
  assign T55 = T44 ^ 1'h1;
  assign io_in_2_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = T63 | T58;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_1_valid;
  assign T60 = T61 | io_in_0_valid;
  assign T61 = T62 | T39;
  assign T62 = T44 | T42;
  assign T63 = T65 & T64;
  assign T64 = last_grant < 2'h2;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T44 | T42;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_6_io_in_2_ready;
  wire LockingRRArbiter_6_io_in_1_ready;
  wire LockingRRArbiter_6_io_in_0_ready;
  wire LockingRRArbiter_6_io_out_valid;
  wire[1:0] LockingRRArbiter_6_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_6_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_6_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_6_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_6_io_out_bits_payload_p_type;
  wire LockingRRArbiter_7_io_in_2_ready;
  wire LockingRRArbiter_7_io_in_1_ready;
  wire LockingRRArbiter_7_io_in_0_ready;
  wire LockingRRArbiter_7_io_out_valid;
  wire[1:0] LockingRRArbiter_7_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_7_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_7_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_7_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_7_io_out_bits_payload_p_type;
  wire LockingRRArbiter_8_io_in_2_ready;
  wire LockingRRArbiter_8_io_in_1_ready;
  wire LockingRRArbiter_8_io_in_0_ready;
  wire LockingRRArbiter_8_io_out_valid;
  wire[1:0] LockingRRArbiter_8_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_8_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_8_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_8_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_8_io_out_bits_payload_p_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_6_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_6_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_6_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_6_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_6_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_6_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_7_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_7_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_7_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_7_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_7_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_7_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_8_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_8_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_8_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_8_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_8_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_8_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_8_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_7_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_6_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_8_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_7_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_6_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_8_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_7_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_6_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_2 LockingRRArbiter_6(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_6_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_6_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_6_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_6_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_6_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_6_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_6_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_6_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_6_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_7(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_7_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_7_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_7_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_7_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_7_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_7_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_7_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_7_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_7_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_8(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_8_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_8_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_8_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_8_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_8_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_8_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_8_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_8_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_8_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T71;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[511:0] T23;
  wire[511:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T71 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_g_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_g_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T15;
  assign T15 = T18 ? io_in_2_bits_payload_master_xact_id : T16;
  assign T16 = T17 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T19;
  assign T19 = T22 ? io_in_2_bits_payload_client_xact_id : T20;
  assign T20 = T21 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T23;
  assign T23 = T26 ? io_in_2_bits_payload_data : T24;
  assign T24 = T25 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T27;
  assign T27 = T30 ? io_in_2_bits_header_dst : T28;
  assign T28 = T29 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T31;
  assign T31 = T34 ? io_in_2_bits_header_src : T32;
  assign T32 = T33 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_valid = T35;
  assign T35 = T38 ? io_in_2_valid : T36;
  assign T36 = T37 ? io_in_1_valid : io_in_0_valid;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_in_0_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T50 | T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T45 | T43;
  assign T43 = io_in_2_valid & T44;
  assign T44 = last_grant < 2'h2;
  assign T45 = T48 | T46;
  assign T46 = io_in_1_valid & T47;
  assign T47 = last_grant < 2'h1;
  assign T48 = io_in_0_valid & T49;
  assign T49 = last_grant < 2'h0;
  assign T50 = last_grant < 2'h0;
  assign io_in_1_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T57 | T53;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T55 | io_in_0_valid;
  assign T55 = T56 | T43;
  assign T56 = T48 | T46;
  assign T57 = T59 & T58;
  assign T58 = last_grant < 2'h1;
  assign T59 = T48 ^ 1'h1;
  assign io_in_2_ready = T60;
  assign T60 = T61 & io_out_ready;
  assign T61 = T67 | T62;
  assign T62 = T63 ^ 1'h1;
  assign T63 = T64 | io_in_1_valid;
  assign T64 = T65 | io_in_0_valid;
  assign T65 = T66 | T43;
  assign T66 = T48 | T46;
  assign T67 = T69 & T68;
  assign T68 = last_grant < 2'h2;
  assign T69 = T70 ^ 1'h1;
  assign T70 = T48 | T46;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[511:0] io_out_2_bits_payload_data,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[3:0] io_out_2_bits_payload_g_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[511:0] io_out_1_bits_payload_data,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[3:0] io_out_1_bits_payload_g_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[511:0] io_out_0_bits_payload_data,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[3:0] io_out_0_bits_payload_g_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_9_io_in_2_ready;
  wire LockingRRArbiter_9_io_in_1_ready;
  wire LockingRRArbiter_9_io_in_0_ready;
  wire LockingRRArbiter_9_io_out_valid;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_9_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_9_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_9_io_out_bits_payload_g_type;
  wire LockingRRArbiter_10_io_in_2_ready;
  wire LockingRRArbiter_10_io_in_1_ready;
  wire LockingRRArbiter_10_io_in_0_ready;
  wire LockingRRArbiter_10_io_out_valid;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_10_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_10_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_10_io_out_bits_payload_g_type;
  wire LockingRRArbiter_11_io_in_2_ready;
  wire LockingRRArbiter_11_io_in_1_ready;
  wire LockingRRArbiter_11_io_in_0_ready;
  wire LockingRRArbiter_11_io_out_valid;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_11_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_11_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_11_io_out_bits_payload_g_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_9_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_9_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_data = LockingRRArbiter_9_io_out_bits_payload_data;
  assign io_out_0_bits_header_dst = LockingRRArbiter_9_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_9_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_9_io_out_valid;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_10_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_10_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_data = LockingRRArbiter_10_io_out_bits_payload_data;
  assign io_out_1_bits_header_dst = LockingRRArbiter_10_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_10_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_10_io_out_valid;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_11_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_11_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_data = LockingRRArbiter_11_io_out_bits_payload_data;
  assign io_out_2_bits_header_dst = LockingRRArbiter_11_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_11_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_11_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_11_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_10_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_9_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_11_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_10_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_9_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_11_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_10_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_9_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_3 LockingRRArbiter_9(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_9_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_9_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_9_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_9_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_9_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_9_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_9_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_9_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_9_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_9_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_10(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_10_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_10_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_10_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_10_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_10_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_10_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_10_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_10_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_10_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_10_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_11(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_11_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_11_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_11_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_11_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_11_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_11_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_11_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_11_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_11_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_11_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T59;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T59 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_master_xact_id = T10;
  assign T10 = T14 ? io_in_2_bits_payload_master_xact_id : T11;
  assign T11 = T12 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T15;
  assign T15 = T18 ? io_in_2_bits_header_dst : T16;
  assign T16 = T17 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T19;
  assign T19 = T22 ? io_in_2_bits_header_src : T20;
  assign T20 = T21 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_valid = T23;
  assign T23 = T26 ? io_in_2_valid : T24;
  assign T24 = T25 ? io_in_1_valid : io_in_0_valid;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_in_0_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T38 | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T33 | T31;
  assign T31 = io_in_2_valid & T32;
  assign T32 = last_grant < 2'h2;
  assign T33 = T36 | T34;
  assign T34 = io_in_1_valid & T35;
  assign T35 = last_grant < 2'h1;
  assign T36 = io_in_0_valid & T37;
  assign T37 = last_grant < 2'h0;
  assign T38 = last_grant < 2'h0;
  assign io_in_1_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T45 | T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T43 | io_in_0_valid;
  assign T43 = T44 | T31;
  assign T44 = T36 | T34;
  assign T45 = T47 & T46;
  assign T46 = last_grant < 2'h1;
  assign T47 = T36 ^ 1'h1;
  assign io_in_2_ready = T48;
  assign T48 = T49 & io_out_ready;
  assign T49 = T55 | T50;
  assign T50 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_1_valid;
  assign T52 = T53 | io_in_0_valid;
  assign T53 = T54 | T31;
  assign T54 = T36 | T34;
  assign T55 = T57 & T56;
  assign T56 = last_grant < 2'h2;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T36 | T34;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[2:0] io_out_0_bits_payload_master_xact_id
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_12_io_in_2_ready;
  wire LockingRRArbiter_12_io_in_1_ready;
  wire LockingRRArbiter_12_io_in_0_ready;
  wire LockingRRArbiter_12_io_out_valid;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_12_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_13_io_in_2_ready;
  wire LockingRRArbiter_13_io_in_1_ready;
  wire LockingRRArbiter_13_io_in_0_ready;
  wire LockingRRArbiter_13_io_out_valid;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_13_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_14_io_in_2_ready;
  wire LockingRRArbiter_14_io_in_1_ready;
  wire LockingRRArbiter_14_io_in_0_ready;
  wire LockingRRArbiter_14_io_out_valid;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_14_io_out_bits_payload_master_xact_id;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_12_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_12_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_12_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_12_io_out_valid;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_13_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_13_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_13_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_13_io_out_valid;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_14_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_14_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_14_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_14_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_14_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_13_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_12_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_14_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_13_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_12_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_14_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_13_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_12_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_4 LockingRRArbiter_12(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_12_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_12_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_12_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_12_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_12_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_12_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_12_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_13(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_13_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_13_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_13_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_13_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_13_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_13_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_13_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_14(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_14_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_14_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_14_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_14_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_14_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_14_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_14_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketChipCrossbarNetwork(input clk, input reset,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [1:0] io_clients_1_acquire_bits_header_src,
    input [1:0] io_clients_1_acquire_bits_header_dst,
    input [25:0] io_clients_1_acquire_bits_payload_addr,
    input [1:0] io_clients_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_1_acquire_bits_payload_data,
    input [2:0] io_clients_1_acquire_bits_payload_a_type,
    input [5:0] io_clients_1_acquire_bits_payload_write_mask,
    input [2:0] io_clients_1_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_1_acquire_bits_payload_atomic_opcode,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_header_src,
    output[1:0] io_clients_1_grant_bits_header_dst,
    output[511:0] io_clients_1_grant_bits_payload_data,
    output[1:0] io_clients_1_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_1_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_1_grant_bits_payload_g_type,
    output io_clients_1_finish_ready,
    input  io_clients_1_finish_valid,
    input [1:0] io_clients_1_finish_bits_header_src,
    input [1:0] io_clients_1_finish_bits_header_dst,
    input [2:0] io_clients_1_finish_bits_payload_master_xact_id,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[1:0] io_clients_1_probe_bits_header_src,
    output[1:0] io_clients_1_probe_bits_header_dst,
    output[25:0] io_clients_1_probe_bits_payload_addr,
    output[2:0] io_clients_1_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_1_probe_bits_payload_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_header_src,
    input [1:0] io_clients_1_release_bits_header_dst,
    input [25:0] io_clients_1_release_bits_payload_addr,
    input [1:0] io_clients_1_release_bits_payload_client_xact_id,
    input [2:0] io_clients_1_release_bits_payload_master_xact_id,
    input [511:0] io_clients_1_release_bits_payload_data,
    input [2:0] io_clients_1_release_bits_payload_r_type,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [1:0] io_clients_0_acquire_bits_header_src,
    input [1:0] io_clients_0_acquire_bits_header_dst,
    input [25:0] io_clients_0_acquire_bits_payload_addr,
    input [1:0] io_clients_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_0_acquire_bits_payload_data,
    input [2:0] io_clients_0_acquire_bits_payload_a_type,
    input [5:0] io_clients_0_acquire_bits_payload_write_mask,
    input [2:0] io_clients_0_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_0_acquire_bits_payload_atomic_opcode,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_header_src,
    output[1:0] io_clients_0_grant_bits_header_dst,
    output[511:0] io_clients_0_grant_bits_payload_data,
    output[1:0] io_clients_0_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_0_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_0_grant_bits_payload_g_type,
    output io_clients_0_finish_ready,
    input  io_clients_0_finish_valid,
    input [1:0] io_clients_0_finish_bits_header_src,
    input [1:0] io_clients_0_finish_bits_header_dst,
    input [2:0] io_clients_0_finish_bits_payload_master_xact_id,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[1:0] io_clients_0_probe_bits_header_src,
    output[1:0] io_clients_0_probe_bits_header_dst,
    output[25:0] io_clients_0_probe_bits_payload_addr,
    output[2:0] io_clients_0_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_0_probe_bits_payload_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_header_src,
    input [1:0] io_clients_0_release_bits_header_dst,
    input [25:0] io_clients_0_release_bits_payload_addr,
    input [1:0] io_clients_0_release_bits_payload_client_xact_id,
    input [2:0] io_clients_0_release_bits_payload_master_xact_id,
    input [511:0] io_clients_0_release_bits_payload_data,
    input [2:0] io_clients_0_release_bits_payload_r_type,
    input  io_masters_0_acquire_ready,
    output io_masters_0_acquire_valid,
    output[1:0] io_masters_0_acquire_bits_header_src,
    output[1:0] io_masters_0_acquire_bits_header_dst,
    output[25:0] io_masters_0_acquire_bits_payload_addr,
    output[1:0] io_masters_0_acquire_bits_payload_client_xact_id,
    output[511:0] io_masters_0_acquire_bits_payload_data,
    output[2:0] io_masters_0_acquire_bits_payload_a_type,
    output[5:0] io_masters_0_acquire_bits_payload_write_mask,
    output[2:0] io_masters_0_acquire_bits_payload_subword_addr,
    output[3:0] io_masters_0_acquire_bits_payload_atomic_opcode,
    output io_masters_0_grant_ready,
    input  io_masters_0_grant_valid,
    input [1:0] io_masters_0_grant_bits_header_src,
    input [1:0] io_masters_0_grant_bits_header_dst,
    input [511:0] io_masters_0_grant_bits_payload_data,
    input [1:0] io_masters_0_grant_bits_payload_client_xact_id,
    input [2:0] io_masters_0_grant_bits_payload_master_xact_id,
    input [3:0] io_masters_0_grant_bits_payload_g_type,
    input  io_masters_0_finish_ready,
    output io_masters_0_finish_valid,
    output[1:0] io_masters_0_finish_bits_header_src,
    output[1:0] io_masters_0_finish_bits_header_dst,
    output[2:0] io_masters_0_finish_bits_payload_master_xact_id,
    output io_masters_0_probe_ready,
    input  io_masters_0_probe_valid,
    input [1:0] io_masters_0_probe_bits_header_src,
    input [1:0] io_masters_0_probe_bits_header_dst,
    input [25:0] io_masters_0_probe_bits_payload_addr,
    input [2:0] io_masters_0_probe_bits_payload_master_xact_id,
    input [1:0] io_masters_0_probe_bits_payload_p_type,
    input  io_masters_0_release_ready,
    output io_masters_0_release_valid,
    output[1:0] io_masters_0_release_bits_header_src,
    output[1:0] io_masters_0_release_bits_header_dst,
    output[25:0] io_masters_0_release_bits_payload_addr,
    output[1:0] io_masters_0_release_bits_payload_client_xact_id,
    output[2:0] io_masters_0_release_bits_payload_master_xact_id,
    output[511:0] io_masters_0_release_bits_payload_data,
    output[2:0] io_masters_0_release_bits_payload_r_type
);

  wire T63;
  wire[2:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[2:0] T69;
  wire[1:0] T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[3:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire[511:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[2:0] T87;
  wire[25:0] T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[511:0] T95;
  wire[2:0] T96;
  wire[1:0] T97;
  wire[25:0] T98;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire[2:0] T103;
  wire[511:0] T104;
  wire[2:0] T105;
  wire[1:0] T106;
  wire[25:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire[1:0] T110;
  wire T111;
  wire T112;
  wire[3:0] T113;
  wire[2:0] T114;
  wire[5:0] T115;
  wire[2:0] T116;
  wire[511:0] T117;
  wire[1:0] T118;
  wire[25:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire[3:0] T124;
  wire[2:0] T125;
  wire[5:0] T126;
  wire[2:0] T127;
  wire[511:0] T128;
  wire[1:0] T129;
  wire[25:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire T134;
  wire[2:0] T0;
  wire[511:0] T1;
  wire[2:0] T2;
  wire[1:0] T3;
  wire[25:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire[2:0] T17;
  wire[5:0] T18;
  wire[2:0] T19;
  wire[511:0] T20;
  wire[1:0] T21;
  wire[25:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire[2:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire[2:0] T37;
  wire[1:0] T38;
  wire[511:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[2:0] T47;
  wire[25:0] T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[3:0] T54;
  wire[2:0] T55;
  wire[1:0] T56;
  wire[511:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire acqNet_io_in_2_ready;
  wire acqNet_io_in_1_ready;
  wire acqNet_io_out_0_valid;
  wire[1:0] acqNet_io_out_0_bits_header_src;
  wire[1:0] acqNet_io_out_0_bits_header_dst;
  wire[25:0] acqNet_io_out_0_bits_payload_addr;
  wire[1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[511:0] acqNet_io_out_0_bits_payload_data;
  wire[2:0] acqNet_io_out_0_bits_payload_a_type;
  wire[5:0] acqNet_io_out_0_bits_payload_write_mask;
  wire[2:0] acqNet_io_out_0_bits_payload_subword_addr;
  wire[3:0] acqNet_io_out_0_bits_payload_atomic_opcode;
  wire relNet_io_in_2_ready;
  wire relNet_io_in_1_ready;
  wire relNet_io_out_0_valid;
  wire[1:0] relNet_io_out_0_bits_header_src;
  wire[1:0] relNet_io_out_0_bits_header_dst;
  wire[25:0] relNet_io_out_0_bits_payload_addr;
  wire[1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire[2:0] relNet_io_out_0_bits_payload_master_xact_id;
  wire[511:0] relNet_io_out_0_bits_payload_data;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire prbNet_io_in_0_ready;
  wire prbNet_io_out_2_valid;
  wire[1:0] prbNet_io_out_2_bits_header_src;
  wire[1:0] prbNet_io_out_2_bits_header_dst;
  wire[25:0] prbNet_io_out_2_bits_payload_addr;
  wire[2:0] prbNet_io_out_2_bits_payload_master_xact_id;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire prbNet_io_out_1_valid;
  wire[1:0] prbNet_io_out_1_bits_header_src;
  wire[1:0] prbNet_io_out_1_bits_header_dst;
  wire[25:0] prbNet_io_out_1_bits_payload_addr;
  wire[2:0] prbNet_io_out_1_bits_payload_master_xact_id;
  wire[1:0] prbNet_io_out_1_bits_payload_p_type;
  wire gntNet_io_in_0_ready;
  wire gntNet_io_out_2_valid;
  wire[1:0] gntNet_io_out_2_bits_header_src;
  wire[1:0] gntNet_io_out_2_bits_header_dst;
  wire[511:0] gntNet_io_out_2_bits_payload_data;
  wire[1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[2:0] gntNet_io_out_2_bits_payload_master_xact_id;
  wire[3:0] gntNet_io_out_2_bits_payload_g_type;
  wire gntNet_io_out_1_valid;
  wire[1:0] gntNet_io_out_1_bits_header_src;
  wire[1:0] gntNet_io_out_1_bits_header_dst;
  wire[511:0] gntNet_io_out_1_bits_payload_data;
  wire[1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire[2:0] gntNet_io_out_1_bits_payload_master_xact_id;
  wire[3:0] gntNet_io_out_1_bits_payload_g_type;
  wire ackNet_io_in_2_ready;
  wire ackNet_io_in_1_ready;
  wire ackNet_io_out_0_valid;
  wire[1:0] ackNet_io_out_0_bits_header_src;
  wire[1:0] ackNet_io_out_0_bits_header_dst;
  wire[2:0] ackNet_io_out_0_bits_payload_master_xact_id;


  assign T63 = io_masters_0_finish_ready;
  assign T64 = io_clients_0_finish_bits_payload_master_xact_id;
  assign T65 = io_clients_0_finish_bits_header_dst;
  assign T66 = T67;
  assign T67 = io_clients_0_finish_bits_header_src + 2'h1;
  assign T68 = io_clients_0_finish_valid;
  assign T69 = io_clients_1_finish_bits_payload_master_xact_id;
  assign T70 = io_clients_1_finish_bits_header_dst;
  assign T71 = T72;
  assign T72 = io_clients_1_finish_bits_header_src + 2'h1;
  assign T73 = io_clients_1_finish_valid;
  assign T74 = io_clients_0_grant_ready;
  assign T75 = io_clients_1_grant_ready;
  assign T76 = io_masters_0_grant_bits_payload_g_type;
  assign T77 = io_masters_0_grant_bits_payload_master_xact_id;
  assign T78 = io_masters_0_grant_bits_payload_client_xact_id;
  assign T79 = io_masters_0_grant_bits_payload_data;
  assign T80 = T81;
  assign T81 = io_masters_0_grant_bits_header_dst + 2'h1;
  assign T82 = io_masters_0_grant_bits_header_src;
  assign T83 = io_masters_0_grant_valid;
  assign T84 = io_clients_0_probe_ready;
  assign T85 = io_clients_1_probe_ready;
  assign T86 = io_masters_0_probe_bits_payload_p_type;
  assign T87 = io_masters_0_probe_bits_payload_master_xact_id;
  assign T88 = io_masters_0_probe_bits_payload_addr;
  assign T89 = T90;
  assign T90 = io_masters_0_probe_bits_header_dst + 2'h1;
  assign T91 = io_masters_0_probe_bits_header_src;
  assign T92 = io_masters_0_probe_valid;
  assign T93 = io_masters_0_release_ready;
  assign T94 = io_clients_0_release_bits_payload_r_type;
  assign T95 = io_clients_0_release_bits_payload_data;
  assign T96 = io_clients_0_release_bits_payload_master_xact_id;
  assign T97 = io_clients_0_release_bits_payload_client_xact_id;
  assign T98 = io_clients_0_release_bits_payload_addr;
  assign T99 = io_clients_0_release_bits_header_dst;
  assign T100 = T101;
  assign T101 = io_clients_0_release_bits_header_src + 2'h1;
  assign T102 = io_clients_0_release_valid;
  assign T103 = io_clients_1_release_bits_payload_r_type;
  assign T104 = io_clients_1_release_bits_payload_data;
  assign T105 = io_clients_1_release_bits_payload_master_xact_id;
  assign T106 = io_clients_1_release_bits_payload_client_xact_id;
  assign T107 = io_clients_1_release_bits_payload_addr;
  assign T108 = io_clients_1_release_bits_header_dst;
  assign T109 = T110;
  assign T110 = io_clients_1_release_bits_header_src + 2'h1;
  assign T111 = io_clients_1_release_valid;
  assign T112 = io_masters_0_acquire_ready;
  assign T113 = io_clients_0_acquire_bits_payload_atomic_opcode;
  assign T114 = io_clients_0_acquire_bits_payload_subword_addr;
  assign T115 = io_clients_0_acquire_bits_payload_write_mask;
  assign T116 = io_clients_0_acquire_bits_payload_a_type;
  assign T117 = io_clients_0_acquire_bits_payload_data;
  assign T118 = io_clients_0_acquire_bits_payload_client_xact_id;
  assign T119 = io_clients_0_acquire_bits_payload_addr;
  assign T120 = io_clients_0_acquire_bits_header_dst;
  assign T121 = T122;
  assign T122 = io_clients_0_acquire_bits_header_src + 2'h1;
  assign T123 = io_clients_0_acquire_valid;
  assign T124 = io_clients_1_acquire_bits_payload_atomic_opcode;
  assign T125 = io_clients_1_acquire_bits_payload_subword_addr;
  assign T126 = io_clients_1_acquire_bits_payload_write_mask;
  assign T127 = io_clients_1_acquire_bits_payload_a_type;
  assign T128 = io_clients_1_acquire_bits_payload_data;
  assign T129 = io_clients_1_acquire_bits_payload_client_xact_id;
  assign T130 = io_clients_1_acquire_bits_payload_addr;
  assign T131 = io_clients_1_acquire_bits_header_dst;
  assign T132 = T133;
  assign T133 = io_clients_1_acquire_bits_header_src + 2'h1;
  assign T134 = io_clients_1_acquire_valid;
  assign io_masters_0_release_bits_payload_r_type = T0;
  assign T0 = relNet_io_out_0_bits_payload_r_type;
  assign io_masters_0_release_bits_payload_data = T1;
  assign T1 = relNet_io_out_0_bits_payload_data;
  assign io_masters_0_release_bits_payload_master_xact_id = T2;
  assign T2 = relNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_release_bits_payload_client_xact_id = T3;
  assign T3 = relNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_release_bits_payload_addr = T4;
  assign T4 = relNet_io_out_0_bits_payload_addr;
  assign io_masters_0_release_bits_header_dst = T5;
  assign T5 = relNet_io_out_0_bits_header_dst;
  assign io_masters_0_release_bits_header_src = T6;
  assign T6 = T7;
  assign T7 = relNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_release_valid = T8;
  assign T8 = relNet_io_out_0_valid;
  assign io_masters_0_probe_ready = T9;
  assign T9 = prbNet_io_in_0_ready;
  assign io_masters_0_finish_bits_payload_master_xact_id = T10;
  assign T10 = ackNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_finish_bits_header_dst = T11;
  assign T11 = ackNet_io_out_0_bits_header_dst;
  assign io_masters_0_finish_bits_header_src = T12;
  assign T12 = T13;
  assign T13 = ackNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_finish_valid = T14;
  assign T14 = ackNet_io_out_0_valid;
  assign io_masters_0_grant_ready = T15;
  assign T15 = gntNet_io_in_0_ready;
  assign io_masters_0_acquire_bits_payload_atomic_opcode = T16;
  assign T16 = acqNet_io_out_0_bits_payload_atomic_opcode;
  assign io_masters_0_acquire_bits_payload_subword_addr = T17;
  assign T17 = acqNet_io_out_0_bits_payload_subword_addr;
  assign io_masters_0_acquire_bits_payload_write_mask = T18;
  assign T18 = acqNet_io_out_0_bits_payload_write_mask;
  assign io_masters_0_acquire_bits_payload_a_type = T19;
  assign T19 = acqNet_io_out_0_bits_payload_a_type;
  assign io_masters_0_acquire_bits_payload_data = T20;
  assign T20 = acqNet_io_out_0_bits_payload_data;
  assign io_masters_0_acquire_bits_payload_client_xact_id = T21;
  assign T21 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_acquire_bits_payload_addr = T22;
  assign T22 = acqNet_io_out_0_bits_payload_addr;
  assign io_masters_0_acquire_bits_header_dst = T23;
  assign T23 = acqNet_io_out_0_bits_header_dst;
  assign io_masters_0_acquire_bits_header_src = T24;
  assign T24 = T25;
  assign T25 = acqNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_acquire_valid = T26;
  assign T26 = acqNet_io_out_0_valid;
  assign io_clients_0_release_ready = T27;
  assign T27 = relNet_io_in_1_ready;
  assign io_clients_0_probe_bits_payload_p_type = T28;
  assign T28 = prbNet_io_out_1_bits_payload_p_type;
  assign io_clients_0_probe_bits_payload_master_xact_id = T29;
  assign T29 = prbNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_probe_bits_payload_addr = T30;
  assign T30 = prbNet_io_out_1_bits_payload_addr;
  assign io_clients_0_probe_bits_header_dst = T31;
  assign T31 = T32;
  assign T32 = prbNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_probe_bits_header_src = T33;
  assign T33 = prbNet_io_out_1_bits_header_src;
  assign io_clients_0_probe_valid = T34;
  assign T34 = prbNet_io_out_1_valid;
  assign io_clients_0_finish_ready = T35;
  assign T35 = ackNet_io_in_1_ready;
  assign io_clients_0_grant_bits_payload_g_type = T36;
  assign T36 = gntNet_io_out_1_bits_payload_g_type;
  assign io_clients_0_grant_bits_payload_master_xact_id = T37;
  assign T37 = gntNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_grant_bits_payload_client_xact_id = T38;
  assign T38 = gntNet_io_out_1_bits_payload_client_xact_id;
  assign io_clients_0_grant_bits_payload_data = T39;
  assign T39 = gntNet_io_out_1_bits_payload_data;
  assign io_clients_0_grant_bits_header_dst = T40;
  assign T40 = T41;
  assign T41 = gntNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_grant_bits_header_src = T42;
  assign T42 = gntNet_io_out_1_bits_header_src;
  assign io_clients_0_grant_valid = T43;
  assign T43 = gntNet_io_out_1_valid;
  assign io_clients_0_acquire_ready = T44;
  assign T44 = acqNet_io_in_1_ready;
  assign io_clients_1_release_ready = T45;
  assign T45 = relNet_io_in_2_ready;
  assign io_clients_1_probe_bits_payload_p_type = T46;
  assign T46 = prbNet_io_out_2_bits_payload_p_type;
  assign io_clients_1_probe_bits_payload_master_xact_id = T47;
  assign T47 = prbNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_probe_bits_payload_addr = T48;
  assign T48 = prbNet_io_out_2_bits_payload_addr;
  assign io_clients_1_probe_bits_header_dst = T49;
  assign T49 = T50;
  assign T50 = prbNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_probe_bits_header_src = T51;
  assign T51 = prbNet_io_out_2_bits_header_src;
  assign io_clients_1_probe_valid = T52;
  assign T52 = prbNet_io_out_2_valid;
  assign io_clients_1_finish_ready = T53;
  assign T53 = ackNet_io_in_2_ready;
  assign io_clients_1_grant_bits_payload_g_type = T54;
  assign T54 = gntNet_io_out_2_bits_payload_g_type;
  assign io_clients_1_grant_bits_payload_master_xact_id = T55;
  assign T55 = gntNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_grant_bits_payload_client_xact_id = T56;
  assign T56 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign io_clients_1_grant_bits_payload_data = T57;
  assign T57 = gntNet_io_out_2_bits_payload_data;
  assign io_clients_1_grant_bits_header_dst = T58;
  assign T58 = T59;
  assign T59 = gntNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_grant_bits_header_src = T60;
  assign T60 = gntNet_io_out_2_bits_header_src;
  assign io_clients_1_grant_valid = T61;
  assign T61 = gntNet_io_out_2_valid;
  assign io_clients_1_acquire_ready = T62;
  assign T62 = acqNet_io_in_2_ready;
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T134 ),
       .io_in_2_bits_header_src( T132 ),
       .io_in_2_bits_header_dst( T131 ),
       .io_in_2_bits_payload_addr( T130 ),
       .io_in_2_bits_payload_client_xact_id( T129 ),
       .io_in_2_bits_payload_data( T128 ),
       .io_in_2_bits_payload_a_type( T127 ),
       .io_in_2_bits_payload_write_mask( T126 ),
       .io_in_2_bits_payload_subword_addr( T125 ),
       .io_in_2_bits_payload_atomic_opcode( T124 ),
       .io_in_1_ready( acqNet_io_in_1_ready ),
       .io_in_1_valid( T123 ),
       .io_in_1_bits_header_src( T121 ),
       .io_in_1_bits_header_dst( T120 ),
       .io_in_1_bits_payload_addr( T119 ),
       .io_in_1_bits_payload_client_xact_id( T118 ),
       .io_in_1_bits_payload_data( T117 ),
       .io_in_1_bits_payload_a_type( T116 ),
       .io_in_1_bits_payload_write_mask( T115 ),
       .io_in_1_bits_payload_subword_addr( T114 ),
       .io_in_1_bits_payload_atomic_opcode( T113 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_write_mask(  )
       //.io_in_0_bits_payload_subword_addr(  )
       //.io_in_0_bits_payload_atomic_opcode(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_write_mask(  )
       //.io_out_2_bits_payload_subword_addr(  )
       //.io_out_2_bits_payload_atomic_opcode(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_a_type(  )
       //.io_out_1_bits_payload_write_mask(  )
       //.io_out_1_bits_payload_subword_addr(  )
       //.io_out_1_bits_payload_atomic_opcode(  )
       .io_out_0_ready( T112 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( acqNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_write_mask( acqNet_io_out_0_bits_payload_write_mask ),
       .io_out_0_bits_payload_subword_addr( acqNet_io_out_0_bits_payload_subword_addr ),
       .io_out_0_bits_payload_atomic_opcode( acqNet_io_out_0_bits_payload_atomic_opcode )
  );
  `ifndef SYNTHESIS
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {16{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_write_mask = {1{$random}};
    assign acqNet.io_in_0_bits_payload_subword_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_atomic_opcode = {1{$random}};
  `endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T111 ),
       .io_in_2_bits_header_src( T109 ),
       .io_in_2_bits_header_dst( T108 ),
       .io_in_2_bits_payload_addr( T107 ),
       .io_in_2_bits_payload_client_xact_id( T106 ),
       .io_in_2_bits_payload_master_xact_id( T105 ),
       .io_in_2_bits_payload_data( T104 ),
       .io_in_2_bits_payload_r_type( T103 ),
       .io_in_1_ready( relNet_io_in_1_ready ),
       .io_in_1_valid( T102 ),
       .io_in_1_bits_header_src( T100 ),
       .io_in_1_bits_header_dst( T99 ),
       .io_in_1_bits_payload_addr( T98 ),
       .io_in_1_bits_payload_client_xact_id( T97 ),
       .io_in_1_bits_payload_master_xact_id( T96 ),
       .io_in_1_bits_payload_data( T95 ),
       .io_in_1_bits_payload_r_type( T94 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_r_type(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_r_type(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_r_type(  )
       .io_out_0_ready( T93 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( relNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_master_xact_id( relNet_io_out_0_bits_payload_master_xact_id ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type )
  );
  `ifndef SYNTHESIS
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {16{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
  `endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_p_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_p_type(  )
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T92 ),
       .io_in_0_bits_header_src( T91 ),
       .io_in_0_bits_header_dst( T89 ),
       .io_in_0_bits_payload_addr( T88 ),
       .io_in_0_bits_payload_master_xact_id( T87 ),
       .io_in_0_bits_payload_p_type( T86 ),
       .io_out_2_ready( T85 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr( prbNet_io_out_2_bits_payload_addr ),
       .io_out_2_bits_payload_master_xact_id( prbNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( T84 ),
       .io_out_1_valid( prbNet_io_out_1_valid ),
       .io_out_1_bits_header_src( prbNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( prbNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr( prbNet_io_out_1_bits_payload_addr ),
       .io_out_1_bits_payload_master_xact_id( prbNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_p_type( prbNet_io_out_1_bits_payload_p_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_p_type(  )
  );
  `ifndef SYNTHESIS
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_1_bits_header_src = {1{$random}};
    assign prbNet.io_in_1_bits_header_dst = {1{$random}};
    assign prbNet.io_in_1_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_1_bits_payload_p_type = {1{$random}};
  `endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_data(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_g_type(  )
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T83 ),
       .io_in_0_bits_header_src( T82 ),
       .io_in_0_bits_header_dst( T80 ),
       .io_in_0_bits_payload_data( T79 ),
       .io_in_0_bits_payload_client_xact_id( T78 ),
       .io_in_0_bits_payload_master_xact_id( T77 ),
       .io_in_0_bits_payload_g_type( T76 ),
       .io_out_2_ready( T75 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_master_xact_id( gntNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_1_ready( T74 ),
       .io_out_1_valid( gntNet_io_out_1_valid ),
       .io_out_1_bits_header_src( gntNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( gntNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_data( gntNet_io_out_1_bits_payload_data ),
       .io_out_1_bits_payload_client_xact_id( gntNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_master_xact_id( gntNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_g_type( gntNet_io_out_1_bits_payload_g_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_data(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_g_type(  )
  );
  `ifndef SYNTHESIS
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {16{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_1_bits_header_src = {1{$random}};
    assign gntNet.io_in_1_bits_header_dst = {1{$random}};
    assign gntNet.io_in_1_bits_payload_data = {16{$random}};
    assign gntNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_g_type = {1{$random}};
  `endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T73 ),
       .io_in_2_bits_header_src( T71 ),
       .io_in_2_bits_header_dst( T70 ),
       .io_in_2_bits_payload_master_xact_id( T69 ),
       .io_in_1_ready( ackNet_io_in_1_ready ),
       .io_in_1_valid( T68 ),
       .io_in_1_bits_header_src( T66 ),
       .io_in_1_bits_header_dst( T65 ),
       .io_in_1_bits_payload_master_xact_id( T64 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       .io_out_0_ready( T63 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_master_xact_id( ackNet_io_out_0_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module VoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[1:0] io_inner_probe_bits_header_src
    //output[1:0] io_inner_probe_bits_header_dst
    //output[25:0] io_inner_probe_bits_payload_addr
    //output[2:0] io_inner_probe_bits_payload_master_xact_id
    //output[1:0] io_inner_probe_bits_payload_p_type
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T38;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [25:0] xact_addr;
  wire[25:0] T20;
  wire[3:0] T21;
  wire[2:0] T22;
  wire[5:0] T23;
  wire[2:0] T24;
  wire[511:0] T25;
  reg [511:0] xact_data;
  wire[511:0] T26;
  wire[2:0] T27;
  wire[25:0] T28;
  wire[3:0] T29;
  wire[3:0] T30;
  wire T31;
  reg [2:0] xact_r_type;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[1:0] T34;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T35;
  wire[511:0] T36;
  wire[1:0] T39;
  reg  init_client_id;
  wire T40;
  wire[1:0] T41;
  wire[1:0] T37;
  wire[1:0] T42;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    xact_r_type = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T19 & T1;
  assign T1 = state != 2'h0;
  assign T38 = reset ? 2'h0 : T2;
  assign T2 = T17 ? 2'h0 : T3;
  assign T3 = T15 ? 2'h2 : T4;
  assign T4 = T13 ? T5 : state;
  assign T5 = T6 ? 2'h1 : 2'h2;
  assign T6 = T8 | T7;
  assign T7 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T8 = T10 | T9;
  assign T9 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T10 = T12 | T11;
  assign T11 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T12 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T13 = T14 & io_inner_release_valid;
  assign T14 = 2'h0 == state;
  assign T15 = T16 & io_outer_acquire_ready;
  assign T16 = 2'h1 == state;
  assign T17 = T18 & io_inner_grant_ready;
  assign T18 = 2'h2 == state;
  assign T19 = xact_addr == io_inner_release_bits_payload_addr;
  assign T20 = T13 ? io_inner_release_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = 1'h0;
  assign io_outer_acquire_bits_payload_atomic_opcode = T21;
  assign T21 = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T22;
  assign T22 = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T23;
  assign T23 = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T24;
  assign T24 = 3'h3;
  assign io_outer_acquire_bits_payload_data = T25;
  assign T25 = xact_data;
  assign T26 = T13 ? io_inner_release_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T27;
  assign T27 = 3'h0;
  assign io_outer_acquire_bits_payload_addr = T28;
  assign T28 = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T16;
  assign io_inner_release_ready = T14;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_grant_bits_payload_g_type = T29;
  assign T29 = T30;
  assign T30 = T31 ? 4'h0 : 4'h3;
  assign T31 = xact_r_type == 3'h0;
  assign T32 = T13 ? io_inner_release_bits_payload_r_type : xact_r_type;
  assign io_inner_grant_bits_payload_master_xact_id = T33;
  assign T33 = 3'h0;
  assign io_inner_grant_bits_payload_client_xact_id = T34;
  assign T34 = xact_client_xact_id;
  assign T35 = T13 ? io_inner_release_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T36;
  assign T36 = 512'h0;
  assign io_inner_grant_bits_header_dst = T39;
  assign T39 = {1'h0, init_client_id};
  assign T40 = T41[1'h0:1'h0];
  assign T41 = reset ? 2'h0 : T37;
  assign T37 = T13 ? io_inner_release_bits_header_src : T42;
  assign T42 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T18;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T17) begin
      state <= 2'h0;
    end else if(T15) begin
      state <= 2'h2;
    end else if(T13) begin
      state <= T5;
    end
    if(T13) begin
      xact_addr <= io_inner_release_bits_payload_addr;
    end
    if(T13) begin
      xact_data <= io_inner_release_bits_payload_data;
    end
    if(T13) begin
      xact_r_type <= io_inner_release_bits_payload_r_type;
    end
    if(T13) begin
      xact_client_xact_id <= io_inner_release_bits_payload_client_xact_id;
    end
    init_client_id <= T40;
  end
endmodule

module AcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h1;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h1;
  assign outer_read_client_xact_id = 3'h1;
  assign outer_write_acq_client_xact_id = 3'h1;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h1;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h1;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h1;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module AcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h2;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h2;
  assign outer_read_client_xact_id = 3'h2;
  assign outer_write_acq_client_xact_id = 3'h2;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h2;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h2;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h2;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module AcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h3;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h3;
  assign outer_read_client_xact_id = 3'h3;
  assign outer_write_acq_client_xact_id = 3'h3;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h3;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h3;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h3;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module AcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h4;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h4;
  assign outer_read_client_xact_id = 3'h4;
  assign outer_write_acq_client_xact_id = 3'h4;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h4;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h4;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h4;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module AcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h5;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h5;
  assign outer_read_client_xact_id = 3'h5;
  assign outer_write_acq_client_xact_id = 3'h5;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h5;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h5;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h5;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module AcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h6;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h6;
  assign outer_read_client_xact_id = 3'h6;
  assign outer_write_acq_client_xact_id = 3'h6;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h6;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h6;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h6;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module AcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T145;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T146;
  wire[1:0] T147;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T148;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T149;
  wire T38;
  wire[1:0] T150;
  wire T39;
  wire[1:0] T151;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [25:0] xact_addr;
  wire[25:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T100;
  wire[2:0] T101;
  wire[2:0] T102;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T103;
  wire[511:0] T104;
  wire[511:0] T105;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[25:0] T110;
  wire[25:0] T111;
  wire[25:0] T112;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  wire[25:0] T126;
  wire[1:0] T152;
  wire T153;
  wire T154;
  reg [1:0] probe_flags;
  wire[1:0] T155;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[2:0] T136;
  wire[1:0] T137;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T138;
  wire[511:0] T139;
  wire[1:0] T156;
  reg  init_client_id;
  wire T157;
  wire[1:0] T158;
  wire[1:0] T140;
  wire[1:0] T159;
  wire T141;
  wire T142;
  wire T143;
  wire T144;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T86 & T1;
  assign T1 = state != 3'h0;
  assign T145 = reset ? 3'h0 : T2;
  assign T2 = T82 ? 3'h0 : T3;
  assign T3 = T80 ? T78 : T4;
  assign T4 = T76 ? T75 : T5;
  assign T5 = T73 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T146 = T147[1'h0:1'h0];
  assign T147 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T151 : T33;
  assign T33 = T52 ? T150 : T34;
  assign T34 = T21 ? T35 : T148;
  assign T148 = {1'h0, release_count};
  assign T35 = T149 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T149 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T150 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T151 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T72 ? 4'h2 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = xact_a_type == 3'h0;
  assign T73 = T74 & io_outer_acquire_ready;
  assign T74 = 3'h2 == state;
  assign T75 = pending_outer_read ? 3'h2 : 3'h4;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h3 == state;
  assign T78 = T79 ? 3'h5 : 3'h0;
  assign T79 = grant_type != 4'h0;
  assign T80 = T81 & io_inner_grant_ready;
  assign T81 = 3'h4 == state;
  assign T82 = T85 & T83;
  assign T83 = io_inner_finish_valid & T84;
  assign T84 = io_inner_finish_bits_payload_master_xact_id == 3'h7;
  assign T85 = 3'h5 == state;
  assign T86 = xact_addr == io_inner_release_bits_payload_addr;
  assign T87 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T88;
  assign T88 = T90 & T89;
  assign T89 = state != 3'h0;
  assign T90 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T91;
  assign T91 = T77 ? outer_write_acq_atomic_opcode : T92;
  assign T92 = T74 ? outer_read_atomic_opcode : T93;
  assign T93 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T94;
  assign T94 = T77 ? outer_write_acq_subword_addr : T95;
  assign T95 = T74 ? outer_read_subword_addr : T96;
  assign T96 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T97;
  assign T97 = T77 ? outer_write_acq_write_mask : T98;
  assign T98 = T74 ? outer_read_write_mask : T99;
  assign T99 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T100;
  assign T100 = T77 ? outer_write_acq_a_type : T101;
  assign T101 = T74 ? outer_read_a_type : T102;
  assign T102 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T103;
  assign T103 = T77 ? outer_write_acq_data : T104;
  assign T104 = T74 ? outer_read_data : T105;
  assign T105 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T106 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T107;
  assign T107 = T77 ? outer_write_acq_client_xact_id : T108;
  assign T108 = T74 ? outer_read_client_xact_id : T109;
  assign T109 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h7;
  assign outer_read_client_xact_id = 3'h7;
  assign outer_write_acq_client_xact_id = 3'h7;
  assign io_outer_acquire_bits_payload_addr = T110;
  assign T110 = T77 ? outer_write_acq_addr : T111;
  assign T111 = T74 ? outer_read_addr : T112;
  assign T112 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T113;
  assign T113 = T77 ? 1'h1 : T114;
  assign T114 = T74 ? 1'h1 : T53;
  assign io_inner_release_ready = T115;
  assign T115 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T116;
  assign T116 = T117;
  assign T117 = T124 ? 2'h1 : T118;
  assign T118 = T123 ? 2'h0 : T119;
  assign T119 = T122 ? 2'h2 : T120;
  assign T120 = T121 ? 2'h0 : 2'h2;
  assign T121 = xact_a_type == 3'h3;
  assign T122 = xact_a_type == 3'h2;
  assign T123 = xact_a_type == 3'h1;
  assign T124 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T125;
  assign T125 = 3'h7;
  assign io_inner_probe_bits_payload_addr = T126;
  assign T126 = xact_addr;
  assign io_inner_probe_bits_header_dst = T152;
  assign T152 = {1'h0, T153};
  assign T153 = T154 == 1'h0;
  assign T154 = probe_flags[1'h0:1'h0];
  assign T155 = reset ? 2'h0 : T127;
  assign T127 = T132 ? T129 : T128;
  assign T128 = T21 ? probe_initial_flags : probe_flags;
  assign T129 = probe_flags & T130;
  assign T130 = ~ T131;
  assign T131 = 1'h1 << T153;
  assign T132 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T133;
  assign T133 = T51 ? T134 : 1'h0;
  assign T134 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T135;
  assign T135 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T136;
  assign T136 = 3'h7;
  assign io_inner_grant_bits_payload_client_xact_id = T137;
  assign T137 = xact_client_xact_id;
  assign T138 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T139;
  assign T139 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T156;
  assign T156 = {1'h0, init_client_id};
  assign T157 = T158[1'h0:1'h0];
  assign T158 = reset ? 2'h0 : T140;
  assign T140 = T21 ? io_inner_acquire_bits_header_src : T159;
  assign T159 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T141;
  assign T141 = T142 ? 1'h1 : T81;
  assign T142 = T85 & T143;
  assign T143 = io_outer_grant_valid & T144;
  assign T144 = io_outer_grant_bits_payload_client_xact_id == 3'h7;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T146;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T132) begin
      probe_flags <= T129;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T157;
  end
endmodule

module Arbiter_11(
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits : io_in_0_bits;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits : io_in_2_bits;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits : io_in_4_bits;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits : io_in_6_bits;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_valid = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_valid : io_in_0_valid;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_valid : io_in_4_valid;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_valid : io_in_6_valid;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T41 ^ 1'h1;
  assign T41 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T45 | io_in_2_valid;
  assign T45 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T46;
  assign T46 = T47 & io_out_ready;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T49 | io_in_3_valid;
  assign T49 = T50 | io_in_2_valid;
  assign T50 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T54 | io_in_4_valid;
  assign T54 = T55 | io_in_3_valid;
  assign T55 = T56 | io_in_2_valid;
  assign T56 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_5_valid;
  assign T60 = T61 | io_in_4_valid;
  assign T61 = T62 | io_in_3_valid;
  assign T62 = T63 | io_in_2_valid;
  assign T63 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_6_valid;
  assign T67 = T68 | io_in_5_valid;
  assign T68 = T69 | io_in_4_valid;
  assign T69 = T70 | io_in_3_valid;
  assign T70 = T71 | io_in_2_valid;
  assign T71 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_12(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input [1:0] io_in_7_bits_payload_p_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input [1:0] io_in_6_bits_payload_p_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input [1:0] io_in_5_bits_payload_p_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[25:0] T37;
  wire[25:0] T38;
  wire[25:0] T39;
  wire T40;
  wire[25:0] T41;
  wire T42;
  wire T43;
  wire[25:0] T44;
  wire[25:0] T45;
  wire T46;
  wire[25:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_p_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_p_type : io_in_4_bits_payload_p_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_p_type : io_in_6_bits_payload_p_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_addr = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_valid = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_valid : io_in_0_valid;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_valid : io_in_4_valid;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_valid : io_in_6_valid;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T95;
  assign T95 = T96 & io_out_ready;
  assign T96 = T97 ^ 1'h1;
  assign T97 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T98;
  assign T98 = T99 & io_out_ready;
  assign T99 = T100 ^ 1'h1;
  assign T100 = T101 | io_in_2_valid;
  assign T101 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T102;
  assign T102 = T103 & io_out_ready;
  assign T103 = T104 ^ 1'h1;
  assign T104 = T105 | io_in_3_valid;
  assign T105 = T106 | io_in_2_valid;
  assign T106 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T110 | io_in_4_valid;
  assign T110 = T111 | io_in_3_valid;
  assign T111 = T112 | io_in_2_valid;
  assign T112 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T113;
  assign T113 = T114 & io_out_ready;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T116 | io_in_5_valid;
  assign T116 = T117 | io_in_4_valid;
  assign T117 = T118 | io_in_3_valid;
  assign T118 = T119 | io_in_2_valid;
  assign T119 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T120;
  assign T120 = T121 & io_out_ready;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T123 | io_in_6_valid;
  assign T123 = T124 | io_in_5_valid;
  assign T124 = T125 | io_in_4_valid;
  assign T125 = T126 | io_in_3_valid;
  assign T126 = T127 | io_in_2_valid;
  assign T127 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_13(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [511:0] io_in_7_bits_payload_data,
    input [1:0] io_in_7_bits_payload_client_xact_id,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input [3:0] io_in_7_bits_payload_g_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [511:0] io_in_6_bits_payload_data,
    input [1:0] io_in_6_bits_payload_client_xact_id,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input [3:0] io_in_6_bits_payload_g_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [511:0] io_in_5_bits_payload_data,
    input [1:0] io_in_5_bits_payload_client_xact_id,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input [3:0] io_in_5_bits_payload_g_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [511:0] io_in_4_bits_payload_data,
    input [1:0] io_in_4_bits_payload_client_xact_id,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input [3:0] io_in_4_bits_payload_g_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [511:0] io_in_3_bits_payload_data,
    input [1:0] io_in_3_bits_payload_client_xact_id,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input [3:0] io_in_3_bits_payload_g_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[511:0] T51;
  wire[511:0] T52;
  wire[511:0] T53;
  wire T54;
  wire[511:0] T55;
  wire T56;
  wire T57;
  wire[511:0] T58;
  wire[511:0] T59;
  wire T60;
  wire[511:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_g_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_g_type : io_in_4_bits_payload_g_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_g_type : io_in_6_bits_payload_g_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_payload_data = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_out_valid = T93;
  assign T93 = T106 ? T100 : T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96 ? io_in_1_valid : io_in_0_valid;
  assign T96 = T12[1'h0:1'h0];
  assign T97 = T98 ? io_in_3_valid : io_in_2_valid;
  assign T98 = T12[1'h0:1'h0];
  assign T99 = T12[1'h1:1'h1];
  assign T100 = T105 ? T103 : T101;
  assign T101 = T102 ? io_in_5_valid : io_in_4_valid;
  assign T102 = T12[1'h0:1'h0];
  assign T103 = T104 ? io_in_7_valid : io_in_6_valid;
  assign T104 = T12[1'h0:1'h0];
  assign T105 = T12[1'h1:1'h1];
  assign T106 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T109;
  assign T109 = T110 & io_out_ready;
  assign T110 = T111 ^ 1'h1;
  assign T111 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T112;
  assign T112 = T113 & io_out_ready;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115 | io_in_2_valid;
  assign T115 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T116;
  assign T116 = T117 & io_out_ready;
  assign T117 = T118 ^ 1'h1;
  assign T118 = T119 | io_in_3_valid;
  assign T119 = T120 | io_in_2_valid;
  assign T120 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T121;
  assign T121 = T122 & io_out_ready;
  assign T122 = T123 ^ 1'h1;
  assign T123 = T124 | io_in_4_valid;
  assign T124 = T125 | io_in_3_valid;
  assign T125 = T126 | io_in_2_valid;
  assign T126 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T127;
  assign T127 = T128 & io_out_ready;
  assign T128 = T129 ^ 1'h1;
  assign T129 = T130 | io_in_5_valid;
  assign T130 = T131 | io_in_4_valid;
  assign T131 = T132 | io_in_3_valid;
  assign T132 = T133 | io_in_2_valid;
  assign T133 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T134;
  assign T134 = T135 & io_out_ready;
  assign T135 = T136 ^ 1'h1;
  assign T136 = T137 | io_in_6_valid;
  assign T137 = T138 | io_in_5_valid;
  assign T138 = T139 | io_in_4_valid;
  assign T139 = T140 | io_in_3_valid;
  assign T140 = T141 | io_in_2_valid;
  assign T141 = io_in_0_valid | io_in_1_valid;
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [2:0] io_in_7_bits_payload_client_xact_id,
    input [511:0] io_in_7_bits_payload_data,
    input [2:0] io_in_7_bits_payload_a_type,
    input [5:0] io_in_7_bits_payload_write_mask,
    input [2:0] io_in_7_bits_payload_subword_addr,
    input [3:0] io_in_7_bits_payload_atomic_opcode,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [2:0] io_in_6_bits_payload_client_xact_id,
    input [511:0] io_in_6_bits_payload_data,
    input [2:0] io_in_6_bits_payload_a_type,
    input [5:0] io_in_6_bits_payload_write_mask,
    input [2:0] io_in_6_bits_payload_subword_addr,
    input [3:0] io_in_6_bits_payload_atomic_opcode,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [2:0] io_in_5_bits_payload_client_xact_id,
    input [511:0] io_in_5_bits_payload_data,
    input [2:0] io_in_5_bits_payload_a_type,
    input [5:0] io_in_5_bits_payload_write_mask,
    input [2:0] io_in_5_bits_payload_subword_addr,
    input [3:0] io_in_5_bits_payload_atomic_opcode,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [2:0] io_in_4_bits_payload_client_xact_id,
    input [511:0] io_in_4_bits_payload_data,
    input [2:0] io_in_4_bits_payload_a_type,
    input [5:0] io_in_4_bits_payload_write_mask,
    input [2:0] io_in_4_bits_payload_subword_addr,
    input [3:0] io_in_4_bits_payload_atomic_opcode,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [2:0] io_in_3_bits_payload_client_xact_id,
    input [511:0] io_in_3_bits_payload_data,
    input [2:0] io_in_3_bits_payload_a_type,
    input [5:0] io_in_3_bits_payload_write_mask,
    input [2:0] io_in_3_bits_payload_subword_addr,
    input [3:0] io_in_3_bits_payload_atomic_opcode,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T340;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire[3:0] T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[2:0] T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire[2:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire T64;
  wire[5:0] T65;
  wire T66;
  wire T67;
  wire[5:0] T68;
  wire[5:0] T69;
  wire T70;
  wire[5:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire T78;
  wire[2:0] T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[2:0] T83;
  wire T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[511:0] T89;
  wire[511:0] T90;
  wire[511:0] T91;
  wire T92;
  wire[511:0] T93;
  wire T94;
  wire T95;
  wire[511:0] T96;
  wire[511:0] T97;
  wire T98;
  wire[511:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire T106;
  wire[2:0] T107;
  wire T108;
  wire T109;
  wire[2:0] T110;
  wire[2:0] T111;
  wire T112;
  wire[2:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[25:0] T117;
  wire[25:0] T118;
  wire[25:0] T119;
  wire T120;
  wire[25:0] T121;
  wire T122;
  wire T123;
  wire[25:0] T124;
  wire[25:0] T125;
  wire T126;
  wire[25:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire T140;
  wire[1:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[1:0] T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire T148;
  wire[1:0] T149;
  wire T150;
  wire T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T30 ? 3'h1 : T2;
  assign T2 = T28 ? 3'h2 : T3;
  assign T3 = T26 ? 3'h3 : T4;
  assign T4 = T24 ? 3'h4 : T5;
  assign T5 = T22 ? 3'h5 : T6;
  assign T6 = T20 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T340 = reset ? 3'h0 : T18;
  assign T18 = T19 ? T0 : R17;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = io_in_6_valid & T21;
  assign T21 = R17 < 3'h6;
  assign T22 = io_in_5_valid & T23;
  assign T23 = R17 < 3'h5;
  assign T24 = io_in_4_valid & T25;
  assign T25 = R17 < 3'h4;
  assign T26 = io_in_3_valid & T27;
  assign T27 = R17 < 3'h3;
  assign T28 = io_in_2_valid & T29;
  assign T29 = R17 < 3'h2;
  assign T30 = io_in_1_valid & T31;
  assign T31 = R17 < 3'h1;
  assign io_out_bits_payload_atomic_opcode = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = T0;
  assign T37 = T38 ? io_in_3_bits_payload_atomic_opcode : io_in_2_bits_payload_atomic_opcode;
  assign T38 = T36[1'h0:1'h0];
  assign T39 = T36[1'h1:1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_payload_atomic_opcode : io_in_4_bits_payload_atomic_opcode;
  assign T42 = T36[1'h0:1'h0];
  assign T43 = T44 ? io_in_7_bits_payload_atomic_opcode : io_in_6_bits_payload_atomic_opcode;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign T46 = T36[2'h2:2'h2];
  assign io_out_bits_payload_subword_addr = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T50 = T36[1'h0:1'h0];
  assign T51 = T52 ? io_in_3_bits_payload_subword_addr : io_in_2_bits_payload_subword_addr;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_payload_subword_addr : io_in_4_bits_payload_subword_addr;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T58 ? io_in_7_bits_payload_subword_addr : io_in_6_bits_payload_subword_addr;
  assign T58 = T36[1'h0:1'h0];
  assign T59 = T36[1'h1:1'h1];
  assign T60 = T36[2'h2:2'h2];
  assign io_out_bits_payload_write_mask = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T66 ? io_in_3_bits_payload_write_mask : io_in_2_bits_payload_write_mask;
  assign T66 = T36[1'h0:1'h0];
  assign T67 = T36[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_payload_write_mask : io_in_4_bits_payload_write_mask;
  assign T70 = T36[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_payload_write_mask : io_in_6_bits_payload_write_mask;
  assign T72 = T36[1'h0:1'h0];
  assign T73 = T36[1'h1:1'h1];
  assign T74 = T36[2'h2:2'h2];
  assign io_out_bits_payload_a_type = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T78 = T36[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T80 = T36[1'h0:1'h0];
  assign T81 = T36[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_bits_payload_a_type : io_in_4_bits_payload_a_type;
  assign T84 = T36[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_bits_payload_a_type : io_in_6_bits_payload_a_type;
  assign T86 = T36[1'h0:1'h0];
  assign T87 = T36[1'h1:1'h1];
  assign T88 = T36[2'h2:2'h2];
  assign io_out_bits_payload_data = T89;
  assign T89 = T102 ? T96 : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T92 = T36[1'h0:1'h0];
  assign T93 = T94 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T94 = T36[1'h0:1'h0];
  assign T95 = T36[1'h1:1'h1];
  assign T96 = T101 ? T99 : T97;
  assign T97 = T98 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T98 = T36[1'h0:1'h0];
  assign T99 = T100 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T100 = T36[1'h0:1'h0];
  assign T101 = T36[1'h1:1'h1];
  assign T102 = T36[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T103;
  assign T103 = T116 ? T110 : T104;
  assign T104 = T109 ? T107 : T105;
  assign T105 = T106 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T106 = T36[1'h0:1'h0];
  assign T107 = T108 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T108 = T36[1'h0:1'h0];
  assign T109 = T36[1'h1:1'h1];
  assign T110 = T115 ? T113 : T111;
  assign T111 = T112 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T112 = T36[1'h0:1'h0];
  assign T113 = T114 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T114 = T36[1'h0:1'h0];
  assign T115 = T36[1'h1:1'h1];
  assign T116 = T36[2'h2:2'h2];
  assign io_out_bits_payload_addr = T117;
  assign T117 = T130 ? T124 : T118;
  assign T118 = T123 ? T121 : T119;
  assign T119 = T120 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T120 = T36[1'h0:1'h0];
  assign T121 = T122 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T122 = T36[1'h0:1'h0];
  assign T123 = T36[1'h1:1'h1];
  assign T124 = T129 ? T127 : T125;
  assign T125 = T126 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T126 = T36[1'h0:1'h0];
  assign T127 = T128 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T128 = T36[1'h0:1'h0];
  assign T129 = T36[1'h1:1'h1];
  assign T130 = T36[2'h2:2'h2];
  assign io_out_bits_header_dst = T131;
  assign T131 = T144 ? T138 : T132;
  assign T132 = T137 ? T135 : T133;
  assign T133 = T134 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T134 = T36[1'h0:1'h0];
  assign T135 = T136 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T136 = T36[1'h0:1'h0];
  assign T137 = T36[1'h1:1'h1];
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T140 = T36[1'h0:1'h0];
  assign T141 = T142 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T142 = T36[1'h0:1'h0];
  assign T143 = T36[1'h1:1'h1];
  assign T144 = T36[2'h2:2'h2];
  assign io_out_bits_header_src = T145;
  assign T145 = T158 ? T152 : T146;
  assign T146 = T151 ? T149 : T147;
  assign T147 = T148 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T148 = T36[1'h0:1'h0];
  assign T149 = T150 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T150 = T36[1'h0:1'h0];
  assign T151 = T36[1'h1:1'h1];
  assign T152 = T157 ? T155 : T153;
  assign T153 = T154 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T154 = T36[1'h0:1'h0];
  assign T155 = T156 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T156 = T36[1'h0:1'h0];
  assign T157 = T36[1'h1:1'h1];
  assign T158 = T36[2'h2:2'h2];
  assign io_out_valid = T159;
  assign T159 = T172 ? T166 : T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162 ? io_in_1_valid : io_in_0_valid;
  assign T162 = T36[1'h0:1'h0];
  assign T163 = T164 ? io_in_3_valid : io_in_2_valid;
  assign T164 = T36[1'h0:1'h0];
  assign T165 = T36[1'h1:1'h1];
  assign T166 = T171 ? T169 : T167;
  assign T167 = T168 ? io_in_5_valid : io_in_4_valid;
  assign T168 = T36[1'h0:1'h0];
  assign T169 = T170 ? io_in_7_valid : io_in_6_valid;
  assign T170 = T36[1'h0:1'h0];
  assign T171 = T36[1'h1:1'h1];
  assign T172 = T36[2'h2:2'h2];
  assign io_in_0_ready = T173;
  assign T173 = T174 & io_out_ready;
  assign T174 = T199 | T175;
  assign T175 = T176 ^ 1'h1;
  assign T176 = T179 | T177;
  assign T177 = io_in_7_valid & T178;
  assign T178 = R17 < 3'h7;
  assign T179 = T182 | T180;
  assign T180 = io_in_6_valid & T181;
  assign T181 = R17 < 3'h6;
  assign T182 = T185 | T183;
  assign T183 = io_in_5_valid & T184;
  assign T184 = R17 < 3'h5;
  assign T185 = T188 | T186;
  assign T186 = io_in_4_valid & T187;
  assign T187 = R17 < 3'h4;
  assign T188 = T191 | T189;
  assign T189 = io_in_3_valid & T190;
  assign T190 = R17 < 3'h3;
  assign T191 = T194 | T192;
  assign T192 = io_in_2_valid & T193;
  assign T193 = R17 < 3'h2;
  assign T194 = T197 | T195;
  assign T195 = io_in_1_valid & T196;
  assign T196 = R17 < 3'h1;
  assign T197 = io_in_0_valid & T198;
  assign T198 = R17 < 3'h0;
  assign T199 = R17 < 3'h0;
  assign io_in_1_ready = T200;
  assign T200 = T201 & io_out_ready;
  assign T201 = T211 | T202;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T204 | io_in_0_valid;
  assign T204 = T205 | T177;
  assign T205 = T206 | T180;
  assign T206 = T207 | T183;
  assign T207 = T208 | T186;
  assign T208 = T209 | T189;
  assign T209 = T210 | T192;
  assign T210 = T197 | T195;
  assign T211 = T213 & T212;
  assign T212 = R17 < 3'h1;
  assign T213 = T197 ^ 1'h1;
  assign io_in_2_ready = T214;
  assign T214 = T215 & io_out_ready;
  assign T215 = T226 | T216;
  assign T216 = T217 ^ 1'h1;
  assign T217 = T218 | io_in_1_valid;
  assign T218 = T219 | io_in_0_valid;
  assign T219 = T220 | T177;
  assign T220 = T221 | T180;
  assign T221 = T222 | T183;
  assign T222 = T223 | T186;
  assign T223 = T224 | T189;
  assign T224 = T225 | T192;
  assign T225 = T197 | T195;
  assign T226 = T228 & T227;
  assign T227 = R17 < 3'h2;
  assign T228 = T229 ^ 1'h1;
  assign T229 = T197 | T195;
  assign io_in_3_ready = T230;
  assign T230 = T231 & io_out_ready;
  assign T231 = T243 | T232;
  assign T232 = T233 ^ 1'h1;
  assign T233 = T234 | io_in_2_valid;
  assign T234 = T235 | io_in_1_valid;
  assign T235 = T236 | io_in_0_valid;
  assign T236 = T237 | T177;
  assign T237 = T238 | T180;
  assign T238 = T239 | T183;
  assign T239 = T240 | T186;
  assign T240 = T241 | T189;
  assign T241 = T242 | T192;
  assign T242 = T197 | T195;
  assign T243 = T245 & T244;
  assign T244 = R17 < 3'h3;
  assign T245 = T246 ^ 1'h1;
  assign T246 = T247 | T192;
  assign T247 = T197 | T195;
  assign io_in_4_ready = T248;
  assign T248 = T249 & io_out_ready;
  assign T249 = T262 | T250;
  assign T250 = T251 ^ 1'h1;
  assign T251 = T252 | io_in_3_valid;
  assign T252 = T253 | io_in_2_valid;
  assign T253 = T254 | io_in_1_valid;
  assign T254 = T255 | io_in_0_valid;
  assign T255 = T256 | T177;
  assign T256 = T257 | T180;
  assign T257 = T258 | T183;
  assign T258 = T259 | T186;
  assign T259 = T260 | T189;
  assign T260 = T261 | T192;
  assign T261 = T197 | T195;
  assign T262 = T264 & T263;
  assign T263 = R17 < 3'h4;
  assign T264 = T265 ^ 1'h1;
  assign T265 = T266 | T189;
  assign T266 = T267 | T192;
  assign T267 = T197 | T195;
  assign io_in_5_ready = T268;
  assign T268 = T269 & io_out_ready;
  assign T269 = T283 | T270;
  assign T270 = T271 ^ 1'h1;
  assign T271 = T272 | io_in_4_valid;
  assign T272 = T273 | io_in_3_valid;
  assign T273 = T274 | io_in_2_valid;
  assign T274 = T275 | io_in_1_valid;
  assign T275 = T276 | io_in_0_valid;
  assign T276 = T277 | T177;
  assign T277 = T278 | T180;
  assign T278 = T279 | T183;
  assign T279 = T280 | T186;
  assign T280 = T281 | T189;
  assign T281 = T282 | T192;
  assign T282 = T197 | T195;
  assign T283 = T285 & T284;
  assign T284 = R17 < 3'h5;
  assign T285 = T286 ^ 1'h1;
  assign T286 = T287 | T186;
  assign T287 = T288 | T189;
  assign T288 = T289 | T192;
  assign T289 = T197 | T195;
  assign io_in_6_ready = T290;
  assign T290 = T291 & io_out_ready;
  assign T291 = T306 | T292;
  assign T292 = T293 ^ 1'h1;
  assign T293 = T294 | io_in_5_valid;
  assign T294 = T295 | io_in_4_valid;
  assign T295 = T296 | io_in_3_valid;
  assign T296 = T297 | io_in_2_valid;
  assign T297 = T298 | io_in_1_valid;
  assign T298 = T299 | io_in_0_valid;
  assign T299 = T300 | T177;
  assign T300 = T301 | T180;
  assign T301 = T302 | T183;
  assign T302 = T303 | T186;
  assign T303 = T304 | T189;
  assign T304 = T305 | T192;
  assign T305 = T197 | T195;
  assign T306 = T308 & T307;
  assign T307 = R17 < 3'h6;
  assign T308 = T309 ^ 1'h1;
  assign T309 = T310 | T183;
  assign T310 = T311 | T186;
  assign T311 = T312 | T189;
  assign T312 = T313 | T192;
  assign T313 = T197 | T195;
  assign io_in_7_ready = T314;
  assign T314 = T315 & io_out_ready;
  assign T315 = T331 | T316;
  assign T316 = T317 ^ 1'h1;
  assign T317 = T318 | io_in_6_valid;
  assign T318 = T319 | io_in_5_valid;
  assign T319 = T320 | io_in_4_valid;
  assign T320 = T321 | io_in_3_valid;
  assign T321 = T322 | io_in_2_valid;
  assign T322 = T323 | io_in_1_valid;
  assign T323 = T324 | io_in_0_valid;
  assign T324 = T325 | T177;
  assign T325 = T326 | T180;
  assign T326 = T327 | T183;
  assign T327 = T328 | T186;
  assign T328 = T329 | T189;
  assign T329 = T330 | T192;
  assign T330 = T197 | T195;
  assign T331 = T333 & T332;
  assign T332 = R17 < 3'h7;
  assign T333 = T334 ^ 1'h1;
  assign T334 = T335 | T180;
  assign T335 = T336 | T183;
  assign T336 = T337 | T186;
  assign T337 = T338 | T189;
  assign T338 = T339 | T192;
  assign T339 = T197 | T195;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T19) begin
      R17 <= T0;
    end
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input  io_in_7_bits_payload_master_xact_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input  io_in_6_bits_payload_master_xact_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input  io_in_5_bits_payload_master_xact_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input  io_in_4_bits_payload_master_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input  io_in_3_bits_payload_master_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input  io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input  io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input  io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output io_out_bits_payload_master_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T256;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[2:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire T64;
  wire[1:0] T65;
  wire T66;
  wire T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire T70;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T30 ? 3'h1 : T2;
  assign T2 = T28 ? 3'h2 : T3;
  assign T3 = T26 ? 3'h3 : T4;
  assign T4 = T24 ? 3'h4 : T5;
  assign T5 = T22 ? 3'h5 : T6;
  assign T6 = T20 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T256 = reset ? 3'h0 : T18;
  assign T18 = T19 ? T0 : R17;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = io_in_6_valid & T21;
  assign T21 = R17 < 3'h6;
  assign T22 = io_in_5_valid & T23;
  assign T23 = R17 < 3'h5;
  assign T24 = io_in_4_valid & T25;
  assign T25 = R17 < 3'h4;
  assign T26 = io_in_3_valid & T27;
  assign T27 = R17 < 3'h3;
  assign T28 = io_in_2_valid & T29;
  assign T29 = R17 < 3'h2;
  assign T30 = io_in_1_valid & T31;
  assign T31 = R17 < 3'h1;
  assign io_out_bits_payload_master_xact_id = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = T0;
  assign T37 = T38 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T38 = T36[1'h0:1'h0];
  assign T39 = T36[1'h1:1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T42 = T36[1'h0:1'h0];
  assign T43 = T44 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign T46 = T36[2'h2:2'h2];
  assign io_out_bits_header_dst = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T50 = T36[1'h0:1'h0];
  assign T51 = T52 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T58 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T58 = T36[1'h0:1'h0];
  assign T59 = T36[1'h1:1'h1];
  assign T60 = T36[2'h2:2'h2];
  assign io_out_bits_header_src = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T66 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T66 = T36[1'h0:1'h0];
  assign T67 = T36[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T70 = T36[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T72 = T36[1'h0:1'h0];
  assign T73 = T36[1'h1:1'h1];
  assign T74 = T36[2'h2:2'h2];
  assign io_out_valid = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_valid : io_in_0_valid;
  assign T78 = T36[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_valid : io_in_2_valid;
  assign T80 = T36[1'h0:1'h0];
  assign T81 = T36[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_valid : io_in_4_valid;
  assign T84 = T36[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_valid : io_in_6_valid;
  assign T86 = T36[1'h0:1'h0];
  assign T87 = T36[1'h1:1'h1];
  assign T88 = T36[2'h2:2'h2];
  assign io_in_0_ready = T89;
  assign T89 = T90 & io_out_ready;
  assign T90 = T115 | T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T95 | T93;
  assign T93 = io_in_7_valid & T94;
  assign T94 = R17 < 3'h7;
  assign T95 = T98 | T96;
  assign T96 = io_in_6_valid & T97;
  assign T97 = R17 < 3'h6;
  assign T98 = T101 | T99;
  assign T99 = io_in_5_valid & T100;
  assign T100 = R17 < 3'h5;
  assign T101 = T104 | T102;
  assign T102 = io_in_4_valid & T103;
  assign T103 = R17 < 3'h4;
  assign T104 = T107 | T105;
  assign T105 = io_in_3_valid & T106;
  assign T106 = R17 < 3'h3;
  assign T107 = T110 | T108;
  assign T108 = io_in_2_valid & T109;
  assign T109 = R17 < 3'h2;
  assign T110 = T113 | T111;
  assign T111 = io_in_1_valid & T112;
  assign T112 = R17 < 3'h1;
  assign T113 = io_in_0_valid & T114;
  assign T114 = R17 < 3'h0;
  assign T115 = R17 < 3'h0;
  assign io_in_1_ready = T116;
  assign T116 = T117 & io_out_ready;
  assign T117 = T127 | T118;
  assign T118 = T119 ^ 1'h1;
  assign T119 = T120 | io_in_0_valid;
  assign T120 = T121 | T93;
  assign T121 = T122 | T96;
  assign T122 = T123 | T99;
  assign T123 = T124 | T102;
  assign T124 = T125 | T105;
  assign T125 = T126 | T108;
  assign T126 = T113 | T111;
  assign T127 = T129 & T128;
  assign T128 = R17 < 3'h1;
  assign T129 = T113 ^ 1'h1;
  assign io_in_2_ready = T130;
  assign T130 = T131 & io_out_ready;
  assign T131 = T142 | T132;
  assign T132 = T133 ^ 1'h1;
  assign T133 = T134 | io_in_1_valid;
  assign T134 = T135 | io_in_0_valid;
  assign T135 = T136 | T93;
  assign T136 = T137 | T96;
  assign T137 = T138 | T99;
  assign T138 = T139 | T102;
  assign T139 = T140 | T105;
  assign T140 = T141 | T108;
  assign T141 = T113 | T111;
  assign T142 = T144 & T143;
  assign T143 = R17 < 3'h2;
  assign T144 = T145 ^ 1'h1;
  assign T145 = T113 | T111;
  assign io_in_3_ready = T146;
  assign T146 = T147 & io_out_ready;
  assign T147 = T159 | T148;
  assign T148 = T149 ^ 1'h1;
  assign T149 = T150 | io_in_2_valid;
  assign T150 = T151 | io_in_1_valid;
  assign T151 = T152 | io_in_0_valid;
  assign T152 = T153 | T93;
  assign T153 = T154 | T96;
  assign T154 = T155 | T99;
  assign T155 = T156 | T102;
  assign T156 = T157 | T105;
  assign T157 = T158 | T108;
  assign T158 = T113 | T111;
  assign T159 = T161 & T160;
  assign T160 = R17 < 3'h3;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T163 | T108;
  assign T163 = T113 | T111;
  assign io_in_4_ready = T164;
  assign T164 = T165 & io_out_ready;
  assign T165 = T178 | T166;
  assign T166 = T167 ^ 1'h1;
  assign T167 = T168 | io_in_3_valid;
  assign T168 = T169 | io_in_2_valid;
  assign T169 = T170 | io_in_1_valid;
  assign T170 = T171 | io_in_0_valid;
  assign T171 = T172 | T93;
  assign T172 = T173 | T96;
  assign T173 = T174 | T99;
  assign T174 = T175 | T102;
  assign T175 = T176 | T105;
  assign T176 = T177 | T108;
  assign T177 = T113 | T111;
  assign T178 = T180 & T179;
  assign T179 = R17 < 3'h4;
  assign T180 = T181 ^ 1'h1;
  assign T181 = T182 | T105;
  assign T182 = T183 | T108;
  assign T183 = T113 | T111;
  assign io_in_5_ready = T184;
  assign T184 = T185 & io_out_ready;
  assign T185 = T199 | T186;
  assign T186 = T187 ^ 1'h1;
  assign T187 = T188 | io_in_4_valid;
  assign T188 = T189 | io_in_3_valid;
  assign T189 = T190 | io_in_2_valid;
  assign T190 = T191 | io_in_1_valid;
  assign T191 = T192 | io_in_0_valid;
  assign T192 = T193 | T93;
  assign T193 = T194 | T96;
  assign T194 = T195 | T99;
  assign T195 = T196 | T102;
  assign T196 = T197 | T105;
  assign T197 = T198 | T108;
  assign T198 = T113 | T111;
  assign T199 = T201 & T200;
  assign T200 = R17 < 3'h5;
  assign T201 = T202 ^ 1'h1;
  assign T202 = T203 | T102;
  assign T203 = T204 | T105;
  assign T204 = T205 | T108;
  assign T205 = T113 | T111;
  assign io_in_6_ready = T206;
  assign T206 = T207 & io_out_ready;
  assign T207 = T222 | T208;
  assign T208 = T209 ^ 1'h1;
  assign T209 = T210 | io_in_5_valid;
  assign T210 = T211 | io_in_4_valid;
  assign T211 = T212 | io_in_3_valid;
  assign T212 = T213 | io_in_2_valid;
  assign T213 = T214 | io_in_1_valid;
  assign T214 = T215 | io_in_0_valid;
  assign T215 = T216 | T93;
  assign T216 = T217 | T96;
  assign T217 = T218 | T99;
  assign T218 = T219 | T102;
  assign T219 = T220 | T105;
  assign T220 = T221 | T108;
  assign T221 = T113 | T111;
  assign T222 = T224 & T223;
  assign T223 = R17 < 3'h6;
  assign T224 = T225 ^ 1'h1;
  assign T225 = T226 | T99;
  assign T226 = T227 | T102;
  assign T227 = T228 | T105;
  assign T228 = T229 | T108;
  assign T229 = T113 | T111;
  assign io_in_7_ready = T230;
  assign T230 = T231 & io_out_ready;
  assign T231 = T247 | T232;
  assign T232 = T233 ^ 1'h1;
  assign T233 = T234 | io_in_6_valid;
  assign T234 = T235 | io_in_5_valid;
  assign T235 = T236 | io_in_4_valid;
  assign T236 = T237 | io_in_3_valid;
  assign T237 = T238 | io_in_2_valid;
  assign T238 = T239 | io_in_1_valid;
  assign T239 = T240 | io_in_0_valid;
  assign T240 = T241 | T93;
  assign T241 = T242 | T96;
  assign T242 = T243 | T99;
  assign T243 = T244 | T102;
  assign T244 = T245 | T105;
  assign T245 = T246 | T108;
  assign T246 = T113 | T111;
  assign T247 = T249 & T248;
  assign T248 = R17 < 3'h7;
  assign T249 = T250 ^ 1'h1;
  assign T250 = T251 | T96;
  assign T251 = T252 | T99;
  assign T252 = T253 | T102;
  assign T253 = T254 | T105;
  assign T254 = T255 | T108;
  assign T255 = T113 | T111;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T19) begin
      R17 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatPassesId(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [1:0] io_in_7_acquire_bits_header_src,
    input [1:0] io_in_7_acquire_bits_header_dst,
    input [25:0] io_in_7_acquire_bits_payload_addr,
    input [2:0] io_in_7_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_7_acquire_bits_payload_data,
    input [2:0] io_in_7_acquire_bits_payload_a_type,
    input [5:0] io_in_7_acquire_bits_payload_write_mask,
    input [2:0] io_in_7_acquire_bits_payload_subword_addr,
    input [3:0] io_in_7_acquire_bits_payload_atomic_opcode,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_header_src,
    output[1:0] io_in_7_grant_bits_header_dst,
    output[511:0] io_in_7_grant_bits_payload_data,
    output[2:0] io_in_7_grant_bits_payload_client_xact_id,
    output io_in_7_grant_bits_payload_master_xact_id,
    output[3:0] io_in_7_grant_bits_payload_g_type,
    output io_in_7_finish_ready,
    input  io_in_7_finish_valid,
    input [1:0] io_in_7_finish_bits_header_src,
    input [1:0] io_in_7_finish_bits_header_dst,
    input  io_in_7_finish_bits_payload_master_xact_id,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [1:0] io_in_6_acquire_bits_header_src,
    input [1:0] io_in_6_acquire_bits_header_dst,
    input [25:0] io_in_6_acquire_bits_payload_addr,
    input [2:0] io_in_6_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_6_acquire_bits_payload_data,
    input [2:0] io_in_6_acquire_bits_payload_a_type,
    input [5:0] io_in_6_acquire_bits_payload_write_mask,
    input [2:0] io_in_6_acquire_bits_payload_subword_addr,
    input [3:0] io_in_6_acquire_bits_payload_atomic_opcode,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_header_src,
    output[1:0] io_in_6_grant_bits_header_dst,
    output[511:0] io_in_6_grant_bits_payload_data,
    output[2:0] io_in_6_grant_bits_payload_client_xact_id,
    output io_in_6_grant_bits_payload_master_xact_id,
    output[3:0] io_in_6_grant_bits_payload_g_type,
    output io_in_6_finish_ready,
    input  io_in_6_finish_valid,
    input [1:0] io_in_6_finish_bits_header_src,
    input [1:0] io_in_6_finish_bits_header_dst,
    input  io_in_6_finish_bits_payload_master_xact_id,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [1:0] io_in_5_acquire_bits_header_src,
    input [1:0] io_in_5_acquire_bits_header_dst,
    input [25:0] io_in_5_acquire_bits_payload_addr,
    input [2:0] io_in_5_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_5_acquire_bits_payload_data,
    input [2:0] io_in_5_acquire_bits_payload_a_type,
    input [5:0] io_in_5_acquire_bits_payload_write_mask,
    input [2:0] io_in_5_acquire_bits_payload_subword_addr,
    input [3:0] io_in_5_acquire_bits_payload_atomic_opcode,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_header_src,
    output[1:0] io_in_5_grant_bits_header_dst,
    output[511:0] io_in_5_grant_bits_payload_data,
    output[2:0] io_in_5_grant_bits_payload_client_xact_id,
    output io_in_5_grant_bits_payload_master_xact_id,
    output[3:0] io_in_5_grant_bits_payload_g_type,
    output io_in_5_finish_ready,
    input  io_in_5_finish_valid,
    input [1:0] io_in_5_finish_bits_header_src,
    input [1:0] io_in_5_finish_bits_header_dst,
    input  io_in_5_finish_bits_payload_master_xact_id,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [1:0] io_in_4_acquire_bits_header_src,
    input [1:0] io_in_4_acquire_bits_header_dst,
    input [25:0] io_in_4_acquire_bits_payload_addr,
    input [2:0] io_in_4_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_4_acquire_bits_payload_data,
    input [2:0] io_in_4_acquire_bits_payload_a_type,
    input [5:0] io_in_4_acquire_bits_payload_write_mask,
    input [2:0] io_in_4_acquire_bits_payload_subword_addr,
    input [3:0] io_in_4_acquire_bits_payload_atomic_opcode,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_header_src,
    output[1:0] io_in_4_grant_bits_header_dst,
    output[511:0] io_in_4_grant_bits_payload_data,
    output[2:0] io_in_4_grant_bits_payload_client_xact_id,
    output io_in_4_grant_bits_payload_master_xact_id,
    output[3:0] io_in_4_grant_bits_payload_g_type,
    output io_in_4_finish_ready,
    input  io_in_4_finish_valid,
    input [1:0] io_in_4_finish_bits_header_src,
    input [1:0] io_in_4_finish_bits_header_dst,
    input  io_in_4_finish_bits_payload_master_xact_id,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [1:0] io_in_3_acquire_bits_header_src,
    input [1:0] io_in_3_acquire_bits_header_dst,
    input [25:0] io_in_3_acquire_bits_payload_addr,
    input [2:0] io_in_3_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_3_acquire_bits_payload_data,
    input [2:0] io_in_3_acquire_bits_payload_a_type,
    input [5:0] io_in_3_acquire_bits_payload_write_mask,
    input [2:0] io_in_3_acquire_bits_payload_subword_addr,
    input [3:0] io_in_3_acquire_bits_payload_atomic_opcode,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_header_src,
    output[1:0] io_in_3_grant_bits_header_dst,
    output[511:0] io_in_3_grant_bits_payload_data,
    output[2:0] io_in_3_grant_bits_payload_client_xact_id,
    output io_in_3_grant_bits_payload_master_xact_id,
    output[3:0] io_in_3_grant_bits_payload_g_type,
    output io_in_3_finish_ready,
    input  io_in_3_finish_valid,
    input [1:0] io_in_3_finish_bits_header_src,
    input [1:0] io_in_3_finish_bits_header_dst,
    input  io_in_3_finish_bits_payload_master_xact_id,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [2:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_2_acquire_bits_payload_data,
    input [2:0] io_in_2_acquire_bits_payload_a_type,
    input [5:0] io_in_2_acquire_bits_payload_write_mask,
    input [2:0] io_in_2_acquire_bits_payload_subword_addr,
    input [3:0] io_in_2_acquire_bits_payload_atomic_opcode,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[511:0] io_in_2_grant_bits_payload_data,
    output[2:0] io_in_2_grant_bits_payload_client_xact_id,
    output io_in_2_grant_bits_payload_master_xact_id,
    output[3:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input  io_in_2_finish_bits_payload_master_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [2:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[2:0] io_in_1_grant_bits_payload_client_xact_id,
    output io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input  io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [2:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[2:0] io_in_0_grant_bits_payload_client_xact_id,
    output io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input  io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[2:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [2:0] io_out_grant_bits_payload_client_xact_id,
    input  io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output io_out_finish_bits_payload_master_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire RRArbiter_2_io_in_7_ready;
  wire RRArbiter_2_io_in_6_ready;
  wire RRArbiter_2_io_in_5_ready;
  wire RRArbiter_2_io_in_4_ready;
  wire RRArbiter_2_io_in_3_ready;
  wire RRArbiter_2_io_in_2_ready;
  wire RRArbiter_2_io_in_1_ready;
  wire RRArbiter_2_io_in_0_ready;
  wire RRArbiter_2_io_out_valid;
  wire[1:0] RRArbiter_2_io_out_bits_header_src;
  wire[1:0] RRArbiter_2_io_out_bits_header_dst;
  wire[25:0] RRArbiter_2_io_out_bits_payload_addr;
  wire[2:0] RRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] RRArbiter_2_io_out_bits_payload_data;
  wire[2:0] RRArbiter_2_io_out_bits_payload_a_type;
  wire[5:0] RRArbiter_2_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_2_io_out_bits_payload_subword_addr;
  wire[3:0] RRArbiter_2_io_out_bits_payload_atomic_opcode;
  wire RRArbiter_3_io_in_7_ready;
  wire RRArbiter_3_io_in_6_ready;
  wire RRArbiter_3_io_in_5_ready;
  wire RRArbiter_3_io_in_4_ready;
  wire RRArbiter_3_io_in_3_ready;
  wire RRArbiter_3_io_in_2_ready;
  wire RRArbiter_3_io_in_1_ready;
  wire RRArbiter_3_io_in_0_ready;
  wire RRArbiter_3_io_out_valid;
  wire[1:0] RRArbiter_3_io_out_bits_header_src;
  wire[1:0] RRArbiter_3_io_out_bits_header_dst;
  wire RRArbiter_3_io_out_bits_payload_master_xact_id;


  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_3_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_3_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_3_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_3_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T15 ? io_in_7_grant_ready : T1;
  assign T1 = T14 ? io_in_6_grant_ready : T2;
  assign T2 = T13 ? io_in_5_grant_ready : T3;
  assign T3 = T12 ? io_in_4_grant_ready : T4;
  assign T4 = T11 ? io_in_3_grant_ready : T5;
  assign T5 = T10 ? io_in_2_grant_ready : T6;
  assign T6 = T9 ? io_in_1_grant_ready : T7;
  assign T7 = T8 ? io_in_0_grant_ready : 1'h0;
  assign T8 = io_out_grant_bits_payload_client_xact_id == 3'h0;
  assign T9 = io_out_grant_bits_payload_client_xact_id == 3'h1;
  assign T10 = io_out_grant_bits_payload_client_xact_id == 3'h2;
  assign T11 = io_out_grant_bits_payload_client_xact_id == 3'h3;
  assign T12 = io_out_grant_bits_payload_client_xact_id == 3'h4;
  assign T13 = io_out_grant_bits_payload_client_xact_id == 3'h5;
  assign T14 = io_out_grant_bits_payload_client_xact_id == 3'h6;
  assign T15 = io_out_grant_bits_payload_client_xact_id == 3'h7;
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_2_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_2_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_2_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_2_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_2_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_2_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_2_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_2_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_3_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T16;
  assign T16 = T8 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_2_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_3_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_2_io_in_1_ready;
  assign io_in_2_finish_ready = RRArbiter_3_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T18;
  assign T18 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = RRArbiter_2_io_in_2_ready;
  assign io_in_3_finish_ready = RRArbiter_3_io_in_3_ready;
  assign io_in_3_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_3_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_3_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_3_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_3_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_3_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_3_grant_valid = T19;
  assign T19 = T11 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = RRArbiter_2_io_in_3_ready;
  assign io_in_4_finish_ready = RRArbiter_3_io_in_4_ready;
  assign io_in_4_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_4_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_4_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_4_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_4_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_4_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_4_grant_valid = T20;
  assign T20 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = RRArbiter_2_io_in_4_ready;
  assign io_in_5_finish_ready = RRArbiter_3_io_in_5_ready;
  assign io_in_5_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_5_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_5_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_5_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_5_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_5_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_5_grant_valid = T21;
  assign T21 = T13 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = RRArbiter_2_io_in_5_ready;
  assign io_in_6_finish_ready = RRArbiter_3_io_in_6_ready;
  assign io_in_6_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_6_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_6_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_6_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_6_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_6_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_6_grant_valid = T22;
  assign T22 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = RRArbiter_2_io_in_6_ready;
  assign io_in_7_finish_ready = RRArbiter_3_io_in_7_ready;
  assign io_in_7_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_7_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_7_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_7_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_7_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_7_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_7_grant_valid = T23;
  assign T23 = T15 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = RRArbiter_2_io_in_7_ready;
  RRArbiter_3 RRArbiter_2(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_2_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_header_src( io_in_7_acquire_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_acquire_bits_header_dst ),
       .io_in_7_bits_payload_addr( io_in_7_acquire_bits_payload_addr ),
       .io_in_7_bits_payload_client_xact_id( io_in_7_acquire_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_data( io_in_7_acquire_bits_payload_data ),
       .io_in_7_bits_payload_a_type( io_in_7_acquire_bits_payload_a_type ),
       .io_in_7_bits_payload_write_mask( io_in_7_acquire_bits_payload_write_mask ),
       .io_in_7_bits_payload_subword_addr( io_in_7_acquire_bits_payload_subword_addr ),
       .io_in_7_bits_payload_atomic_opcode( io_in_7_acquire_bits_payload_atomic_opcode ),
       .io_in_6_ready( RRArbiter_2_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_header_src( io_in_6_acquire_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_acquire_bits_header_dst ),
       .io_in_6_bits_payload_addr( io_in_6_acquire_bits_payload_addr ),
       .io_in_6_bits_payload_client_xact_id( io_in_6_acquire_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_data( io_in_6_acquire_bits_payload_data ),
       .io_in_6_bits_payload_a_type( io_in_6_acquire_bits_payload_a_type ),
       .io_in_6_bits_payload_write_mask( io_in_6_acquire_bits_payload_write_mask ),
       .io_in_6_bits_payload_subword_addr( io_in_6_acquire_bits_payload_subword_addr ),
       .io_in_6_bits_payload_atomic_opcode( io_in_6_acquire_bits_payload_atomic_opcode ),
       .io_in_5_ready( RRArbiter_2_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_header_src( io_in_5_acquire_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_acquire_bits_header_dst ),
       .io_in_5_bits_payload_addr( io_in_5_acquire_bits_payload_addr ),
       .io_in_5_bits_payload_client_xact_id( io_in_5_acquire_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_data( io_in_5_acquire_bits_payload_data ),
       .io_in_5_bits_payload_a_type( io_in_5_acquire_bits_payload_a_type ),
       .io_in_5_bits_payload_write_mask( io_in_5_acquire_bits_payload_write_mask ),
       .io_in_5_bits_payload_subword_addr( io_in_5_acquire_bits_payload_subword_addr ),
       .io_in_5_bits_payload_atomic_opcode( io_in_5_acquire_bits_payload_atomic_opcode ),
       .io_in_4_ready( RRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_header_src( io_in_4_acquire_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_acquire_bits_header_dst ),
       .io_in_4_bits_payload_addr( io_in_4_acquire_bits_payload_addr ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_acquire_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_data( io_in_4_acquire_bits_payload_data ),
       .io_in_4_bits_payload_a_type( io_in_4_acquire_bits_payload_a_type ),
       .io_in_4_bits_payload_write_mask( io_in_4_acquire_bits_payload_write_mask ),
       .io_in_4_bits_payload_subword_addr( io_in_4_acquire_bits_payload_subword_addr ),
       .io_in_4_bits_payload_atomic_opcode( io_in_4_acquire_bits_payload_atomic_opcode ),
       .io_in_3_ready( RRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_header_src( io_in_3_acquire_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_acquire_bits_header_dst ),
       .io_in_3_bits_payload_addr( io_in_3_acquire_bits_payload_addr ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_acquire_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_data( io_in_3_acquire_bits_payload_data ),
       .io_in_3_bits_payload_a_type( io_in_3_acquire_bits_payload_a_type ),
       .io_in_3_bits_payload_write_mask( io_in_3_acquire_bits_payload_write_mask ),
       .io_in_3_bits_payload_subword_addr( io_in_3_acquire_bits_payload_subword_addr ),
       .io_in_3_bits_payload_atomic_opcode( io_in_3_acquire_bits_payload_atomic_opcode ),
       .io_in_2_ready( RRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_acquire_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_acquire_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_acquire_bits_payload_atomic_opcode ),
       .io_in_1_ready( RRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_2_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_2_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_2_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_4 RRArbiter_3(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_3_io_in_7_ready ),
       .io_in_7_valid( io_in_7_finish_valid ),
       .io_in_7_bits_header_src( io_in_7_finish_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_finish_bits_header_dst ),
       .io_in_7_bits_payload_master_xact_id( io_in_7_finish_bits_payload_master_xact_id ),
       .io_in_6_ready( RRArbiter_3_io_in_6_ready ),
       .io_in_6_valid( io_in_6_finish_valid ),
       .io_in_6_bits_header_src( io_in_6_finish_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_finish_bits_header_dst ),
       .io_in_6_bits_payload_master_xact_id( io_in_6_finish_bits_payload_master_xact_id ),
       .io_in_5_ready( RRArbiter_3_io_in_5_ready ),
       .io_in_5_valid( io_in_5_finish_valid ),
       .io_in_5_bits_header_src( io_in_5_finish_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_finish_bits_header_dst ),
       .io_in_5_bits_payload_master_xact_id( io_in_5_finish_bits_payload_master_xact_id ),
       .io_in_4_ready( RRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( io_in_4_finish_valid ),
       .io_in_4_bits_header_src( io_in_4_finish_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_finish_bits_header_dst ),
       .io_in_4_bits_payload_master_xact_id( io_in_4_finish_bits_payload_master_xact_id ),
       .io_in_3_ready( RRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( io_in_3_finish_valid ),
       .io_in_3_bits_header_src( io_in_3_finish_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_finish_bits_header_dst ),
       .io_in_3_bits_payload_master_xact_id( io_in_3_finish_bits_payload_master_xact_id ),
       .io_in_2_ready( RRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_finish_bits_payload_master_xact_id ),
       .io_in_1_ready( RRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_3_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module L2CoherenceAgent(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    output[1:0] io_outer_acquire_bits_header_dst,
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[2:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [2:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    output io_outer_finish_valid,
    output[1:0] io_outer_finish_bits_header_src,
    output[1:0] io_outer_finish_bits_header_dst,
    output io_outer_finish_bits_payload_master_xact_id,
    input  io_incoherent_1,
    input  io_incoherent_0
);

  wire T30;
  wire T31;
  wire any_acquire_conflict;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[2:0] release_idx;
  wire voluntary;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire VoluntaryReleaseTracker_io_inner_acquire_ready;
  wire VoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_src;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_dst;
  wire[511:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_data;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type;
  wire VoluntaryReleaseTracker_io_inner_probe_valid;
  wire VoluntaryReleaseTracker_io_inner_release_ready;
  wire VoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_header_src;
  wire[25:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type;
  wire[5:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode;
  wire VoluntaryReleaseTracker_io_outer_grant_ready;
  wire VoluntaryReleaseTracker_io_has_acquire_conflict;
  wire AcquireTracker_0_io_inner_acquire_ready;
  wire AcquireTracker_0_io_inner_grant_valid;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_0_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_0_io_inner_probe_valid;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_0_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_0_io_inner_release_ready;
  wire AcquireTracker_0_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_0_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_0_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_0_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_0_io_outer_grant_ready;
  wire AcquireTracker_0_io_has_acquire_conflict;
  wire AcquireTracker_1_io_inner_acquire_ready;
  wire AcquireTracker_1_io_inner_grant_valid;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_1_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_1_io_inner_probe_valid;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_1_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_1_io_inner_release_ready;
  wire AcquireTracker_1_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_1_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_1_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_1_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_1_io_outer_grant_ready;
  wire AcquireTracker_1_io_has_acquire_conflict;
  wire AcquireTracker_2_io_inner_acquire_ready;
  wire AcquireTracker_2_io_inner_grant_valid;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_2_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_2_io_inner_probe_valid;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_2_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_2_io_inner_release_ready;
  wire AcquireTracker_2_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_2_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_2_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_2_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_2_io_outer_grant_ready;
  wire AcquireTracker_2_io_has_acquire_conflict;
  wire AcquireTracker_3_io_inner_acquire_ready;
  wire AcquireTracker_3_io_inner_grant_valid;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_3_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_3_io_inner_probe_valid;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_3_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_3_io_inner_release_ready;
  wire AcquireTracker_3_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_3_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_3_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_3_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_3_io_outer_grant_ready;
  wire AcquireTracker_3_io_has_acquire_conflict;
  wire AcquireTracker_4_io_inner_acquire_ready;
  wire AcquireTracker_4_io_inner_grant_valid;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_4_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_4_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_4_io_inner_probe_valid;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_4_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_4_io_inner_release_ready;
  wire AcquireTracker_4_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_4_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_4_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_4_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_4_io_outer_grant_ready;
  wire AcquireTracker_4_io_has_acquire_conflict;
  wire AcquireTracker_5_io_inner_acquire_ready;
  wire AcquireTracker_5_io_inner_grant_valid;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_5_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_5_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_5_io_inner_probe_valid;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_5_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_5_io_inner_release_ready;
  wire AcquireTracker_5_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_5_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_5_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_5_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_5_io_outer_grant_ready;
  wire AcquireTracker_5_io_has_acquire_conflict;
  wire AcquireTracker_6_io_inner_acquire_ready;
  wire AcquireTracker_6_io_inner_grant_valid;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_6_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_6_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_6_io_inner_probe_valid;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_6_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_6_io_inner_release_ready;
  wire AcquireTracker_6_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_6_io_outer_acquire_bits_payload_addr;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_6_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_6_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_6_io_outer_grant_ready;
  wire AcquireTracker_6_io_has_acquire_conflict;
  wire alloc_arb_io_in_7_ready;
  wire alloc_arb_io_in_6_ready;
  wire alloc_arb_io_in_5_ready;
  wire alloc_arb_io_in_4_ready;
  wire alloc_arb_io_in_3_ready;
  wire alloc_arb_io_in_2_ready;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire probe_arb_io_in_7_ready;
  wire probe_arb_io_in_6_ready;
  wire probe_arb_io_in_5_ready;
  wire probe_arb_io_in_4_ready;
  wire probe_arb_io_in_3_ready;
  wire probe_arb_io_in_2_ready;
  wire probe_arb_io_in_1_ready;
  wire probe_arb_io_in_0_ready;
  wire probe_arb_io_out_valid;
  wire[1:0] probe_arb_io_out_bits_header_src;
  wire[1:0] probe_arb_io_out_bits_header_dst;
  wire[25:0] probe_arb_io_out_bits_payload_addr;
  wire[2:0] probe_arb_io_out_bits_payload_master_xact_id;
  wire[1:0] probe_arb_io_out_bits_payload_p_type;
  wire grant_arb_io_in_7_ready;
  wire grant_arb_io_in_6_ready;
  wire grant_arb_io_in_5_ready;
  wire grant_arb_io_in_4_ready;
  wire grant_arb_io_in_3_ready;
  wire grant_arb_io_in_2_ready;
  wire grant_arb_io_in_1_ready;
  wire grant_arb_io_in_0_ready;
  wire grant_arb_io_out_valid;
  wire[1:0] grant_arb_io_out_bits_header_src;
  wire[1:0] grant_arb_io_out_bits_header_dst;
  wire[511:0] grant_arb_io_out_bits_payload_data;
  wire[1:0] grant_arb_io_out_bits_payload_client_xact_id;
  wire[2:0] grant_arb_io_out_bits_payload_master_xact_id;
  wire[3:0] grant_arb_io_out_bits_payload_g_type;
  wire outer_arb_io_in_7_acquire_ready;
  wire outer_arb_io_in_7_grant_valid;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_7_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_7_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_7_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_7_grant_bits_payload_g_type;
  wire outer_arb_io_in_7_finish_ready;
  wire outer_arb_io_in_6_acquire_ready;
  wire outer_arb_io_in_6_grant_valid;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_6_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_6_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_6_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_6_grant_bits_payload_g_type;
  wire outer_arb_io_in_6_finish_ready;
  wire outer_arb_io_in_5_acquire_ready;
  wire outer_arb_io_in_5_grant_valid;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_5_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_5_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_5_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_5_grant_bits_payload_g_type;
  wire outer_arb_io_in_5_finish_ready;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_4_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_4_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_g_type;
  wire outer_arb_io_in_4_finish_ready;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_3_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_3_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_g_type;
  wire outer_arb_io_in_3_finish_ready;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_2_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_2_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_g_type;
  wire outer_arb_io_in_2_finish_ready;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_1_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_1_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_g_type;
  wire outer_arb_io_in_1_finish_ready;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_0_grant_bits_payload_data;
  wire[2:0] outer_arb_io_in_0_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_g_type;
  wire outer_arb_io_in_0_finish_ready;
  wire outer_arb_io_out_acquire_valid;
  wire[1:0] outer_arb_io_out_acquire_bits_header_src;
  wire[1:0] outer_arb_io_out_acquire_bits_header_dst;
  wire[25:0] outer_arb_io_out_acquire_bits_payload_addr;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_out_acquire_bits_payload_data;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_a_type;
  wire[5:0] outer_arb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_subword_addr;
  wire[3:0] outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  wire outer_arb_io_out_grant_ready;
  wire outer_arb_io_out_finish_valid;
  wire[1:0] outer_arb_io_out_finish_bits_header_src;
  wire[1:0] outer_arb_io_out_finish_bits_header_dst;
  wire outer_arb_io_out_finish_bits_payload_master_xact_id;


  assign T30 = io_inner_acquire_valid & T31;
  assign T31 = any_acquire_conflict ^ 1'h1;
  assign any_acquire_conflict = T17 | AcquireTracker_6_io_has_acquire_conflict;
  assign T17 = T18 | AcquireTracker_5_io_has_acquire_conflict;
  assign T18 = T19 | AcquireTracker_4_io_has_acquire_conflict;
  assign T19 = T20 | AcquireTracker_3_io_has_acquire_conflict;
  assign T20 = T21 | AcquireTracker_2_io_has_acquire_conflict;
  assign T21 = T22 | AcquireTracker_1_io_has_acquire_conflict;
  assign T22 = VoluntaryReleaseTracker_io_has_acquire_conflict | AcquireTracker_0_io_has_acquire_conflict;
  assign T32 = T33;
  assign T33 = {io_incoherent_1, io_incoherent_0};
  assign T34 = io_inner_release_valid & T35;
  assign T35 = release_idx == 3'h7;
  assign release_idx = voluntary ? 3'h0 : io_inner_release_bits_payload_master_xact_id;
  assign voluntary = io_inner_release_bits_payload_r_type == 3'h0;
  assign T36 = T33;
  assign T37 = io_inner_release_valid & T38;
  assign T38 = release_idx == 3'h6;
  assign T39 = T33;
  assign T40 = io_inner_release_valid & T41;
  assign T41 = release_idx == 3'h5;
  assign T42 = T33;
  assign T43 = io_inner_release_valid & T44;
  assign T44 = release_idx == 3'h4;
  assign T45 = T33;
  assign T46 = io_inner_release_valid & T47;
  assign T47 = release_idx == 3'h3;
  assign T48 = T33;
  assign T49 = io_inner_release_valid & T50;
  assign T50 = release_idx == 3'h2;
  assign T51 = T33;
  assign T52 = io_inner_release_valid & T53;
  assign T53 = release_idx == 3'h1;
  assign T54 = T33;
  assign T55 = io_inner_release_valid & T56;
  assign T56 = release_idx == 3'h0;
  assign io_outer_finish_bits_payload_master_xact_id = outer_arb_io_out_finish_bits_payload_master_xact_id;
  assign io_outer_finish_bits_header_dst = outer_arb_io_out_finish_bits_header_dst;
  assign io_outer_finish_bits_header_src = outer_arb_io_out_finish_bits_header_src;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_outer_acquire_bits_payload_subword_addr = outer_arb_io_out_acquire_bits_payload_subword_addr;
  assign io_outer_acquire_bits_payload_write_mask = outer_arb_io_out_acquire_bits_payload_write_mask;
  assign io_outer_acquire_bits_payload_a_type = outer_arb_io_out_acquire_bits_payload_a_type;
  assign io_outer_acquire_bits_payload_data = outer_arb_io_out_acquire_bits_payload_data;
  assign io_outer_acquire_bits_payload_client_xact_id = outer_arb_io_out_acquire_bits_payload_client_xact_id;
  assign io_outer_acquire_bits_payload_addr = outer_arb_io_out_acquire_bits_payload_addr;
  assign io_outer_acquire_bits_header_dst = outer_arb_io_out_acquire_bits_header_dst;
  assign io_outer_acquire_bits_header_src = outer_arb_io_out_acquire_bits_header_src;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T0;
  assign T0 = T14 ? T8 : T1;
  assign T1 = T7 ? T5 : T2;
  assign T2 = T3 ? AcquireTracker_0_io_inner_release_ready : VoluntaryReleaseTracker_io_inner_release_ready;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = release_idx;
  assign T5 = T6 ? AcquireTracker_2_io_inner_release_ready : AcquireTracker_1_io_inner_release_ready;
  assign T6 = T4[1'h0:1'h0];
  assign T7 = T4[1'h1:1'h1];
  assign T8 = T13 ? T11 : T9;
  assign T9 = T10 ? AcquireTracker_4_io_inner_release_ready : AcquireTracker_3_io_inner_release_ready;
  assign T10 = T4[1'h0:1'h0];
  assign T11 = T12 ? AcquireTracker_6_io_inner_release_ready : AcquireTracker_5_io_inner_release_ready;
  assign T12 = T4[1'h0:1'h0];
  assign T13 = T4[1'h1:1'h1];
  assign T14 = T4[2'h2:2'h2];
  assign io_inner_probe_bits_payload_p_type = probe_arb_io_out_bits_payload_p_type;
  assign io_inner_probe_bits_payload_master_xact_id = probe_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_probe_bits_payload_addr = probe_arb_io_out_bits_payload_addr;
  assign io_inner_probe_bits_header_dst = probe_arb_io_out_bits_header_dst;
  assign io_inner_probe_bits_header_src = probe_arb_io_out_bits_header_src;
  assign io_inner_probe_valid = probe_arb_io_out_valid;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_grant_bits_payload_g_type = grant_arb_io_out_bits_payload_g_type;
  assign io_inner_grant_bits_payload_master_xact_id = grant_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_grant_bits_payload_client_xact_id = grant_arb_io_out_bits_payload_client_xact_id;
  assign io_inner_grant_bits_payload_data = grant_arb_io_out_bits_payload_data;
  assign io_inner_grant_bits_header_dst = grant_arb_io_out_bits_header_dst;
  assign io_inner_grant_bits_header_src = grant_arb_io_out_bits_header_src;
  assign io_inner_grant_valid = grant_arb_io_out_valid;
  assign io_inner_acquire_ready = T15;
  assign T15 = T23 & T16;
  assign T16 = any_acquire_conflict ^ 1'h1;
  assign T23 = T24 | AcquireTracker_6_io_inner_acquire_ready;
  assign T24 = T25 | AcquireTracker_5_io_inner_acquire_ready;
  assign T25 = T26 | AcquireTracker_4_io_inner_acquire_ready;
  assign T26 = T27 | AcquireTracker_3_io_inner_acquire_ready;
  assign T27 = T28 | AcquireTracker_2_io_inner_acquire_ready;
  assign T28 = T29 | AcquireTracker_1_io_inner_acquire_ready;
  assign T29 = VoluntaryReleaseTracker_io_inner_acquire_ready | AcquireTracker_0_io_inner_acquire_ready;
  VoluntaryReleaseTracker VoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_0_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_0_ready ),
       .io_inner_grant_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_0_ready ),
       .io_inner_probe_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_header_src(  )
       //.io_inner_probe_bits_header_dst(  )
       //.io_inner_probe_bits_payload_addr(  )
       //.io_inner_probe_bits_payload_master_xact_id(  )
       //.io_inner_probe_bits_payload_p_type(  )
       .io_inner_release_ready( VoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T55 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T54 ),
       .io_has_acquire_conflict( VoluntaryReleaseTracker_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_0 AcquireTracker_0(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_0_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_1_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_1_ready ),
       .io_inner_grant_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_1_ready ),
       .io_inner_probe_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_0_io_inner_release_ready ),
       .io_inner_release_valid( T52 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T51 ),
       .io_has_acquire_conflict( AcquireTracker_0_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_1 AcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_2_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_2_ready ),
       .io_inner_grant_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_2_ready ),
       .io_inner_probe_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T49 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T48 ),
       .io_has_acquire_conflict( AcquireTracker_1_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_2 AcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_3_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_3_ready ),
       .io_inner_grant_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_3_ready ),
       .io_inner_probe_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T46 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T45 ),
       .io_has_acquire_conflict( AcquireTracker_2_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_3 AcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_4_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_4_ready ),
       .io_inner_grant_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_4_ready ),
       .io_inner_probe_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T43 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T42 ),
       .io_has_acquire_conflict( AcquireTracker_3_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_4 AcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_5_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_5_ready ),
       .io_inner_grant_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_5_ready ),
       .io_inner_probe_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( T40 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_4_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T39 ),
       .io_has_acquire_conflict( AcquireTracker_4_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_5 AcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_6_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_6_ready ),
       .io_inner_grant_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_6_ready ),
       .io_inner_probe_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( T37 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_5_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T36 ),
       .io_has_acquire_conflict( AcquireTracker_5_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_6 AcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_7_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_7_ready ),
       .io_inner_grant_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_7_ready ),
       .io_inner_probe_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( T34 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_6_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T32 ),
       .io_has_acquire_conflict( AcquireTracker_6_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  Arbiter_11 alloc_arb(
       .io_in_7_ready( alloc_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_acquire_ready ),
       //.io_in_7_bits(  )
       .io_in_6_ready( alloc_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_acquire_ready ),
       //.io_in_6_bits(  )
       .io_in_5_ready( alloc_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_acquire_ready ),
       //.io_in_5_bits(  )
       .io_in_4_ready( alloc_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_acquire_ready ),
       //.io_in_4_bits(  )
       .io_in_3_ready( alloc_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_acquire_ready ),
       //.io_in_3_bits(  )
       .io_in_2_ready( alloc_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_acquire_ready ),
       //.io_in_2_bits(  )
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_acquire_ready ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T30 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_7_bits = {1{$random}};
    assign alloc_arb.io_in_6_bits = {1{$random}};
    assign alloc_arb.io_in_5_bits = {1{$random}};
    assign alloc_arb.io_in_4_bits = {1{$random}};
    assign alloc_arb.io_in_3_bits = {1{$random}};
    assign alloc_arb.io_in_2_bits = {1{$random}};
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  Arbiter_12 probe_arb(
       .io_in_7_ready( probe_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_in_7_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_in_6_ready( probe_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_in_6_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_in_5_ready( probe_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_in_5_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_in_4_ready( probe_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_in_4_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_in_3_ready( probe_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_in_3_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_in_2_ready( probe_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_in_2_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_in_1_ready( probe_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_in_1_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_in_0_ready( probe_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_p_type(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( probe_arb_io_out_valid ),
       .io_out_bits_header_src( probe_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( probe_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( probe_arb_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( probe_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( probe_arb_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign probe_arb.io_in_0_bits_header_src = {1{$random}};
    assign probe_arb.io_in_0_bits_header_dst = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_addr = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_p_type = {1{$random}};
  `endif
  Arbiter_13 grant_arb(
       .io_in_7_ready( grant_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_in_7_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_in_7_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       .io_in_6_ready( grant_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_in_6_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_in_6_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       .io_in_5_ready( grant_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_in_5_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_in_5_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       .io_in_4_ready( grant_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_in_4_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_in_4_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       .io_in_3_ready( grant_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_in_3_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_in_3_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       .io_in_2_ready( grant_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_in_2_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       .io_in_1_ready( grant_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_in_1_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       .io_in_0_ready( grant_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_in_0_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_in_0_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( grant_arb_io_out_valid ),
       .io_out_bits_header_src( grant_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( grant_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_data( grant_arb_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( grant_arb_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( grant_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( grant_arb_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  UncachedTileLinkIOArbiterThatPassesId outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_in_7_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_in_7_acquire_bits_header_dst(  )
       .io_in_7_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_in_7_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_7_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_in_7_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_in_7_acquire_bits_payload_write_mask( AcquireTracker_6_io_outer_acquire_bits_payload_write_mask ),
       .io_in_7_acquire_bits_payload_subword_addr( AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_7_acquire_bits_payload_atomic_opcode( AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_7_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_in_7_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_in_7_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_in_7_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_in_7_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_in_7_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_in_7_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_in_7_finish_valid(  )
       //.io_in_7_finish_bits_header_src(  )
       //.io_in_7_finish_bits_header_dst(  )
       //.io_in_7_finish_bits_payload_master_xact_id(  )
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_in_6_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_in_6_acquire_bits_header_dst(  )
       .io_in_6_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_in_6_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_6_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_in_6_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_in_6_acquire_bits_payload_write_mask( AcquireTracker_5_io_outer_acquire_bits_payload_write_mask ),
       .io_in_6_acquire_bits_payload_subword_addr( AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_6_acquire_bits_payload_atomic_opcode( AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_6_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_in_6_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_in_6_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_in_6_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_in_6_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_in_6_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_in_6_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_in_6_finish_valid(  )
       //.io_in_6_finish_bits_header_src(  )
       //.io_in_6_finish_bits_header_dst(  )
       //.io_in_6_finish_bits_payload_master_xact_id(  )
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_in_5_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_in_5_acquire_bits_header_dst(  )
       .io_in_5_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_in_5_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_5_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_in_5_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_in_5_acquire_bits_payload_write_mask( AcquireTracker_4_io_outer_acquire_bits_payload_write_mask ),
       .io_in_5_acquire_bits_payload_subword_addr( AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_5_acquire_bits_payload_atomic_opcode( AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_5_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_in_5_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_in_5_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_in_5_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_in_5_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_in_5_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_in_5_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_in_5_finish_valid(  )
       //.io_in_5_finish_bits_header_src(  )
       //.io_in_5_finish_bits_header_dst(  )
       //.io_in_5_finish_bits_payload_master_xact_id(  )
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_in_4_acquire_bits_header_dst(  )
       .io_in_4_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_in_4_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_4_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_in_4_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_in_4_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_in_4_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_4_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_4_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_in_4_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_in_4_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_in_4_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_in_4_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_in_4_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_in_4_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_in_4_finish_valid(  )
       //.io_in_4_finish_bits_header_src(  )
       //.io_in_4_finish_bits_header_dst(  )
       //.io_in_4_finish_bits_payload_master_xact_id(  )
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_in_3_acquire_bits_header_dst(  )
       .io_in_3_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_in_3_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_3_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_in_3_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_in_3_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_in_3_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_3_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_3_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_in_3_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_in_3_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_in_3_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_in_3_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_in_3_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_in_3_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_in_3_finish_valid(  )
       //.io_in_3_finish_bits_header_src(  )
       //.io_in_3_finish_bits_header_dst(  )
       //.io_in_3_finish_bits_payload_master_xact_id(  )
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_in_2_acquire_bits_header_dst(  )
       .io_in_2_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_in_2_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_2_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_2_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_in_2_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_in_2_finish_valid(  )
       //.io_in_2_finish_bits_header_src(  )
       //.io_in_2_finish_bits_header_dst(  )
       //.io_in_2_finish_bits_payload_master_xact_id(  )
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_in_1_finish_valid(  )
       //.io_in_1_finish_bits_header_src(  )
       //.io_in_1_finish_bits_header_dst(  )
       //.io_in_1_finish_bits_payload_master_xact_id(  )
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_in_0_acquire_bits_header_dst(  )
       .io_in_0_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_in_0_finish_valid(  )
       //.io_in_0_finish_bits_header_src(  )
       //.io_in_0_finish_bits_header_dst(  )
       //.io_in_0_finish_bits_payload_master_xact_id(  )
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( outer_arb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( outer_arb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( outer_arb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( outer_arb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( outer_arb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( outer_arb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( outer_arb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( outer_arb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( outer_arb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_header_src( io_outer_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_outer_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_outer_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_outer_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_outer_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_outer_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_outer_finish_ready ),
       .io_out_finish_valid( outer_arb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( outer_arb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( outer_arb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( outer_arb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign outer_arb.io_in_7_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_valid = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_6_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_valid = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_5_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_valid = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_4_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_valid = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_valid = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_valid = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_valid = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_valid = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[5:0] T15;
  wire[4:0] T16;
  wire[25:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_rw = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_addr, T15};
  assign T15 = {io_enq_bits_tag, io_enq_bits_rw};
  assign io_deq_bits_tag = T16;
  assign T16 = T11[3'h5:1'h1];
  assign io_deq_bits_addr = T17;
  assign T17 = T11[5'h1f:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T16;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T17;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T18;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[127:0] T11;
  reg [127:0] ram [1:0];
  wire[127:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T16 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T17 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T18 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_data;
  end
endmodule

module MemIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [2:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input [2:0] io_uncached_acquire_bits_payload_a_type,
    input [5:0] io_uncached_acquire_bits_payload_write_mask,
    input [2:0] io_uncached_acquire_bits_payload_subword_addr,
    input [3:0] io_uncached_acquire_bits_payload_atomic_opcode,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[2:0] io_uncached_grant_bits_payload_client_xact_id,
    output io_uncached_grant_bits_payload_master_xact_id,
    output[3:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input  io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire[127:0] T56;
  reg [511:0] buf_out;
  wire[511:0] T57;
  wire[511:0] T58;
  wire T29;
  wire T30;
  reg  active_out;
  wire T53;
  wire T27;
  wire T28;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg [2:0] cnt_out;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T40;
  reg  has_data;
  wire T54;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg  cmd_sent_out;
  wire T55;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[511:0] T59;
  wire[383:0] T60;
  wire T38;
  wire T39;
  wire T61;
  wire T62;
  wire T63;
  wire[4:0] T64;
  reg [2:0] tag_out;
  wire[2:0] T65;
  reg [25:0] addr_out;
  wire[25:0] T66;
  wire T67;
  wire T68;
  wire T0;
  wire T1;
  reg [2:0] cnt_in;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  wire T5;
  reg  active_in;
  wire T51;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[3:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T52;
  reg [4:0] tag_in;
  wire[4:0] T17;
  wire[511:0] T18;
  reg [511:0] buf_in;
  wire[511:0] T19;
  wire[511:0] T20;
  wire[511:0] T21;
  wire[511:0] T22;
  wire[383:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire mem_cmd_q_io_enq_ready;
  wire mem_cmd_q_io_deq_valid;
  wire[25:0] mem_cmd_q_io_deq_bits_addr;
  wire[4:0] mem_cmd_q_io_deq_bits_tag;
  wire mem_cmd_q_io_deq_bits_rw;
  wire mem_data_q_io_enq_ready;
  wire mem_data_q_io_deq_valid;
  wire[127:0] mem_data_q_io_deq_bits_data;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    buf_out = {16{$random}};
    active_out = {1{$random}};
    cnt_out = {1{$random}};
    has_data = {1{$random}};
    cmd_sent_out = {1{$random}};
    tag_out = {1{$random}};
    addr_out = {1{$random}};
    cnt_in = {1{$random}};
    active_in = {1{$random}};
    tag_in = {1{$random}};
    buf_in = {16{$random}};
  end
`endif

  assign T56 = buf_out[7'h7f:1'h0];
  assign T57 = T38 ? T59 : T58;
  assign T58 = T29 ? io_uncached_acquire_bits_payload_data : buf_out;
  assign T29 = T30 & io_uncached_acquire_valid;
  assign T30 = active_out ^ 1'h1;
  assign T53 = reset ? 1'h0 : T27;
  assign T27 = T31 ? 1'h0 : T28;
  assign T28 = T29 ? 1'h1 : active_out;
  assign T31 = active_out & T32;
  assign T32 = cmd_sent_out & T33;
  assign T33 = T40 | T34;
  assign T34 = cnt_out == 3'h4;
  assign T35 = T38 ? T37 : T36;
  assign T36 = T29 ? 3'h0 : cnt_out;
  assign T37 = cnt_out + 3'h1;
  assign T40 = has_data ^ 1'h1;
  assign T54 = reset ? 1'h0 : T41;
  assign T41 = T29 ? T42 : has_data;
  assign T42 = T44 | T43;
  assign T43 = 3'h6 == io_uncached_acquire_bits_payload_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h5 == io_uncached_acquire_bits_payload_a_type;
  assign T46 = 3'h3 == io_uncached_acquire_bits_payload_a_type;
  assign T55 = reset ? 1'h0 : T47;
  assign T47 = T49 ? 1'h1 : T48;
  assign T48 = T29 ? 1'h0 : cmd_sent_out;
  assign T49 = active_out & T50;
  assign T50 = mem_cmd_q_io_enq_ready & T67;
  assign T59 = {128'h0, T60};
  assign T60 = buf_out >> 8'h80;
  assign T38 = active_out & T39;
  assign T39 = mem_data_q_io_enq_ready & T61;
  assign T61 = T63 & T62;
  assign T62 = cnt_out < 3'h4;
  assign T63 = active_out & has_data;
  assign T64 = {2'h0, tag_out};
  assign T65 = T29 ? io_uncached_acquire_bits_payload_client_xact_id : tag_out;
  assign T66 = T29 ? io_uncached_acquire_bits_payload_addr : addr_out;
  assign T67 = active_out & T68;
  assign T68 = cmd_sent_out ^ 1'h1;
  assign io_mem_resp_ready = T0;
  assign T0 = T13 | T1;
  assign T1 = cnt_in < 3'h4;
  assign T2 = T11 ? T10 : T3;
  assign T3 = T4 ? 3'h1 : cnt_in;
  assign T4 = T5 & io_mem_resp_valid;
  assign T5 = active_in ^ 1'h1;
  assign T51 = reset ? 1'h0 : T6;
  assign T6 = T8 ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : active_in;
  assign T8 = active_in & T9;
  assign T9 = io_uncached_grant_ready & io_uncached_grant_valid;
  assign T10 = cnt_in + 3'h1;
  assign T11 = active_in & T12;
  assign T12 = io_mem_resp_ready & io_mem_resp_valid;
  assign T13 = active_in ^ 1'h1;
  assign io_mem_req_data_bits_data = mem_data_q_io_deq_bits_data;
  assign io_mem_req_data_valid = mem_data_q_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = mem_cmd_q_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = mem_cmd_q_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = mem_cmd_q_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = mem_cmd_q_io_deq_valid;
  assign io_uncached_grant_bits_payload_g_type = T14;
  assign T14 = 4'h0;
  assign io_uncached_grant_bits_payload_master_xact_id = T15;
  assign T15 = 1'h0;
  assign io_uncached_grant_bits_payload_client_xact_id = T16;
  assign T16 = T52;
  assign T52 = tag_in[2'h2:1'h0];
  assign T17 = T4 ? io_mem_resp_bits_tag : tag_in;
  assign io_uncached_grant_bits_payload_data = T18;
  assign T18 = buf_in;
  assign T19 = T11 ? T22 : T20;
  assign T20 = T4 ? T21 : buf_in;
  assign T21 = io_mem_resp_bits_data << 9'h180;
  assign T22 = {io_mem_resp_bits_data, T23};
  assign T23 = buf_in[9'h1ff:8'h80];
  assign io_uncached_grant_valid = T24;
  assign T24 = active_in & T25;
  assign T25 = cnt_in == 3'h4;
  assign io_uncached_acquire_ready = T26;
  assign T26 = active_out ^ 1'h1;
  Queue_13 mem_cmd_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_cmd_q_io_enq_ready ),
       .io_enq_valid( T67 ),
       .io_enq_bits_addr( addr_out ),
       .io_enq_bits_tag( T64 ),
       .io_enq_bits_rw( has_data ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( mem_cmd_q_io_deq_valid ),
       .io_deq_bits_addr( mem_cmd_q_io_deq_bits_addr ),
       .io_deq_bits_tag( mem_cmd_q_io_deq_bits_tag ),
       .io_deq_bits_rw( mem_cmd_q_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_14 mem_data_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_data_q_io_enq_ready ),
       .io_enq_valid( T61 ),
       .io_enq_bits_data( T56 ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( mem_data_q_io_deq_valid ),
       .io_deq_bits_data( mem_data_q_io_deq_bits_data )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T38) begin
      buf_out <= T59;
    end else if(T29) begin
      buf_out <= io_uncached_acquire_bits_payload_data;
    end
    if(reset) begin
      active_out <= 1'h0;
    end else if(T31) begin
      active_out <= 1'h0;
    end else if(T29) begin
      active_out <= 1'h1;
    end
    if(T38) begin
      cnt_out <= T37;
    end else if(T29) begin
      cnt_out <= 3'h0;
    end
    if(reset) begin
      has_data <= 1'h0;
    end else if(T29) begin
      has_data <= T42;
    end
    if(reset) begin
      cmd_sent_out <= 1'h0;
    end else if(T49) begin
      cmd_sent_out <= 1'h1;
    end else if(T29) begin
      cmd_sent_out <= 1'h0;
    end
    if(T29) begin
      tag_out <= io_uncached_acquire_bits_payload_client_xact_id;
    end
    if(T29) begin
      addr_out <= io_uncached_acquire_bits_payload_addr;
    end
    if(T11) begin
      cnt_in <= T10;
    end else if(T4) begin
      cnt_in <= 3'h1;
    end
    if(reset) begin
      active_in <= 1'h0;
    end else if(T8) begin
      active_in <= 1'h0;
    end else if(T4) begin
      active_in <= 1'h1;
    end
    if(T4) begin
      tag_in <= io_mem_resp_bits_tag;
    end
    if(T11) begin
      buf_in <= T22;
    end else if(T4) begin
      buf_in <= T21;
    end
  end
endmodule

module HellaFlowQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[6:0] io_count
);

  wire[4:0] T0;
  wire[4:0] T1;
  wire[132:0] T2;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire atLeastTwo;
  wire T23;
  wire[5:0] T24;
  reg [5:0] deq_ptr;
  wire[5:0] T32;
  wire[5:0] T13;
  wire[5:0] T14;
  wire do_deq;
  wire T15;
  wire do_flow;
  wire T7;
  wire T16;
  reg [5:0] enq_ptr;
  wire[5:0] T33;
  wire[5:0] T9;
  wire[5:0] T10;
  wire do_enq;
  wire T6;
  wire T8;
  wire full;
  reg  maybe_full;
  wire T34;
  wire T25;
  wire T26;
  wire ptr_match;
  wire[5:0] T12;
  wire[5:0] T17;
  wire[132:0] T3;
  wire[132:0] T4;
  wire[132:0] T5;
  reg [5:0] ram_addr;
  wire[5:0] T11;
  wire empty;
  wire T27;
  wire[127:0] T28;
  wire[127:0] T29;
  wire T30;
  reg  ram_out_valid;
  wire T31;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    ram_addr = {1{$random}};
    ram_out_valid = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = empty ? io_enq_bits_tag : T1;
  assign T1 = T2[3'h4:1'h0];
  assign T18 = io_deq_ready & T19;
  assign T19 = atLeastTwo | T20;
  assign T20 = T22 & T21;
  assign T21 = empty ^ 1'h1;
  assign T22 = io_deq_valid ^ 1'h1;
  assign atLeastTwo = full | T23;
  assign T23 = 6'h2 <= T24;
  assign T24 = enq_ptr - deq_ptr;
  assign T32 = reset ? 6'h0 : T13;
  assign T13 = do_deq ? T14 : deq_ptr;
  assign T14 = deq_ptr + 6'h1;
  assign do_deq = T16 & T15;
  assign T15 = do_flow ^ 1'h1;
  assign do_flow = T7;
  assign T7 = empty & io_deq_ready;
  assign T16 = io_deq_ready & io_deq_valid;
  assign T33 = reset ? 6'h0 : T9;
  assign T9 = do_enq ? T10 : enq_ptr;
  assign T10 = enq_ptr + 6'h1;
  assign do_enq = T8 & T6;
  assign T6 = do_flow ^ 1'h1;
  assign T8 = io_enq_ready & io_enq_valid;
  assign full = ptr_match & maybe_full;
  assign T34 = reset ? 1'h0 : T25;
  assign T25 = T26 ? do_enq : maybe_full;
  assign T26 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = io_deq_valid ? T17 : deq_ptr;
  assign T17 = deq_ptr + 6'h1;
  HellaFlowQueue_ram ram (
    .CLK(clk),
    .W0A(enq_ptr),
    .W0E(do_enq),
    .W0I(T4),
    .R1A(T12),
    .R1E(T18),
    .R1O(T2)
  );
  assign T4 = T5;
  assign T5 = {io_enq_bits_data, io_enq_bits_tag};
  assign T11 = T18 ? T12 : ram_addr;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_deq_bits_data = T28;
  assign T28 = empty ? io_enq_bits_data : T29;
  assign T29 = T2[8'h84:3'h5];
  assign io_deq_valid = T30;
  assign T30 = empty ? io_enq_valid : ram_out_valid;
  assign io_enq_ready = T31;
  assign T31 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 6'h0;
    end else if(do_deq) begin
      deq_ptr <= T14;
    end
    if(reset) begin
      enq_ptr <= 6'h0;
    end else if(do_enq) begin
      enq_ptr <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T26) begin
      maybe_full <= do_enq;
    end
    if(T18) begin
      ram_addr <= T12;
    end
    ram_out_valid <= T18;
  end
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
);

  wire[4:0] T0;
  wire[132:0] T1;
  reg [132:0] ram [0:0];
  wire[132:0] T2;
  wire[132:0] T3;
  wire[132:0] T4;
  wire do_enq;
  wire[127:0] T5;
  wire T6;
  wire empty;
  reg  full;
  wire T11;
  wire T7;
  wire T8;
  wire do_deq;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {5{$random}};
    full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[3'h4:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {io_enq_bits_data, io_enq_bits_tag};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_data = T5;
  assign T5 = T1[8'h84:3'h5];
  assign io_deq_valid = T6;
  assign T6 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign T11 = reset ? 1'h0 : T7;
  assign T7 = T8 ? do_enq : full;
  assign T8 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T9;
  assign T9 = T10 | io_deq_ready;
  assign T10 = full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      full <= 1'h0;
    end else if(T8) begin
      full <= do_enq;
    end
  end
endmodule

module HellaQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[6:0] io_count
);

  wire fq_io_enq_ready;
  wire fq_io_deq_valid;
  wire[127:0] fq_io_deq_bits_data;
  wire[4:0] fq_io_deq_bits_tag;
  wire Queue_16_io_enq_ready;
  wire Queue_16_io_deq_valid;
  wire[127:0] Queue_16_io_deq_bits_data;
  wire[4:0] Queue_16_io_deq_bits_tag;


  assign io_deq_bits_tag = Queue_16_io_deq_bits_tag;
  assign io_deq_bits_data = Queue_16_io_deq_bits_data;
  assign io_deq_valid = Queue_16_io_deq_valid;
  assign io_enq_ready = fq_io_enq_ready;
  HellaFlowQueue fq(.clk(clk), .reset(reset),
       .io_enq_ready( fq_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_data( io_enq_bits_data ),
       .io_enq_bits_tag( io_enq_bits_tag ),
       .io_deq_ready( Queue_16_io_enq_ready ),
       .io_deq_valid( fq_io_deq_valid ),
       .io_deq_bits_data( fq_io_deq_bits_data ),
       .io_deq_bits_tag( fq_io_deq_bits_tag )
       //.io_count(  )
  );
  Queue_15 Queue_16(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_16_io_enq_ready ),
       .io_enq_valid( fq_io_deq_valid ),
       .io_enq_bits_data( fq_io_deq_bits_data ),
       .io_enq_bits_tag( fq_io_deq_bits_tag ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( Queue_16_io_deq_valid ),
       .io_deq_bits_data( Queue_16_io_deq_bits_data ),
       .io_deq_bits_tag( Queue_16_io_deq_bits_tag )
  );
endmodule

module MemPipeIOMemIOConverter(input clk, input reset,
    output io_cpu_req_cmd_ready,
    input  io_cpu_req_cmd_valid,
    input [25:0] io_cpu_req_cmd_bits_addr,
    input [4:0] io_cpu_req_cmd_bits_tag,
    input  io_cpu_req_cmd_bits_rw,
    output io_cpu_req_data_ready,
    input  io_cpu_req_data_valid,
    input [127:0] io_cpu_req_data_bits_data,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[127:0] io_cpu_resp_bits_data,
    output[4:0] io_cpu_resp_bits_tag,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire T0;
  wire cmdq_mask;
  wire watermark;
  reg [6:0] count;
  wire[6:0] T17;
  wire[6:0] T1;
  wire[6:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire T5;
  wire T6;
  wire dec;
  wire T7;
  wire T8;
  wire T9;
  wire inc;
  wire T10;
  wire[6:0] T11;
  wire T12;
  wire T13;
  wire[6:0] T14;
  wire T15;
  wire T16;
  wire resp_dataq_io_deq_valid;
  wire[127:0] resp_dataq_io_deq_bits_data;
  wire[4:0] resp_dataq_io_deq_bits_tag;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    count = {1{$random}};
  end
`endif

  assign io_mem_req_data_bits_data = io_cpu_req_data_bits_data;
  assign io_mem_req_data_valid = io_cpu_req_data_valid;
  assign io_mem_req_cmd_bits_rw = io_cpu_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = io_cpu_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = io_cpu_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = T0;
  assign T0 = io_cpu_req_cmd_valid & cmdq_mask;
  assign cmdq_mask = io_cpu_req_cmd_bits_rw | watermark;
  assign watermark = 7'h4 <= count;
  assign T17 = reset ? 7'h40 : T1;
  assign T1 = T15 ? T14 : T2;
  assign T2 = T12 ? T11 : T3;
  assign T3 = T5 ? T4 : count;
  assign T4 = count + 7'h1;
  assign T5 = inc & T6;
  assign T6 = dec ^ 1'h1;
  assign dec = T7;
  assign T7 = T9 & T8;
  assign T8 = io_mem_req_cmd_bits_rw ^ 1'h1;
  assign T9 = io_mem_req_cmd_ready & io_mem_req_cmd_valid;
  assign inc = T10;
  assign T10 = io_cpu_resp_ready & resp_dataq_io_deq_valid;
  assign T11 = count - 7'h4;
  assign T12 = T13 & dec;
  assign T13 = inc ^ 1'h1;
  assign T14 = count - 7'h3;
  assign T15 = inc & dec;
  assign io_cpu_resp_bits_tag = resp_dataq_io_deq_bits_tag;
  assign io_cpu_resp_bits_data = resp_dataq_io_deq_bits_data;
  assign io_cpu_resp_valid = resp_dataq_io_deq_valid;
  assign io_cpu_req_data_ready = io_mem_req_data_ready;
  assign io_cpu_req_cmd_ready = T16;
  assign T16 = io_mem_req_cmd_ready & cmdq_mask;
  HellaQueue resp_dataq(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_data( io_mem_resp_bits_data ),
       .io_enq_bits_tag( io_mem_resp_bits_tag ),
       .io_deq_ready( io_cpu_resp_ready ),
       .io_deq_valid( resp_dataq_io_deq_valid ),
       .io_deq_bits_data( resp_dataq_io_deq_bits_data ),
       .io_deq_bits_tag( resp_dataq_io_deq_bits_tag )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      count <= 7'h40;
    end else if(T15) begin
      count <= T14;
    end else if(T12) begin
      count <= T11;
    end else if(T5) begin
      count <= T4;
    end
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] ram [1:0];
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[5:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[4:0] T12;
  wire[25:0] T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_rw = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_addr, T5};
  assign T5 = {io_enq_bits_tag, io_enq_bits_rw};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_tag = T12;
  assign T12 = T1[3'h5:1'h1];
  assign io_deq_bits_addr = T13;
  assign T13 = T1[5'h1f:3'h6];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
);

  wire[127:0] T0;
  wire[127:0] T1;
  reg [127:0] ram [3:0];
  wire[127:0] T2;
  wire do_enq;
  reg [1:0] R3;
  wire[1:0] T14;
  wire[1:0] T4;
  wire[1:0] T5;
  reg [1:0] R6;
  wire[1:0] T15;
  wire[1:0] T7;
  wire[1:0] T8;
  wire do_deq;
  wire T9;
  wire empty;
  wire T10;
  reg  maybe_full;
  wire T16;
  wire T11;
  wire T12;
  wire ptr_match;
  wire T13;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {4{$random}};
    R3 = {1{$random}};
    R6 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[7'h7f:1'h0];
  assign T1 = ram[R6];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T14 = reset ? 2'h0 : T4;
  assign T4 = do_enq ? T5 : R3;
  assign T5 = R3 + 2'h1;
  assign T15 = reset ? 2'h0 : T7;
  assign T7 = do_deq ? T8 : R6;
  assign T8 = R6 + 2'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T9;
  assign T9 = empty ^ 1'h1;
  assign empty = ptr_match & T10;
  assign T10 = maybe_full ^ 1'h1;
  assign T16 = reset ? 1'h0 : T11;
  assign T11 = T12 ? do_enq : maybe_full;
  assign T12 = do_enq != do_deq;
  assign ptr_match = R3 == R6;
  assign io_enq_ready = T13;
  assign T13 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R3] <= io_enq_bits_data;
    if(reset) begin
      R3 <= 2'h0;
    end else if(do_enq) begin
      R3 <= T5;
    end
    if(reset) begin
      R6 <= 2'h0;
    end else if(do_deq) begin
      R6 <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T12) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module MemPipeIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [2:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input [2:0] io_uncached_acquire_bits_payload_a_type,
    input [5:0] io_uncached_acquire_bits_payload_write_mask,
    input [2:0] io_uncached_acquire_bits_payload_subword_addr,
    input [3:0] io_uncached_acquire_bits_payload_atomic_opcode,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[2:0] io_uncached_grant_bits_payload_client_xact_id,
    output io_uncached_grant_bits_payload_master_xact_id,
    output[3:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input  io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire Queue_14_io_enq_ready;
  wire Queue_14_io_deq_valid;
  wire[25:0] Queue_14_io_deq_bits_addr;
  wire[4:0] Queue_14_io_deq_bits_tag;
  wire Queue_14_io_deq_bits_rw;
  wire Queue_15_io_enq_ready;
  wire Queue_15_io_deq_valid;
  wire[127:0] Queue_15_io_deq_bits_data;
  wire a_io_uncached_acquire_ready;
  wire a_io_uncached_grant_valid;
  wire[511:0] a_io_uncached_grant_bits_payload_data;
  wire[2:0] a_io_uncached_grant_bits_payload_client_xact_id;
  wire a_io_uncached_grant_bits_payload_master_xact_id;
  wire[3:0] a_io_uncached_grant_bits_payload_g_type;
  wire a_io_mem_req_cmd_valid;
  wire[25:0] a_io_mem_req_cmd_bits_addr;
  wire[4:0] a_io_mem_req_cmd_bits_tag;
  wire a_io_mem_req_cmd_bits_rw;
  wire a_io_mem_req_data_valid;
  wire[127:0] a_io_mem_req_data_bits_data;
  wire a_io_mem_resp_ready;
  wire b_io_cpu_req_cmd_ready;
  wire b_io_cpu_req_data_ready;
  wire b_io_cpu_resp_valid;
  wire[127:0] b_io_cpu_resp_bits_data;
  wire[4:0] b_io_cpu_resp_bits_tag;
  wire b_io_mem_req_cmd_valid;
  wire[25:0] b_io_mem_req_cmd_bits_addr;
  wire[4:0] b_io_mem_req_cmd_bits_tag;
  wire b_io_mem_req_cmd_bits_rw;
  wire b_io_mem_req_data_valid;
  wire[127:0] b_io_mem_req_data_bits_data;


  assign io_mem_req_data_bits_data = b_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = b_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = b_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = b_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = b_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = b_io_mem_req_cmd_valid;
  assign io_uncached_grant_bits_payload_g_type = a_io_uncached_grant_bits_payload_g_type;
  assign io_uncached_grant_bits_payload_master_xact_id = a_io_uncached_grant_bits_payload_master_xact_id;
  assign io_uncached_grant_bits_payload_client_xact_id = a_io_uncached_grant_bits_payload_client_xact_id;
  assign io_uncached_grant_bits_payload_data = a_io_uncached_grant_bits_payload_data;
  assign io_uncached_grant_valid = a_io_uncached_grant_valid;
  assign io_uncached_acquire_ready = a_io_uncached_acquire_ready;
  MemIOUncachedTileLinkIOConverter a(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( a_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( io_uncached_acquire_valid ),
       .io_uncached_acquire_bits_header_src( io_uncached_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( io_uncached_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( io_uncached_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( io_uncached_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( io_uncached_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_a_type( io_uncached_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_write_mask( io_uncached_acquire_bits_payload_write_mask ),
       .io_uncached_acquire_bits_payload_subword_addr( io_uncached_acquire_bits_payload_subword_addr ),
       .io_uncached_acquire_bits_payload_atomic_opcode( io_uncached_acquire_bits_payload_atomic_opcode ),
       .io_uncached_grant_ready( io_uncached_grant_ready ),
       .io_uncached_grant_valid( a_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( a_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( a_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( a_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_g_type( a_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( io_uncached_finish_valid ),
       .io_uncached_finish_bits_header_src( io_uncached_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( io_uncached_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( io_uncached_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( Queue_14_io_enq_ready ),
       .io_mem_req_cmd_valid( a_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( a_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( a_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( a_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( Queue_15_io_enq_ready ),
       .io_mem_req_data_valid( a_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( a_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( a_io_mem_resp_ready ),
       .io_mem_resp_valid( b_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( b_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_tag( b_io_cpu_resp_bits_tag )
  );
  MemPipeIOMemIOConverter b(.clk(clk), .reset(reset),
       .io_cpu_req_cmd_ready( b_io_cpu_req_cmd_ready ),
       .io_cpu_req_cmd_valid( Queue_14_io_deq_valid ),
       .io_cpu_req_cmd_bits_addr( Queue_14_io_deq_bits_addr ),
       .io_cpu_req_cmd_bits_tag( Queue_14_io_deq_bits_tag ),
       .io_cpu_req_cmd_bits_rw( Queue_14_io_deq_bits_rw ),
       .io_cpu_req_data_ready( b_io_cpu_req_data_ready ),
       .io_cpu_req_data_valid( Queue_15_io_deq_valid ),
       .io_cpu_req_data_bits_data( Queue_15_io_deq_bits_data ),
       .io_cpu_resp_ready( a_io_mem_resp_ready ),
       .io_cpu_resp_valid( b_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( b_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_tag( b_io_cpu_resp_bits_tag ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( b_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( b_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( b_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( b_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( b_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( b_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
  Queue_10 Queue_14(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_14_io_enq_ready ),
       .io_enq_valid( a_io_mem_req_cmd_valid ),
       .io_enq_bits_addr( a_io_mem_req_cmd_bits_addr ),
       .io_enq_bits_tag( a_io_mem_req_cmd_bits_tag ),
       .io_enq_bits_rw( a_io_mem_req_cmd_bits_rw ),
       .io_deq_ready( b_io_cpu_req_cmd_ready ),
       .io_deq_valid( Queue_14_io_deq_valid ),
       .io_deq_bits_addr( Queue_14_io_deq_bits_addr ),
       .io_deq_bits_tag( Queue_14_io_deq_bits_tag ),
       .io_deq_bits_rw( Queue_14_io_deq_bits_rw )
  );
  Queue_11 Queue_15(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_15_io_enq_ready ),
       .io_enq_valid( a_io_mem_req_data_valid ),
       .io_enq_bits_data( a_io_mem_req_data_bits_data ),
       .io_deq_ready( b_io_cpu_req_data_ready ),
       .io_deq_valid( Queue_15_io_deq_valid ),
       .io_deq_bits_data( Queue_15_io_deq_bits_data )
  );
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[2:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [2:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_acquire_ready,
    input  io_htif_acquire_valid,
    input [1:0] io_htif_acquire_bits_header_src,
    input [1:0] io_htif_acquire_bits_header_dst,
    input [25:0] io_htif_acquire_bits_payload_addr,
    input [1:0] io_htif_acquire_bits_payload_client_xact_id,
    input [511:0] io_htif_acquire_bits_payload_data,
    input [2:0] io_htif_acquire_bits_payload_a_type,
    input [5:0] io_htif_acquire_bits_payload_write_mask,
    input [2:0] io_htif_acquire_bits_payload_subword_addr,
    input [3:0] io_htif_acquire_bits_payload_atomic_opcode,
    input  io_htif_grant_ready,
    output io_htif_grant_valid,
    output[1:0] io_htif_grant_bits_header_src,
    output[1:0] io_htif_grant_bits_header_dst,
    output[511:0] io_htif_grant_bits_payload_data,
    output[1:0] io_htif_grant_bits_payload_client_xact_id,
    output[2:0] io_htif_grant_bits_payload_master_xact_id,
    output[3:0] io_htif_grant_bits_payload_g_type,
    output io_htif_finish_ready,
    input  io_htif_finish_valid,
    input [1:0] io_htif_finish_bits_header_src,
    input [1:0] io_htif_finish_bits_header_dst,
    input [2:0] io_htif_finish_bits_payload_master_xact_id,
    input  io_htif_probe_ready,
    output io_htif_probe_valid,
    output[1:0] io_htif_probe_bits_header_src,
    output[1:0] io_htif_probe_bits_header_dst,
    output[25:0] io_htif_probe_bits_payload_addr,
    output[2:0] io_htif_probe_bits_payload_master_xact_id,
    output[1:0] io_htif_probe_bits_payload_p_type,
    output io_htif_release_ready,
    input  io_htif_release_valid,
    input [1:0] io_htif_release_bits_header_src,
    input [1:0] io_htif_release_bits_header_dst,
    input [25:0] io_htif_release_bits_payload_addr,
    input [1:0] io_htif_release_bits_payload_client_xact_id,
    input [2:0] io_htif_release_bits_payload_master_xact_id,
    input [511:0] io_htif_release_bits_payload_data,
    input [2:0] io_htif_release_bits_payload_r_type,
    input  io_incoherent_1,
    input  io_incoherent_0,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire net_io_clients_1_acquire_ready;
  wire net_io_clients_1_grant_valid;
  wire[1:0] net_io_clients_1_grant_bits_header_src;
  wire[1:0] net_io_clients_1_grant_bits_header_dst;
  wire[511:0] net_io_clients_1_grant_bits_payload_data;
  wire[1:0] net_io_clients_1_grant_bits_payload_client_xact_id;
  wire[2:0] net_io_clients_1_grant_bits_payload_master_xact_id;
  wire[3:0] net_io_clients_1_grant_bits_payload_g_type;
  wire net_io_clients_1_finish_ready;
  wire net_io_clients_1_probe_valid;
  wire[1:0] net_io_clients_1_probe_bits_header_src;
  wire[1:0] net_io_clients_1_probe_bits_header_dst;
  wire[25:0] net_io_clients_1_probe_bits_payload_addr;
  wire[2:0] net_io_clients_1_probe_bits_payload_master_xact_id;
  wire[1:0] net_io_clients_1_probe_bits_payload_p_type;
  wire net_io_clients_1_release_ready;
  wire net_io_clients_0_acquire_ready;
  wire net_io_clients_0_grant_valid;
  wire[1:0] net_io_clients_0_grant_bits_header_src;
  wire[1:0] net_io_clients_0_grant_bits_header_dst;
  wire[511:0] net_io_clients_0_grant_bits_payload_data;
  wire[1:0] net_io_clients_0_grant_bits_payload_client_xact_id;
  wire[2:0] net_io_clients_0_grant_bits_payload_master_xact_id;
  wire[3:0] net_io_clients_0_grant_bits_payload_g_type;
  wire net_io_clients_0_finish_ready;
  wire net_io_clients_0_probe_valid;
  wire[1:0] net_io_clients_0_probe_bits_header_src;
  wire[1:0] net_io_clients_0_probe_bits_header_dst;
  wire[25:0] net_io_clients_0_probe_bits_payload_addr;
  wire[2:0] net_io_clients_0_probe_bits_payload_master_xact_id;
  wire[1:0] net_io_clients_0_probe_bits_payload_p_type;
  wire net_io_clients_0_release_ready;
  wire net_io_masters_0_acquire_valid;
  wire[1:0] net_io_masters_0_acquire_bits_header_src;
  wire[1:0] net_io_masters_0_acquire_bits_header_dst;
  wire[25:0] net_io_masters_0_acquire_bits_payload_addr;
  wire[1:0] net_io_masters_0_acquire_bits_payload_client_xact_id;
  wire[511:0] net_io_masters_0_acquire_bits_payload_data;
  wire[2:0] net_io_masters_0_acquire_bits_payload_a_type;
  wire[5:0] net_io_masters_0_acquire_bits_payload_write_mask;
  wire[2:0] net_io_masters_0_acquire_bits_payload_subword_addr;
  wire[3:0] net_io_masters_0_acquire_bits_payload_atomic_opcode;
  wire net_io_masters_0_grant_ready;
  wire net_io_masters_0_finish_valid;
  wire[1:0] net_io_masters_0_finish_bits_header_src;
  wire[1:0] net_io_masters_0_finish_bits_header_dst;
  wire[2:0] net_io_masters_0_finish_bits_payload_master_xact_id;
  wire net_io_masters_0_probe_ready;
  wire net_io_masters_0_release_valid;
  wire[1:0] net_io_masters_0_release_bits_header_src;
  wire[1:0] net_io_masters_0_release_bits_header_dst;
  wire[25:0] net_io_masters_0_release_bits_payload_addr;
  wire[1:0] net_io_masters_0_release_bits_payload_client_xact_id;
  wire[2:0] net_io_masters_0_release_bits_payload_master_xact_id;
  wire[511:0] net_io_masters_0_release_bits_payload_data;
  wire[2:0] net_io_masters_0_release_bits_payload_r_type;
  wire L2CoherenceAgent_io_inner_acquire_ready;
  wire L2CoherenceAgent_io_inner_grant_valid;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_dst;
  wire[511:0] L2CoherenceAgent_io_inner_grant_bits_payload_data;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] L2CoherenceAgent_io_inner_grant_bits_payload_g_type;
  wire L2CoherenceAgent_io_inner_finish_ready;
  wire L2CoherenceAgent_io_inner_probe_valid;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_dst;
  wire[25:0] L2CoherenceAgent_io_inner_probe_bits_payload_addr;
  wire[2:0] L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_payload_p_type;
  wire L2CoherenceAgent_io_inner_release_ready;
  wire L2CoherenceAgent_io_outer_acquire_valid;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_dst;
  wire[25:0] L2CoherenceAgent_io_outer_acquire_bits_payload_addr;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] L2CoherenceAgent_io_outer_acquire_bits_payload_data;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_a_type;
  wire[5:0] L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode;
  wire L2CoherenceAgent_io_outer_grant_ready;
  wire L2CoherenceAgent_io_outer_finish_valid;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_dst;
  wire L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id;
  wire conv_io_uncached_acquire_ready;
  wire conv_io_uncached_grant_valid;
  wire[511:0] conv_io_uncached_grant_bits_payload_data;
  wire[2:0] conv_io_uncached_grant_bits_payload_client_xact_id;
  wire conv_io_uncached_grant_bits_payload_master_xact_id;
  wire[3:0] conv_io_uncached_grant_bits_payload_g_type;
  wire conv_io_mem_req_cmd_valid;
  wire[25:0] conv_io_mem_req_cmd_bits_addr;
  wire[4:0] conv_io_mem_req_cmd_bits_tag;
  wire conv_io_mem_req_cmd_bits_rw;
  wire conv_io_mem_req_data_valid;
  wire[127:0] conv_io_mem_req_data_bits_data;


  assign io_mem_req_data_bits_data = conv_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = conv_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = conv_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = conv_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = conv_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = conv_io_mem_req_cmd_valid;
  assign io_htif_release_ready = net_io_clients_1_release_ready;
  assign io_htif_probe_bits_payload_p_type = net_io_clients_1_probe_bits_payload_p_type;
  assign io_htif_probe_bits_payload_master_xact_id = net_io_clients_1_probe_bits_payload_master_xact_id;
  assign io_htif_probe_bits_payload_addr = net_io_clients_1_probe_bits_payload_addr;
  assign io_htif_probe_bits_header_dst = net_io_clients_1_probe_bits_header_dst;
  assign io_htif_probe_bits_header_src = net_io_clients_1_probe_bits_header_src;
  assign io_htif_probe_valid = net_io_clients_1_probe_valid;
  assign io_htif_finish_ready = net_io_clients_1_finish_ready;
  assign io_htif_grant_bits_payload_g_type = net_io_clients_1_grant_bits_payload_g_type;
  assign io_htif_grant_bits_payload_master_xact_id = net_io_clients_1_grant_bits_payload_master_xact_id;
  assign io_htif_grant_bits_payload_client_xact_id = net_io_clients_1_grant_bits_payload_client_xact_id;
  assign io_htif_grant_bits_payload_data = net_io_clients_1_grant_bits_payload_data;
  assign io_htif_grant_bits_header_dst = net_io_clients_1_grant_bits_header_dst;
  assign io_htif_grant_bits_header_src = net_io_clients_1_grant_bits_header_src;
  assign io_htif_grant_valid = net_io_clients_1_grant_valid;
  assign io_htif_acquire_ready = net_io_clients_1_acquire_ready;
  assign io_tiles_0_release_ready = net_io_clients_0_release_ready;
  assign io_tiles_0_probe_bits_payload_p_type = net_io_clients_0_probe_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = net_io_clients_0_probe_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = net_io_clients_0_probe_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = net_io_clients_0_probe_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = net_io_clients_0_probe_bits_header_src;
  assign io_tiles_0_probe_valid = net_io_clients_0_probe_valid;
  assign io_tiles_0_finish_ready = net_io_clients_0_finish_ready;
  assign io_tiles_0_grant_bits_payload_g_type = net_io_clients_0_grant_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = net_io_clients_0_grant_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = net_io_clients_0_grant_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = net_io_clients_0_grant_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = net_io_clients_0_grant_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = net_io_clients_0_grant_bits_header_src;
  assign io_tiles_0_grant_valid = net_io_clients_0_grant_valid;
  assign io_tiles_0_acquire_ready = net_io_clients_0_acquire_ready;
  RocketChipCrossbarNetwork net(.clk(clk), .reset(reset),
       .io_clients_1_acquire_ready( net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( io_htif_acquire_valid ),
       .io_clients_1_acquire_bits_header_src( io_htif_acquire_bits_header_src ),
       .io_clients_1_acquire_bits_header_dst( io_htif_acquire_bits_header_dst ),
       .io_clients_1_acquire_bits_payload_addr( io_htif_acquire_bits_payload_addr ),
       .io_clients_1_acquire_bits_payload_client_xact_id( io_htif_acquire_bits_payload_client_xact_id ),
       .io_clients_1_acquire_bits_payload_data( io_htif_acquire_bits_payload_data ),
       .io_clients_1_acquire_bits_payload_a_type( io_htif_acquire_bits_payload_a_type ),
       .io_clients_1_acquire_bits_payload_write_mask( io_htif_acquire_bits_payload_write_mask ),
       .io_clients_1_acquire_bits_payload_subword_addr( io_htif_acquire_bits_payload_subword_addr ),
       .io_clients_1_acquire_bits_payload_atomic_opcode( io_htif_acquire_bits_payload_atomic_opcode ),
       .io_clients_1_grant_ready( io_htif_grant_ready ),
       .io_clients_1_grant_valid( net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_header_src( net_io_clients_1_grant_bits_header_src ),
       .io_clients_1_grant_bits_header_dst( net_io_clients_1_grant_bits_header_dst ),
       .io_clients_1_grant_bits_payload_data( net_io_clients_1_grant_bits_payload_data ),
       .io_clients_1_grant_bits_payload_client_xact_id( net_io_clients_1_grant_bits_payload_client_xact_id ),
       .io_clients_1_grant_bits_payload_master_xact_id( net_io_clients_1_grant_bits_payload_master_xact_id ),
       .io_clients_1_grant_bits_payload_g_type( net_io_clients_1_grant_bits_payload_g_type ),
       .io_clients_1_finish_ready( net_io_clients_1_finish_ready ),
       .io_clients_1_finish_valid( io_htif_finish_valid ),
       .io_clients_1_finish_bits_header_src( io_htif_finish_bits_header_src ),
       .io_clients_1_finish_bits_header_dst( io_htif_finish_bits_header_dst ),
       .io_clients_1_finish_bits_payload_master_xact_id( io_htif_finish_bits_payload_master_xact_id ),
       .io_clients_1_probe_ready( io_htif_probe_ready ),
       .io_clients_1_probe_valid( net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_header_src( net_io_clients_1_probe_bits_header_src ),
       .io_clients_1_probe_bits_header_dst( net_io_clients_1_probe_bits_header_dst ),
       .io_clients_1_probe_bits_payload_addr( net_io_clients_1_probe_bits_payload_addr ),
       .io_clients_1_probe_bits_payload_master_xact_id( net_io_clients_1_probe_bits_payload_master_xact_id ),
       .io_clients_1_probe_bits_payload_p_type( net_io_clients_1_probe_bits_payload_p_type ),
       .io_clients_1_release_ready( net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( io_htif_release_valid ),
       .io_clients_1_release_bits_header_src( io_htif_release_bits_header_src ),
       .io_clients_1_release_bits_header_dst( io_htif_release_bits_header_dst ),
       .io_clients_1_release_bits_payload_addr( io_htif_release_bits_payload_addr ),
       .io_clients_1_release_bits_payload_client_xact_id( io_htif_release_bits_payload_client_xact_id ),
       .io_clients_1_release_bits_payload_master_xact_id( io_htif_release_bits_payload_master_xact_id ),
       .io_clients_1_release_bits_payload_data( io_htif_release_bits_payload_data ),
       .io_clients_1_release_bits_payload_r_type( io_htif_release_bits_payload_r_type ),
       .io_clients_0_acquire_ready( net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_0_acquire_valid ),
       .io_clients_0_acquire_bits_header_src( io_tiles_0_acquire_bits_header_src ),
       .io_clients_0_acquire_bits_header_dst( io_tiles_0_acquire_bits_header_dst ),
       .io_clients_0_acquire_bits_payload_addr( io_tiles_0_acquire_bits_payload_addr ),
       .io_clients_0_acquire_bits_payload_client_xact_id( io_tiles_0_acquire_bits_payload_client_xact_id ),
       .io_clients_0_acquire_bits_payload_data( io_tiles_0_acquire_bits_payload_data ),
       .io_clients_0_acquire_bits_payload_a_type( io_tiles_0_acquire_bits_payload_a_type ),
       .io_clients_0_acquire_bits_payload_write_mask( io_tiles_0_acquire_bits_payload_write_mask ),
       .io_clients_0_acquire_bits_payload_subword_addr( io_tiles_0_acquire_bits_payload_subword_addr ),
       .io_clients_0_acquire_bits_payload_atomic_opcode( io_tiles_0_acquire_bits_payload_atomic_opcode ),
       .io_clients_0_grant_ready( io_tiles_0_grant_ready ),
       .io_clients_0_grant_valid( net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_header_src( net_io_clients_0_grant_bits_header_src ),
       .io_clients_0_grant_bits_header_dst( net_io_clients_0_grant_bits_header_dst ),
       .io_clients_0_grant_bits_payload_data( net_io_clients_0_grant_bits_payload_data ),
       .io_clients_0_grant_bits_payload_client_xact_id( net_io_clients_0_grant_bits_payload_client_xact_id ),
       .io_clients_0_grant_bits_payload_master_xact_id( net_io_clients_0_grant_bits_payload_master_xact_id ),
       .io_clients_0_grant_bits_payload_g_type( net_io_clients_0_grant_bits_payload_g_type ),
       .io_clients_0_finish_ready( net_io_clients_0_finish_ready ),
       .io_clients_0_finish_valid( io_tiles_0_finish_valid ),
       .io_clients_0_finish_bits_header_src( io_tiles_0_finish_bits_header_src ),
       .io_clients_0_finish_bits_header_dst( io_tiles_0_finish_bits_header_dst ),
       .io_clients_0_finish_bits_payload_master_xact_id( io_tiles_0_finish_bits_payload_master_xact_id ),
       .io_clients_0_probe_ready( io_tiles_0_probe_ready ),
       .io_clients_0_probe_valid( net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_header_src( net_io_clients_0_probe_bits_header_src ),
       .io_clients_0_probe_bits_header_dst( net_io_clients_0_probe_bits_header_dst ),
       .io_clients_0_probe_bits_payload_addr( net_io_clients_0_probe_bits_payload_addr ),
       .io_clients_0_probe_bits_payload_master_xact_id( net_io_clients_0_probe_bits_payload_master_xact_id ),
       .io_clients_0_probe_bits_payload_p_type( net_io_clients_0_probe_bits_payload_p_type ),
       .io_clients_0_release_ready( net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_0_release_valid ),
       .io_clients_0_release_bits_header_src( io_tiles_0_release_bits_header_src ),
       .io_clients_0_release_bits_header_dst( io_tiles_0_release_bits_header_dst ),
       .io_clients_0_release_bits_payload_addr( io_tiles_0_release_bits_payload_addr ),
       .io_clients_0_release_bits_payload_client_xact_id( io_tiles_0_release_bits_payload_client_xact_id ),
       .io_clients_0_release_bits_payload_master_xact_id( io_tiles_0_release_bits_payload_master_xact_id ),
       .io_clients_0_release_bits_payload_data( io_tiles_0_release_bits_payload_data ),
       .io_clients_0_release_bits_payload_r_type( io_tiles_0_release_bits_payload_r_type ),
       .io_masters_0_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_masters_0_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_masters_0_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_masters_0_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_masters_0_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_masters_0_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_masters_0_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_masters_0_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_masters_0_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_masters_0_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_masters_0_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_masters_0_grant_ready( net_io_masters_0_grant_ready ),
       .io_masters_0_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_masters_0_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_masters_0_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_masters_0_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_masters_0_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_masters_0_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_masters_0_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_masters_0_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_masters_0_finish_valid( net_io_masters_0_finish_valid ),
       .io_masters_0_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_masters_0_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_masters_0_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_masters_0_probe_ready( net_io_masters_0_probe_ready ),
       .io_masters_0_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_masters_0_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_masters_0_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_masters_0_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_masters_0_probe_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id ),
       .io_masters_0_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_masters_0_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_masters_0_release_valid( net_io_masters_0_release_valid ),
       .io_masters_0_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_masters_0_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_masters_0_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_masters_0_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_masters_0_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_masters_0_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_masters_0_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type )
  );
  L2CoherenceAgent L2CoherenceAgent(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_inner_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_inner_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( net_io_masters_0_grant_ready ),
       .io_inner_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_inner_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_inner_finish_valid( net_io_masters_0_finish_valid ),
       .io_inner_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( net_io_masters_0_probe_ready ),
       .io_inner_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_inner_release_valid( net_io_masters_0_release_valid ),
       .io_inner_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_inner_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type ),
       .io_outer_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_outer_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_outer_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_outer_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_outer_grant_valid( conv_io_uncached_grant_valid ),
       //.io_outer_grant_bits_header_src(  )
       //.io_outer_grant_bits_header_dst(  )
       .io_outer_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_outer_finish_ready(  )
       .io_outer_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_outer_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_outer_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_outer_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_incoherent_1( io_incoherent_1 ),
       .io_incoherent_0( io_incoherent_0 )
  );
  `ifndef SYNTHESIS
    assign L2CoherenceAgent.io_outer_grant_bits_header_src = {1{$random}};
    assign L2CoherenceAgent.io_outer_grant_bits_header_dst = {1{$random}};
    assign L2CoherenceAgent.io_outer_finish_ready = {1{$random}};
  `endif
  MemPipeIOUncachedTileLinkIOConverter conv(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_uncached_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_write_mask( L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask ),
       .io_uncached_acquire_bits_payload_subword_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr ),
       .io_uncached_acquire_bits_payload_atomic_opcode( L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_uncached_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_uncached_grant_valid( conv_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_uncached_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( conv_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( conv_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( conv_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_a_type,
    input [5:0] io_enq_bits_payload_write_mask,
    input [2:0] io_enq_bits_payload_subword_addr,
    input [3:0] io_enq_bits_payload_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_a_type,
    output[5:0] io_deq_bits_payload_write_mask,
    output[2:0] io_deq_bits_payload_subword_addr,
    output[3:0] io_deq_bits_payload_atomic_opcode
);

  wire[3:0] T0;
  wire[559:0] T1;
  reg [559:0] ram [1:0];
  wire[559:0] T2;
  wire[559:0] T3;
  wire[559:0] T4;
  wire[527:0] T5;
  wire[12:0] T6;
  wire[6:0] T7;
  wire[514:0] T8;
  wire[31:0] T9;
  wire[27:0] T10;
  wire[3:0] T11;
  wire do_enq;
  reg  R12;
  wire T31;
  wire T13;
  wire T14;
  reg  R15;
  wire T32;
  wire T16;
  wire T17;
  wire do_deq;
  wire[2:0] T18;
  wire[5:0] T19;
  wire[2:0] T20;
  wire[511:0] T21;
  wire[1:0] T22;
  wire[25:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire empty;
  wire T27;
  reg  maybe_full;
  wire T33;
  wire T28;
  wire T29;
  wire ptr_match;
  wire T30;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R12 = {1{$random}};
    R15 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_atomic_opcode = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[R15];
  assign T3 = T4;
  assign T4 = {T9, T5};
  assign T5 = {T8, T6};
  assign T6 = {io_enq_bits_payload_write_mask, T7};
  assign T7 = {io_enq_bits_payload_subword_addr, io_enq_bits_payload_atomic_opcode};
  assign T8 = {io_enq_bits_payload_data, io_enq_bits_payload_a_type};
  assign T9 = {T11, T10};
  assign T10 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T11 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T31 = reset ? 1'h0 : T13;
  assign T13 = do_enq ? T14 : R12;
  assign T14 = R12 + 1'h1;
  assign T32 = reset ? 1'h0 : T16;
  assign T16 = do_deq ? T17 : R15;
  assign T17 = R15 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_subword_addr = T18;
  assign T18 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_write_mask = T19;
  assign T19 = T1[4'hc:3'h7];
  assign io_deq_bits_payload_a_type = T20;
  assign T20 = T1[4'hf:4'hd];
  assign io_deq_bits_payload_data = T21;
  assign T21 = T1[10'h20f:5'h10];
  assign io_deq_bits_payload_client_xact_id = T22;
  assign T22 = T1[10'h211:10'h210];
  assign io_deq_bits_payload_addr = T23;
  assign T23 = T1[10'h22b:10'h212];
  assign io_deq_bits_header_dst = T24;
  assign T24 = T1[10'h22d:10'h22c];
  assign io_deq_bits_header_src = T25;
  assign T25 = T1[10'h22f:10'h22e];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign T33 = reset ? 1'h0 : T28;
  assign T28 = T29 ? do_enq : maybe_full;
  assign T29 = do_enq != do_deq;
  assign ptr_match = R12 == R15;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R12] <= T3;
    if(reset) begin
      R12 <= 1'h0;
    end else if(do_enq) begin
      R12 <= T14;
    end
    if(reset) begin
      R15 <= 1'h0;
    end else if(do_deq) begin
      R15 <= T17;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T29) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type
);

  wire[2:0] T0;
  wire[549:0] T1;
  reg [549:0] ram [1:0];
  wire[549:0] T2;
  wire[549:0] T3;
  wire[549:0] T4;
  wire[519:0] T5;
  wire[514:0] T6;
  wire[4:0] T7;
  wire[29:0] T8;
  wire[27:0] T9;
  wire do_enq;
  reg  R10;
  wire T27;
  wire T11;
  wire T12;
  reg  R13;
  wire T28;
  wire T14;
  wire T15;
  wire do_deq;
  wire[511:0] T16;
  wire[2:0] T17;
  wire[1:0] T18;
  wire[25:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire empty;
  wire T23;
  reg  maybe_full;
  wire T29;
  wire T24;
  wire T25;
  wire ptr_match;
  wire T26;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R10 = {1{$random}};
    R13 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_r_type = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R13];
  assign T3 = T4;
  assign T4 = {T8, T5};
  assign T5 = {T7, T6};
  assign T6 = {io_enq_bits_payload_data, io_enq_bits_payload_r_type};
  assign T7 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_master_xact_id};
  assign T8 = {io_enq_bits_header_src, T9};
  assign T9 = {io_enq_bits_header_dst, io_enq_bits_payload_addr};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T27 = reset ? 1'h0 : T11;
  assign T11 = do_enq ? T12 : R10;
  assign T12 = R10 + 1'h1;
  assign T28 = reset ? 1'h0 : T14;
  assign T14 = do_deq ? T15 : R13;
  assign T15 = R13 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T16;
  assign T16 = T1[10'h202:2'h3];
  assign io_deq_bits_payload_master_xact_id = T17;
  assign T17 = T1[10'h205:10'h203];
  assign io_deq_bits_payload_client_xact_id = T18;
  assign T18 = T1[10'h207:10'h206];
  assign io_deq_bits_payload_addr = T19;
  assign T19 = T1[10'h221:10'h208];
  assign io_deq_bits_header_dst = T20;
  assign T20 = T1[10'h223:10'h222];
  assign io_deq_bits_header_src = T21;
  assign T21 = T1[10'h225:10'h224];
  assign io_deq_valid = T22;
  assign T22 = empty ^ 1'h1;
  assign empty = ptr_match & T23;
  assign T23 = maybe_full ^ 1'h1;
  assign T29 = reset ? 1'h0 : T24;
  assign T24 = T25 ? do_enq : maybe_full;
  assign T25 = do_enq != do_deq;
  assign ptr_match = R10 == R13;
  assign io_enq_ready = T26;
  assign T26 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R10] <= T3;
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_enq) begin
      R10 <= T12;
    end
    if(reset) begin
      R13 <= 1'h0;
    end else if(do_deq) begin
      R13 <= T15;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T25) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id
);

  wire[2:0] T0;
  wire[6:0] T1;
  reg [6:0] ram [1:0];
  wire[6:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire[4:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_master_xact_id = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_header_src, T5};
  assign T5 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_header_dst = T12;
  assign T12 = T1[3'h4:2'h3];
  assign io_deq_bits_header_src = T13;
  assign T13 = T1[3'h6:3'h5];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [511:0] io_enq_bits_payload_data,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [3:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[511:0] io_deq_bits_payload_data,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[3:0] io_deq_bits_payload_g_type
);

  wire[3:0] T0;
  wire[524:0] T1;
  reg [524:0] ram [0:0];
  wire[524:0] T2;
  wire[524:0] T3;
  wire[524:0] T4;
  wire[8:0] T5;
  wire[6:0] T6;
  wire[515:0] T7;
  wire[513:0] T8;
  wire do_enq;
  wire[2:0] T9;
  wire[1:0] T10;
  wire[511:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire empty;
  reg  full;
  wire T19;
  wire T15;
  wire T16;
  wire do_deq;
  wire T17;
  wire T18;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {17{$random}};
    full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_g_type = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_client_xact_id, T6};
  assign T6 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_g_type};
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_payload_master_xact_id = T9;
  assign T9 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_client_xact_id = T10;
  assign T10 = T1[4'h8:3'h7];
  assign io_deq_bits_payload_data = T11;
  assign T11 = T1[10'h208:4'h9];
  assign io_deq_bits_header_dst = T12;
  assign T12 = T1[10'h20a:10'h209];
  assign io_deq_bits_header_src = T13;
  assign T13 = T1[10'h20c:10'h20b];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign T19 = reset ? 1'h0 : T15;
  assign T15 = T16 ? do_enq : full;
  assign T16 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T17;
  assign T17 = T18 | io_deq_ready;
  assign T18 = full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      full <= 1'h0;
    end else if(T16) begin
      full <= do_enq;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[1:0] io_deq_bits_payload_p_type
);

  wire[1:0] T0;
  wire[34:0] T1;
  reg [34:0] ram [1:0];
  wire[34:0] T2;
  wire[34:0] T3;
  wire[34:0] T4;
  wire[30:0] T5;
  wire[4:0] T6;
  wire[3:0] T7;
  wire do_enq;
  reg  R8;
  wire T23;
  wire T9;
  wire T10;
  reg  R11;
  wire T24;
  wire T12;
  wire T13;
  wire do_deq;
  wire[2:0] T14;
  wire[25:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  reg  maybe_full;
  wire T25;
  wire T20;
  wire T21;
  wire ptr_match;
  wire T22;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R8 = {1{$random}};
    R11 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_p_type = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = ram[R11];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_addr, T6};
  assign T6 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_p_type};
  assign T7 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T23 = reset ? 1'h0 : T9;
  assign T9 = do_enq ? T10 : R8;
  assign T10 = R8 + 1'h1;
  assign T24 = reset ? 1'h0 : T12;
  assign T12 = do_deq ? T13 : R11;
  assign T13 = R11 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T14;
  assign T14 = T1[3'h4:2'h2];
  assign io_deq_bits_payload_addr = T15;
  assign T15 = T1[5'h1e:3'h5];
  assign io_deq_bits_header_dst = T16;
  assign T16 = T1[6'h20:5'h1f];
  assign io_deq_bits_header_src = T17;
  assign T17 = T1[6'h22:6'h21];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign T25 = reset ? 1'h0 : T20;
  assign T20 = T21 ? do_enq : maybe_full;
  assign T21 = do_enq != do_deq;
  assign ptr_match = R8 == R11;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R8] <= T3;
    if(reset) begin
      R8 <= 1'h0;
    end else if(do_enq) begin
      R8 <= T10;
    end
    if(reset) begin
      R11 <= 1'h0;
    end else if(do_deq) begin
      R11 <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T21) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[2:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [2:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[4:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr,
    input  io_incoherent_0
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire[2:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[511:0] T8;
  wire[2:0] T9;
  wire[1:0] T10;
  wire[25:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire[3:0] T15;
  wire[2:0] T16;
  wire[5:0] T17;
  wire[2:0] T18;
  wire[511:0] T19;
  wire[1:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire[2:0] T29;
  wire[511:0] T30;
  wire[2:0] T31;
  wire[1:0] T32;
  wire[25:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire T36;
  wire[3:0] T37;
  wire[2:0] T38;
  wire[5:0] T39;
  wire[2:0] T40;
  wire[511:0] T41;
  wire[1:0] T42;
  wire[25:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T0;
  wire T1;
  wire T2;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[25:0] Queue_4_io_deq_bits_payload_addr;
  wire[1:0] Queue_4_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_4_io_deq_bits_payload_data;
  wire[2:0] Queue_4_io_deq_bits_payload_a_type;
  wire[5:0] Queue_4_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_4_io_deq_bits_payload_subword_addr;
  wire[3:0] Queue_4_io_deq_bits_payload_atomic_opcode;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[1:0] Queue_5_io_deq_bits_header_src;
  wire[1:0] Queue_5_io_deq_bits_header_dst;
  wire[25:0] Queue_5_io_deq_bits_payload_addr;
  wire[1:0] Queue_5_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_5_io_deq_bits_payload_master_xact_id;
  wire[511:0] Queue_5_io_deq_bits_payload_data;
  wire[2:0] Queue_5_io_deq_bits_payload_r_type;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[1:0] Queue_6_io_deq_bits_header_src;
  wire[1:0] Queue_6_io_deq_bits_header_dst;
  wire[2:0] Queue_6_io_deq_bits_payload_master_xact_id;
  wire Queue_7_io_enq_ready;
  wire Queue_7_io_deq_valid;
  wire[1:0] Queue_7_io_deq_bits_header_src;
  wire[1:0] Queue_7_io_deq_bits_header_dst;
  wire[511:0] Queue_7_io_deq_bits_payload_data;
  wire[1:0] Queue_7_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_7_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_7_io_deq_bits_payload_g_type;
  wire Queue_8_io_enq_ready;
  wire Queue_8_io_deq_valid;
  wire[1:0] Queue_8_io_deq_bits_header_src;
  wire[1:0] Queue_8_io_deq_bits_header_dst;
  wire[25:0] Queue_8_io_deq_bits_payload_addr;
  wire[2:0] Queue_8_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_8_io_deq_bits_payload_p_type;
  wire Queue_9_io_enq_ready;
  wire Queue_9_io_deq_valid;
  wire[1:0] Queue_9_io_deq_bits_header_src;
  wire[1:0] Queue_9_io_deq_bits_header_dst;
  wire[25:0] Queue_9_io_deq_bits_payload_addr;
  wire[1:0] Queue_9_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_9_io_deq_bits_payload_data;
  wire[2:0] Queue_9_io_deq_bits_payload_a_type;
  wire[5:0] Queue_9_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_9_io_deq_bits_payload_subword_addr;
  wire[3:0] Queue_9_io_deq_bits_payload_atomic_opcode;
  wire Queue_10_io_enq_ready;
  wire Queue_10_io_deq_valid;
  wire[1:0] Queue_10_io_deq_bits_header_src;
  wire[1:0] Queue_10_io_deq_bits_header_dst;
  wire[25:0] Queue_10_io_deq_bits_payload_addr;
  wire[1:0] Queue_10_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_10_io_deq_bits_payload_master_xact_id;
  wire[511:0] Queue_10_io_deq_bits_payload_data;
  wire[2:0] Queue_10_io_deq_bits_payload_r_type;
  wire Queue_11_io_enq_ready;
  wire Queue_11_io_deq_valid;
  wire[1:0] Queue_11_io_deq_bits_header_src;
  wire[1:0] Queue_11_io_deq_bits_header_dst;
  wire[2:0] Queue_11_io_deq_bits_payload_master_xact_id;
  wire Queue_12_io_enq_ready;
  wire Queue_12_io_deq_valid;
  wire[1:0] Queue_12_io_deq_bits_header_src;
  wire[1:0] Queue_12_io_deq_bits_header_dst;
  wire[511:0] Queue_12_io_deq_bits_payload_data;
  wire[1:0] Queue_12_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_12_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_12_io_deq_bits_payload_g_type;
  wire Queue_13_io_enq_ready;
  wire Queue_13_io_deq_valid;
  wire[1:0] Queue_13_io_deq_bits_header_src;
  wire[1:0] Queue_13_io_deq_bits_header_dst;
  wire[25:0] Queue_13_io_deq_bits_payload_addr;
  wire[2:0] Queue_13_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_13_io_deq_bits_payload_p_type;
  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_pcr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire[4:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_payload_addr;
  wire[1:0] htif_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] htif_io_mem_acquire_bits_payload_data;
  wire[2:0] htif_io_mem_acquire_bits_payload_a_type;
  wire[5:0] htif_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] htif_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] htif_io_mem_acquire_bits_payload_atomic_opcode;
  wire htif_io_mem_grant_ready;
  wire htif_io_mem_finish_valid;
  wire[1:0] htif_io_mem_finish_bits_header_dst;
  wire[2:0] htif_io_mem_finish_bits_payload_master_xact_id;
  wire htif_io_mem_probe_ready;
  wire htif_io_mem_release_valid;
  wire[25:0] htif_io_mem_release_bits_payload_addr;
  wire[1:0] htif_io_mem_release_bits_payload_client_xact_id;
  wire[2:0] htif_io_mem_release_bits_payload_master_xact_id;
  wire[511:0] htif_io_mem_release_bits_payload_data;
  wire[2:0] htif_io_mem_release_bits_payload_r_type;
  wire outmemsys_io_tiles_0_acquire_ready;
  wire outmemsys_io_tiles_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_dst;
  wire[511:0] outmemsys_io_tiles_0_grant_bits_payload_data;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[2:0] outmemsys_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_g_type;
  wire outmemsys_io_tiles_0_finish_ready;
  wire outmemsys_io_tiles_0_probe_valid;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_dst;
  wire[25:0] outmemsys_io_tiles_0_probe_bits_payload_addr;
  wire[2:0] outmemsys_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_payload_p_type;
  wire outmemsys_io_tiles_0_release_ready;
  wire outmemsys_io_htif_acquire_ready;
  wire outmemsys_io_htif_grant_valid;
  wire[1:0] outmemsys_io_htif_grant_bits_header_src;
  wire[1:0] outmemsys_io_htif_grant_bits_header_dst;
  wire[511:0] outmemsys_io_htif_grant_bits_payload_data;
  wire[1:0] outmemsys_io_htif_grant_bits_payload_client_xact_id;
  wire[2:0] outmemsys_io_htif_grant_bits_payload_master_xact_id;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_g_type;
  wire outmemsys_io_htif_finish_ready;
  wire outmemsys_io_htif_probe_valid;
  wire[1:0] outmemsys_io_htif_probe_bits_header_src;
  wire[1:0] outmemsys_io_htif_probe_bits_header_dst;
  wire[25:0] outmemsys_io_htif_probe_bits_payload_addr;
  wire[2:0] outmemsys_io_htif_probe_bits_payload_master_xact_id;
  wire[1:0] outmemsys_io_htif_probe_bits_payload_p_type;
  wire outmemsys_io_htif_release_ready;
  wire outmemsys_io_mem_req_cmd_valid;
  wire[25:0] outmemsys_io_mem_req_cmd_bits_addr;
  wire[4:0] outmemsys_io_mem_req_cmd_bits_tag;
  wire outmemsys_io_mem_req_cmd_bits_rw;
  wire outmemsys_io_mem_req_data_valid;
  wire[127:0] outmemsys_io_mem_req_data_bits_data;


  assign T3 = htif_io_mem_finish_bits_payload_master_xact_id;
  assign T4 = htif_io_mem_finish_bits_header_dst;
  assign T5 = 2'h1;
  assign T6 = htif_io_mem_finish_valid;
  assign T7 = htif_io_mem_release_bits_payload_r_type;
  assign T8 = htif_io_mem_release_bits_payload_data;
  assign T9 = htif_io_mem_release_bits_payload_master_xact_id;
  assign T10 = htif_io_mem_release_bits_payload_client_xact_id;
  assign T11 = htif_io_mem_release_bits_payload_addr;
  assign T12 = 2'h0;
  assign T13 = 2'h1;
  assign T14 = htif_io_mem_release_valid;
  assign T15 = htif_io_mem_acquire_bits_payload_atomic_opcode;
  assign T16 = htif_io_mem_acquire_bits_payload_subword_addr;
  assign T17 = htif_io_mem_acquire_bits_payload_write_mask;
  assign T18 = htif_io_mem_acquire_bits_payload_a_type;
  assign T19 = htif_io_mem_acquire_bits_payload_data;
  assign T20 = htif_io_mem_acquire_bits_payload_client_xact_id;
  assign T21 = htif_io_mem_acquire_bits_payload_addr;
  assign T22 = 2'h0;
  assign T23 = 2'h1;
  assign T24 = htif_io_mem_acquire_valid;
  assign T25 = io_tiles_0_finish_bits_payload_master_xact_id;
  assign T26 = io_tiles_0_finish_bits_header_dst;
  assign T27 = 2'h0;
  assign T28 = io_tiles_0_finish_valid;
  assign T29 = io_tiles_0_release_bits_payload_r_type;
  assign T30 = io_tiles_0_release_bits_payload_data;
  assign T31 = io_tiles_0_release_bits_payload_master_xact_id;
  assign T32 = io_tiles_0_release_bits_payload_client_xact_id;
  assign T33 = io_tiles_0_release_bits_payload_addr;
  assign T34 = 2'h0;
  assign T35 = 2'h0;
  assign T36 = io_tiles_0_release_valid;
  assign T37 = io_tiles_0_acquire_bits_payload_atomic_opcode;
  assign T38 = io_tiles_0_acquire_bits_payload_subword_addr;
  assign T39 = io_tiles_0_acquire_bits_payload_write_mask;
  assign T40 = io_tiles_0_acquire_bits_payload_a_type;
  assign T41 = io_tiles_0_acquire_bits_payload_data;
  assign T42 = io_tiles_0_acquire_bits_payload_client_xact_id;
  assign T43 = io_tiles_0_acquire_bits_payload_addr;
  assign T44 = 2'h0;
  assign T45 = 2'h0;
  assign T46 = io_tiles_0_acquire_valid;
  assign T47 = Queue_10_io_enq_ready;
  assign T48 = Queue_11_io_enq_ready;
  assign T49 = Queue_9_io_enq_ready;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_tiles_0_release_ready = T0;
  assign T0 = Queue_5_io_enq_ready;
  assign io_tiles_0_probe_bits_payload_p_type = Queue_8_io_deq_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = Queue_8_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = Queue_8_io_deq_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = Queue_8_io_deq_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = Queue_8_io_deq_bits_header_src;
  assign io_tiles_0_probe_valid = Queue_8_io_deq_valid;
  assign io_tiles_0_finish_ready = T1;
  assign T1 = Queue_6_io_enq_ready;
  assign io_tiles_0_grant_bits_payload_g_type = Queue_7_io_deq_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = Queue_7_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = Queue_7_io_deq_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = Queue_7_io_deq_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = Queue_7_io_deq_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = Queue_7_io_deq_bits_header_src;
  assign io_tiles_0_grant_valid = Queue_7_io_deq_valid;
  assign io_tiles_0_acquire_ready = T2;
  assign T2 = Queue_4_io_enq_ready;
  assign io_mem_req_data_bits_data = outmemsys_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = outmemsys_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = outmemsys_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = outmemsys_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = outmemsys_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = outmemsys_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = htif_io_host_debug_stats_pcr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_pcr( htif_io_host_debug_stats_pcr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( T49 ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( htif_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( htif_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( htif_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( htif_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( htif_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( htif_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( htif_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( Queue_12_io_deq_valid ),
       .io_mem_grant_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_mem_grant_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_mem_grant_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( Queue_12_io_deq_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type ),
       .io_mem_finish_ready( T48 ),
       .io_mem_finish_valid( htif_io_mem_finish_valid ),
       //.io_mem_finish_bits_header_src(  )
       .io_mem_finish_bits_header_dst( htif_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( htif_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( htif_io_mem_probe_ready ),
       .io_mem_probe_valid( Queue_13_io_deq_valid ),
       .io_mem_probe_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_mem_probe_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( Queue_13_io_deq_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type ),
       .io_mem_release_ready( T47 ),
       .io_mem_release_valid( htif_io_mem_release_valid ),
       //.io_mem_release_bits_header_src(  )
       //.io_mem_release_bits_header_dst(  )
       .io_mem_release_bits_payload_addr( htif_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( htif_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( htif_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( htif_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( htif_io_mem_release_bits_payload_r_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
  `ifndef SYNTHESIS
    assign htif.io_mem_release_bits_payload_addr = {1{$random}};
    assign htif.io_mem_release_bits_payload_client_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_master_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_data = {16{$random}};
    assign htif.io_mem_release_bits_payload_r_type = {1{$random}};
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
  `endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_0_acquire_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Queue_4_io_deq_valid ),
       .io_tiles_0_acquire_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Queue_4_io_deq_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Queue_4_io_deq_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Queue_4_io_deq_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Queue_7_io_enq_ready ),
       .io_tiles_0_grant_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Queue_6_io_deq_valid ),
       .io_tiles_0_finish_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Queue_8_io_enq_ready ),
       .io_tiles_0_probe_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( outmemsys_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Queue_5_io_deq_valid ),
       .io_tiles_0_release_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Queue_5_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type ),
       .io_htif_acquire_ready( outmemsys_io_htif_acquire_ready ),
       .io_htif_acquire_valid( Queue_9_io_deq_valid ),
       .io_htif_acquire_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_htif_acquire_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_htif_acquire_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_htif_acquire_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_htif_acquire_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_htif_acquire_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_htif_acquire_bits_payload_write_mask( Queue_9_io_deq_bits_payload_write_mask ),
       .io_htif_acquire_bits_payload_subword_addr( Queue_9_io_deq_bits_payload_subword_addr ),
       .io_htif_acquire_bits_payload_atomic_opcode( Queue_9_io_deq_bits_payload_atomic_opcode ),
       .io_htif_grant_ready( Queue_12_io_enq_ready ),
       .io_htif_grant_valid( outmemsys_io_htif_grant_valid ),
       .io_htif_grant_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_htif_grant_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_htif_grant_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_htif_grant_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_htif_grant_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_htif_grant_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_htif_finish_ready( outmemsys_io_htif_finish_ready ),
       .io_htif_finish_valid( Queue_11_io_deq_valid ),
       .io_htif_finish_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_htif_finish_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_htif_finish_bits_payload_master_xact_id( Queue_11_io_deq_bits_payload_master_xact_id ),
       .io_htif_probe_ready( Queue_13_io_enq_ready ),
       .io_htif_probe_valid( outmemsys_io_htif_probe_valid ),
       .io_htif_probe_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_htif_probe_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_htif_probe_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_htif_probe_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_htif_probe_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_htif_release_ready( outmemsys_io_htif_release_ready ),
       .io_htif_release_valid( Queue_10_io_deq_valid ),
       .io_htif_release_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_htif_release_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_htif_release_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_htif_release_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_htif_release_bits_payload_master_xact_id( Queue_10_io_deq_bits_payload_master_xact_id ),
       .io_htif_release_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_htif_release_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type ),
       .io_incoherent_1( 1'h1 ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( outmemsys_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( outmemsys_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( outmemsys_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( outmemsys_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( outmemsys_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( outmemsys_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( T46 ),
       .io_enq_bits_header_src( T45 ),
       .io_enq_bits_header_dst( T44 ),
       .io_enq_bits_payload_addr( T43 ),
       .io_enq_bits_payload_client_xact_id( T42 ),
       .io_enq_bits_payload_data( T41 ),
       .io_enq_bits_payload_a_type( T40 ),
       .io_enq_bits_payload_write_mask( T39 ),
       .io_enq_bits_payload_subword_addr( T38 ),
       .io_enq_bits_payload_atomic_opcode( T37 ),
       .io_deq_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_4_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_4_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_4_io_deq_bits_payload_atomic_opcode )
  );
  Queue_4 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( T36 ),
       .io_enq_bits_header_src( T35 ),
       .io_enq_bits_header_dst( T34 ),
       .io_enq_bits_payload_addr( T33 ),
       .io_enq_bits_payload_client_xact_id( T32 ),
       .io_enq_bits_payload_master_xact_id( T31 ),
       .io_enq_bits_payload_data( T30 ),
       .io_enq_bits_payload_r_type( T29 ),
       .io_deq_ready( outmemsys_io_tiles_0_release_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_5_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type )
  );
  Queue_5 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( T28 ),
       .io_enq_bits_header_src( T27 ),
       .io_enq_bits_header_dst( T26 ),
       .io_enq_bits_payload_master_xact_id( T25 ),
       .io_deq_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id )
  );
  Queue_6 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_deq_ready( io_tiles_0_grant_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_7_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_7_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_7_io_deq_bits_payload_g_type )
  );
  Queue_7 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_deq_ready( io_tiles_0_probe_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_8_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_8_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_8_io_deq_bits_payload_p_type )
  );
  Queue_3 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( T24 ),
       .io_enq_bits_header_src( T23 ),
       .io_enq_bits_header_dst( T22 ),
       .io_enq_bits_payload_addr( T21 ),
       .io_enq_bits_payload_client_xact_id( T20 ),
       .io_enq_bits_payload_data( T19 ),
       .io_enq_bits_payload_a_type( T18 ),
       .io_enq_bits_payload_write_mask( T17 ),
       .io_enq_bits_payload_subword_addr( T16 ),
       .io_enq_bits_payload_atomic_opcode( T15 ),
       .io_deq_ready( outmemsys_io_htif_acquire_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_9_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_9_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_9_io_deq_bits_payload_atomic_opcode )
  );
  Queue_4 Queue_10(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_10_io_enq_ready ),
       .io_enq_valid( T14 ),
       .io_enq_bits_header_src( T13 ),
       .io_enq_bits_header_dst( T12 ),
       .io_enq_bits_payload_addr( T11 ),
       .io_enq_bits_payload_client_xact_id( T10 ),
       .io_enq_bits_payload_master_xact_id( T9 ),
       .io_enq_bits_payload_data( T8 ),
       .io_enq_bits_payload_r_type( T7 ),
       .io_deq_ready( outmemsys_io_htif_release_ready ),
       .io_deq_valid( Queue_10_io_deq_valid ),
       .io_deq_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_10_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type )
  );
  Queue_5 Queue_11(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_11_io_enq_ready ),
       .io_enq_valid( T6 ),
       .io_enq_bits_header_src( T5 ),
       .io_enq_bits_header_dst( T4 ),
       .io_enq_bits_payload_master_xact_id( T3 ),
       .io_deq_ready( outmemsys_io_htif_finish_ready ),
       .io_deq_valid( Queue_11_io_deq_valid ),
       .io_deq_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_11_io_deq_bits_payload_master_xact_id )
  );
  Queue_6 Queue_12(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_12_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_deq_ready( htif_io_mem_grant_ready ),
       .io_deq_valid( Queue_12_io_deq_valid ),
       .io_deq_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_12_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type )
  );
  Queue_7 Queue_13(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_13_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_deq_ready( htif_io_mem_probe_ready ),
       .io_deq_valid( Queue_13_io_deq_valid ),
       .io_deq_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_13_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type )
  );
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [4:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[4:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data
);

  wire[63:0] T0;
  wire[69:0] T1;
  reg [69:0] ram [1:0];
  wire[69:0] T2;
  wire[69:0] T3;
  wire[69:0] T4;
  wire[68:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[4:0] T12;
  wire T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_rw, T5};
  assign T5 = {io_enq_bits_addr, io_enq_bits_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_addr = T12;
  assign T12 = T1[7'h44:7'h40];
  assign io_deq_bits_rw = T13;
  assign T13 = T1[7'h45:7'h45];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits
);

  wire[63:0] T0;
  reg [63:0] ram [1:0];
  wire[63:0] T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits
);

  wire T0;
  reg [0:0] ram [1:0];
  wire T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    input  io_mem_backup_en,
    output io_in_mem_ready,
    input  io_in_mem_valid,
    input  io_out_mem_ready,
    output io_out_mem_valid,
    input [7:0] io_temac_rx_axis_fifo_tdata,
    input  io_temac_rx_axis_fifo_tvalid,
    output io_temac_rx_axis_fifo_tready,
    input  io_temac_rx_axis_fifo_tlast,
    output[7:0] io_temac_tx_axis_fifo_tdata,
    output io_temac_tx_axis_fifo_tvalid,
    input  io_temac_tx_axis_fifo_tready,
    output io_temac_tx_axis_fifo_tlast,
    output[11:0] io_temac_s_axi_awaddr,
    output io_temac_s_axi_awvalid,
    input  io_temac_s_axi_awready,
    output[31:0] io_temac_s_axi_wdata,
    output io_temac_s_axi_wvalid,
    input  io_temac_s_axi_wready,
    input [1:0] io_temac_s_axi_bresp,
    input  io_temac_s_axi_bvalid,
    output io_temac_s_axi_bready,
    output[11:0] io_temac_s_axi_araddr,
    output io_temac_s_axi_arvalid,
    input  io_temac_s_axi_arready,
    input [31:0] io_temac_s_axi_rdata,
    input [1:0] io_temac_s_axi_rresp,
    input  io_temac_s_axi_rvalid,
    output io_temac_s_axi_rready
);

  wire resetSigs_0;
  reg  R0;
  reg  R1;
  wire Queue_0_io_enq_ready;
  wire Queue_0_io_deq_valid;
  wire Queue_0_io_deq_bits_rw;
  wire[4:0] Queue_0_io_deq_bits_addr;
  wire[63:0] Queue_0_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire Queue_2_io_deq_bits;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire Queue_3_io_deq_bits;
  wire RocketTile_io_tilelink_acquire_valid;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_header_src;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_header_dst;
  wire[25:0] RocketTile_io_tilelink_acquire_bits_payload_addr;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_payload_client_xact_id;
  wire[511:0] RocketTile_io_tilelink_acquire_bits_payload_data;
  wire[2:0] RocketTile_io_tilelink_acquire_bits_payload_a_type;
  wire[5:0] RocketTile_io_tilelink_acquire_bits_payload_write_mask;
  wire[2:0] RocketTile_io_tilelink_acquire_bits_payload_subword_addr;
  wire[3:0] RocketTile_io_tilelink_acquire_bits_payload_atomic_opcode;
  wire RocketTile_io_tilelink_grant_ready;
  wire RocketTile_io_tilelink_finish_valid;
  wire[1:0] RocketTile_io_tilelink_finish_bits_header_src;
  wire[1:0] RocketTile_io_tilelink_finish_bits_header_dst;
  wire[2:0] RocketTile_io_tilelink_finish_bits_payload_master_xact_id;
  wire RocketTile_io_tilelink_probe_ready;
  wire RocketTile_io_tilelink_release_valid;
  wire[1:0] RocketTile_io_tilelink_release_bits_header_src;
  wire[1:0] RocketTile_io_tilelink_release_bits_header_dst;
  wire[25:0] RocketTile_io_tilelink_release_bits_payload_addr;
  wire[1:0] RocketTile_io_tilelink_release_bits_payload_client_xact_id;
  wire[2:0] RocketTile_io_tilelink_release_bits_payload_master_xact_id;
  wire[511:0] RocketTile_io_tilelink_release_bits_payload_data;
  wire[2:0] RocketTile_io_tilelink_release_bits_payload_r_type;
  wire RocketTile_io_host_pcr_req_ready;
  wire RocketTile_io_host_pcr_rep_valid;
  wire[63:0] RocketTile_io_host_pcr_rep_bits;
  wire RocketTile_io_host_ipi_req_valid;
  wire RocketTile_io_host_ipi_req_bits;
  wire RocketTile_io_host_ipi_rep_ready;
  wire RocketTile_io_host_debug_stats_pcr;
  wire RocketTile_io_temac_rx_axis_fifo_tready;
  wire[7:0] RocketTile_io_temac_tx_axis_fifo_tdata;
  wire RocketTile_io_temac_tx_axis_fifo_tvalid;
  wire RocketTile_io_temac_tx_axis_fifo_tlast;
  wire[11:0] RocketTile_io_temac_s_axi_awaddr;
  wire RocketTile_io_temac_s_axi_awvalid;
  wire[31:0] RocketTile_io_temac_s_axi_wdata;
  wire RocketTile_io_temac_s_axi_wvalid;
  wire RocketTile_io_temac_s_axi_bready;
  wire[11:0] RocketTile_io_temac_s_axi_araddr;
  wire RocketTile_io_temac_s_axi_arvalid;
  wire RocketTile_io_temac_s_axi_rready;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_pcr;
  wire uncore_io_mem_req_cmd_valid;
  wire[25:0] uncore_io_mem_req_cmd_bits_addr;
  wire[4:0] uncore_io_mem_req_cmd_bits_tag;
  wire uncore_io_mem_req_cmd_bits_rw;
  wire uncore_io_mem_req_data_valid;
  wire[127:0] uncore_io_mem_req_data_bits_data;
  wire uncore_io_tiles_0_acquire_ready;
  wire uncore_io_tiles_0_grant_valid;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_src;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_dst;
  wire[511:0] uncore_io_tiles_0_grant_bits_payload_data;
  wire[1:0] uncore_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[2:0] uncore_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_g_type;
  wire uncore_io_tiles_0_finish_ready;
  wire uncore_io_tiles_0_probe_valid;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_src;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_dst;
  wire[25:0] uncore_io_tiles_0_probe_bits_payload_addr;
  wire[2:0] uncore_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[1:0] uncore_io_tiles_0_probe_bits_payload_p_type;
  wire uncore_io_tiles_0_release_ready;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_pcr_req_valid;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire[4:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire uncore_io_htif_0_ipi_req_ready;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_rep_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
`endif

  assign resetSigs_0 = uncore_io_htif_0_reset;
  assign io_temac_s_axi_rready = RocketTile_io_temac_s_axi_rready;
  assign io_temac_s_axi_arvalid = RocketTile_io_temac_s_axi_arvalid;
  assign io_temac_s_axi_araddr = RocketTile_io_temac_s_axi_araddr;
  assign io_temac_s_axi_bready = RocketTile_io_temac_s_axi_bready;
  assign io_temac_s_axi_wvalid = RocketTile_io_temac_s_axi_wvalid;
  assign io_temac_s_axi_wdata = RocketTile_io_temac_s_axi_wdata;
  assign io_temac_s_axi_awvalid = RocketTile_io_temac_s_axi_awvalid;
  assign io_temac_s_axi_awaddr = RocketTile_io_temac_s_axi_awaddr;
  assign io_temac_tx_axis_fifo_tlast = RocketTile_io_temac_tx_axis_fifo_tlast;
  assign io_temac_tx_axis_fifo_tvalid = RocketTile_io_temac_tx_axis_fifo_tvalid;
  assign io_temac_tx_axis_fifo_tdata = RocketTile_io_temac_tx_axis_fifo_tdata;
  assign io_temac_rx_axis_fifo_tready = RocketTile_io_temac_rx_axis_fifo_tready;
  assign io_mem_req_data_bits_data = uncore_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = uncore_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = uncore_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = uncore_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = uncore_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = uncore_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = uncore_io_host_debug_stats_pcr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  RocketTile RocketTile(.clk(clk), .reset(resetSigs_0),
       .io_tilelink_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tilelink_acquire_valid( RocketTile_io_tilelink_acquire_valid ),
       .io_tilelink_acquire_bits_header_src( RocketTile_io_tilelink_acquire_bits_header_src ),
       .io_tilelink_acquire_bits_header_dst( RocketTile_io_tilelink_acquire_bits_header_dst ),
       .io_tilelink_acquire_bits_payload_addr( RocketTile_io_tilelink_acquire_bits_payload_addr ),
       .io_tilelink_acquire_bits_payload_client_xact_id( RocketTile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tilelink_acquire_bits_payload_data( RocketTile_io_tilelink_acquire_bits_payload_data ),
       .io_tilelink_acquire_bits_payload_a_type( RocketTile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tilelink_acquire_bits_payload_write_mask( RocketTile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tilelink_acquire_bits_payload_subword_addr( RocketTile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tilelink_acquire_bits_payload_atomic_opcode( RocketTile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tilelink_grant_ready( RocketTile_io_tilelink_grant_ready ),
       .io_tilelink_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tilelink_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tilelink_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tilelink_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tilelink_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tilelink_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tilelink_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tilelink_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tilelink_finish_valid( RocketTile_io_tilelink_finish_valid ),
       .io_tilelink_finish_bits_header_src( RocketTile_io_tilelink_finish_bits_header_src ),
       .io_tilelink_finish_bits_header_dst( RocketTile_io_tilelink_finish_bits_header_dst ),
       .io_tilelink_finish_bits_payload_master_xact_id( RocketTile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tilelink_probe_ready( RocketTile_io_tilelink_probe_ready ),
       .io_tilelink_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tilelink_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tilelink_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tilelink_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tilelink_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tilelink_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tilelink_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tilelink_release_valid( RocketTile_io_tilelink_release_valid ),
       .io_tilelink_release_bits_header_src( RocketTile_io_tilelink_release_bits_header_src ),
       .io_tilelink_release_bits_header_dst( RocketTile_io_tilelink_release_bits_header_dst ),
       .io_tilelink_release_bits_payload_addr( RocketTile_io_tilelink_release_bits_payload_addr ),
       .io_tilelink_release_bits_payload_client_xact_id( RocketTile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tilelink_release_bits_payload_master_xact_id( RocketTile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tilelink_release_bits_payload_data( RocketTile_io_tilelink_release_bits_payload_data ),
       .io_tilelink_release_bits_payload_r_type( RocketTile_io_tilelink_release_bits_payload_r_type ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( RocketTile_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_0_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_0_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( RocketTile_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( RocketTile_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( RocketTile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( RocketTile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_pcr( RocketTile_io_host_debug_stats_pcr ),
       .io_temac_rx_axis_fifo_tdata( io_temac_rx_axis_fifo_tdata ),
       .io_temac_rx_axis_fifo_tvalid( io_temac_rx_axis_fifo_tvalid ),
       .io_temac_rx_axis_fifo_tready( RocketTile_io_temac_rx_axis_fifo_tready ),
       .io_temac_rx_axis_fifo_tlast( io_temac_rx_axis_fifo_tlast ),
       .io_temac_tx_axis_fifo_tdata( RocketTile_io_temac_tx_axis_fifo_tdata ),
       .io_temac_tx_axis_fifo_tvalid( RocketTile_io_temac_tx_axis_fifo_tvalid ),
       .io_temac_tx_axis_fifo_tready( io_temac_tx_axis_fifo_tready ),
       .io_temac_tx_axis_fifo_tlast( RocketTile_io_temac_tx_axis_fifo_tlast ),
       .io_temac_s_axi_awaddr( RocketTile_io_temac_s_axi_awaddr ),
       .io_temac_s_axi_awvalid( RocketTile_io_temac_s_axi_awvalid ),
       .io_temac_s_axi_awready( io_temac_s_axi_awready ),
       .io_temac_s_axi_wdata( RocketTile_io_temac_s_axi_wdata ),
       .io_temac_s_axi_wvalid( RocketTile_io_temac_s_axi_wvalid ),
       .io_temac_s_axi_wready( io_temac_s_axi_wready ),
       .io_temac_s_axi_bresp( io_temac_s_axi_bresp ),
       .io_temac_s_axi_bvalid( io_temac_s_axi_bvalid ),
       .io_temac_s_axi_bready( RocketTile_io_temac_s_axi_bready ),
       .io_temac_s_axi_araddr( RocketTile_io_temac_s_axi_araddr ),
       .io_temac_s_axi_arvalid( RocketTile_io_temac_s_axi_arvalid ),
       .io_temac_s_axi_arready( io_temac_s_axi_arready ),
       .io_temac_s_axi_rdata( io_temac_s_axi_rdata ),
       .io_temac_s_axi_rresp( io_temac_s_axi_rresp ),
       .io_temac_s_axi_rvalid( io_temac_s_axi_rvalid ),
       .io_temac_s_axi_rready( RocketTile_io_temac_s_axi_rready )
  );
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_pcr( uncore_io_host_debug_stats_pcr ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( uncore_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( uncore_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( uncore_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( uncore_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( uncore_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( uncore_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_tiles_0_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( RocketTile_io_tilelink_acquire_valid ),
       .io_tiles_0_acquire_bits_header_src( RocketTile_io_tilelink_acquire_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( RocketTile_io_tilelink_acquire_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( RocketTile_io_tilelink_acquire_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( RocketTile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( RocketTile_io_tilelink_acquire_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( RocketTile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( RocketTile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( RocketTile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( RocketTile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( RocketTile_io_tilelink_grant_ready ),
       .io_tiles_0_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( RocketTile_io_tilelink_finish_valid ),
       .io_tiles_0_finish_bits_header_src( RocketTile_io_tilelink_finish_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( RocketTile_io_tilelink_finish_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( RocketTile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( RocketTile_io_tilelink_probe_ready ),
       .io_tiles_0_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( RocketTile_io_tilelink_release_valid ),
       .io_tiles_0_release_bits_header_src( RocketTile_io_tilelink_release_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( RocketTile_io_tilelink_release_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( RocketTile_io_tilelink_release_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( RocketTile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( RocketTile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( RocketTile_io_tilelink_release_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( RocketTile_io_tilelink_release_bits_payload_r_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_0_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_pcr( RocketTile_io_host_debug_stats_pcr ),
       .io_incoherent_0( uncore_io_htif_0_reset )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  `ifndef SYNTHESIS
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
  `endif
  Queue_0 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( RocketTile_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_0_io_deq_bits_data )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_pcr_rep_valid ),
       .io_enq_bits( RocketTile_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_ipi_req_valid ),
       .io_enq_bits( RocketTile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [6:0] W0A,
  input W0E,
  input [83:0] W0I,
  input [83:0] W0M,
  input [6:0] R1A,
  input R1E,
  output [83:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<4; i=i+21) begin
    for (j=1; j<21; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [83:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
    end
  `endif
  reg [6:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][20:0] <= W0I[20:0];
  if (W0E && W0M[21]) ram[W0A][41:21] <= W0I[41:21];
  if (W0E && W0M[42]) ram[W0A][62:42] <= W0I[62:42];
  if (W0E && W0M[63]) ram[W0A][83:63] <= W0I[83:63];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [6:0] RW0A,
  input RW0E,
  input RW0W,
  input [37:0] RW0M,
  input [37:0] RW0I,
  output [37:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+19) begin
    for (j=1; j<19; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [37:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {2 {$random}};
    end
  `endif
  reg [6:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][18:0] <= RW0I[18:0];
  if (RW0E && RW0W && RW0M[19]) ram[RW0A][37:19] <= RW0I[37:19];
end
assign RW0O = ram[reg_RW0A];

endmodule


module HellaFlowQueue_ram(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [132:0] W0I,
  input [5:0] R1A,
  input R1E,
  output [132:0] R1O
);

reg [132:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {5 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module DataArray_T6(
  input CLK,
  input RST,
  input init,
  input [8:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [8:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [511:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [8:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_T157(
  input CLK,
  input RST,
  input init,
  input [8:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [511:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [8:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


